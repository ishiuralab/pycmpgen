module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd22b34e767208bd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1a55ff12dabb4bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h960ed8d8b4fcc41b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2295a07da58876e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h518679ccffc503b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcfc827006c9b2a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f114de6b1c0a680;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca0ccd448ea6fb1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h112a92b51ea32b9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h281430ef7e900b36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he94e0e8ba39c7652;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9976e21c1c09f3d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e641d5d72aea462;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbeb3391bab0d2c07;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74654824590085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4feb9a97006fc58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1b6fa6a825ac84b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9df254277c53c8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha851d47f28a3af02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacb04b8dededc216;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50bac01f8f8971a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h522c721ffd906ebf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe2273ffcee70060;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53a4f8139b62331a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h830a1fd1a53655b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a75d8d31fa6d211;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82505f9a993fed3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ae3bf283c466761;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7942ff7b85060536;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1006efeb53361100;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd64324837cd35053;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf563ff6d06b4fb10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf3e56e64e139397;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce442a43990b5e0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fd5a20015b587fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d2ca4a9a91c8a80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he196eb2810d184b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a34b7f6b2de2deb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0fa8bc5314185e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1b3eb9d727a81f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ab5f89ed9d2ca7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c9033a42a544b7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79a3c4c78365fc83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55ebe98b992b7de9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h578124bb547bf1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b7f1c489acf59d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf44d487ab8307789;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8bf458bf7924bbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86ca60afbedd8a5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4326ded1d6a0fca4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48b1b9078c902c16;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22ca9792d2607725;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee49151ad3a6c9b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd67111515811d0a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fa337e7a145fafb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b13c4e2e17783c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb5f9093593823b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20122add0d052754;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26e4961d3d1f7f8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ba1679379c7af1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3efd2feb00faf96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h785d233d4bd6e51e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d0d67c4cb011e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef2f712876094536;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h992579324e809d78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3caca32c5c5325c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc50c45ee6b6f5657;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23d527d14565476c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec9153332216bb10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf6ea82a3cfc0209;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf96b50b03829a43c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcea00d18b09a0aaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c5fcbee8eb6b060;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef1fbdc1dd8355b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b39ae12884cbfab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9b32ba344f8279d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3732e6b019b6e83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3272d7d6ac2f2801;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4285595ddfe42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h969879ca7691ee1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc037c9ad9daf1dc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95d5ad7853f89ab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a4cc896239921d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd90cf425e496008b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h148ace7286b8eb7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd52269b0324ead50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h827eb2ffc6fd7b67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba12ec144b0518;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha07e93d656d53e7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec144ab52beb55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f429ab74012c211;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43456a65a2fe77ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h399e7fdf23e4f36a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaf1de6771d00add;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd11a0634886f65ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb557222fe8d59aaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb286c7900fd7cfd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h503dd32dca16535e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h340a5b81048599b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b2a45c95b0c902e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f9d27d76eb96d58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h370af7e62c21ae75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b91b98b546959cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d02d02a67878c7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefa28e9b8e33fd62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ceda826651d1f28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17229a5bba3a9196;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12cf13f1d6f01965;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h394d704d3f259fdf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bd3b0be70f3db13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h926c6b2bccabf53a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h749a1ae0c45e06f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44ecd118648aa893;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7dadeed9eacb25c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf014abcd9ae6a0cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h387322d75da90fe1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5321734b7ab8acb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd61f625e16735b1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8503fcd0cea16644;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h917d72276e6de758;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf39a576581e460e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7992b87c94a56ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeb8327d2d9e2615;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ceb2e96df68cee5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2939d902af974193;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d7f1081ecfb157c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f49e4ff5411003a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h132e134466638469;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1d56ad749d9962f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ac8e07b11ef6620;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf84190517fcb24bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had94ebb45d842100;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a59715d045c3bbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdad225b7e6f6887f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb0dbb21cb313fda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cff709cd56a239d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f22eeb041c42667;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe0f99d81ae641f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc307f649d3a9423b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0346ac234cd6452;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha715500109ee37d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97fbaa17d6a1ad9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd7d193dd967161d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf17b1e3d515eb141;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dffd6c0d29f4ebb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc123645ea3fbe660;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had4b3ccbe56385b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfd7e07ad84ec4f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1b47c04b04a0b4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71c85935ac2808d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1da9722a1d719e45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2eb37161ceece6c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce50dcfcc36d92f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6120be31f35c9da3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48e906b46efbac0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66b19ef07c6ac4e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcde542ebe0cad69f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea3ca9f5343763a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed6a5179f567d4e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde65a21296a53974;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e3f24ca40eec9aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h911afaa9804545f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42b00ca7a8fae369;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h609f68d9ee70d682;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5359ffc562fc993;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda34dabe0e5429fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d016c4feeec8257;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9d3eb8beaa3ee0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1265029960d3e0ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3892ed46250855e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54831aa78ed8fda2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37e35f42cce23e83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a5fca22d13de72a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h224df9060967623e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea3c7b5fa9b77c04;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d3589282e7e945e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1179391d86b4a79a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85782c27ba383b8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2f2b82a9bf3e5a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fdf37c648d63023;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81e35540a4309bc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c12b9222be24a87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79db011fd2bdf0b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60daa5c921d1faa6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdca80da262af6979;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99b9ff09c84f82e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc151eea6cc8ef08b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e9c87327fdf4c01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4341a0eb2bf5e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0bf27ca78ea4243;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf05658178caa288;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36511abcccc2ee9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha31a14c9d49d9efa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h707be90317bd7803;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1b4e9c7c9b78c6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6308a72f74b53f22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dba27566e5391d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaf2c16124d08e5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he83488cbf5b176f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h744a31a229a9e633;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9dea78d856edc47c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h831fe6205c30c9c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h313f5064dfee9f7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30639ee833a93124;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b82c47cc635ebe3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8ac80e851efe23a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ad8ea46047c03d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6ee4bd74415ee17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3ef0a72a5ee3aee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b8de2c5c655f0e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6297e0e7136d987;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53a9dad3293061c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c5a047e415ee193;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf936ff89e78c82f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde52f354b24e8f72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a1fa3ece6b2e97c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8afeae9468e6d9e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde272075ddec54ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedd663005d3c0a34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2ead107e171215b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d44c2d0a5084ebe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h613c7688aeef274f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ee20c49e4317a90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc81599943fb7b2d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fa75e2d90e92f83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2236823d3ee6a9e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefc30def23f6cfc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf466ac6600bd8ebe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d718cb5a79e37e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21b6089bc43b1f70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h338e2b4e0d4bb8fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86e70a6c828c7014;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h316ff7dbdacf4e72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e57cfdd818af081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he360ff232aa3408e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h644e2611a46ea2d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h587c84b092843691;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc641b39b9e6c1e0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d721fb407263ad6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cd484391041580b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6f352f10ec3ff08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h353ab3f5a11cfbe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0e79d2231b52744;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf60eb06bae2e2aa5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2b7a594bcfb63cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haea85b923ac9d2cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2fe1a8ff4dda5da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5355a02fc5c2f4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd269736e7e7c8114;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd6549d3f93c8b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7237522ca990faf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h378f4d11d6d0d050;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8399331b95dc90ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd090d05fee78e39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f25afbe0165a2f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h964f817c9b3f28f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f945f641538963d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceb6698ec7990968;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7df7f380defb44e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93d9a0d0e23a9fa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf58054cea3d69b37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30efef79990bdb1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93915094879cae18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he65982969b7c0a67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had85e0b3a6c85394;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f0658106c46a273;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haccf60d56d2ee42b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a43bc5d6d6d0aee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6256cb3e555511b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1534f218c520d2cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc53ce7d294a77e43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h609740c033a1083e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c8fb5a7e59084e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16fb7b634c1eb0ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25bdc689de0525e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe5f52084a5d9c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b340c417c3994c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h375784e68a0ff3c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f2b443ecd66234;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1c0f9fc53d28f98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea9e3f7386863c8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49344fdf7e34d2e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dbda7d923540919;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9d154ad63dad8c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d2865133ee6a2be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ff409c8a79ee68d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h190e97bc6dbdb030;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50768839f65811cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40c4c34fdc6d4305;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d6bdee644254180;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7443f55c2f948c06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef53099fdb616c67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb38fa20421576ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb45a978eeaa5a91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf5b7058d2abea10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdecdf1572cc479f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe6769aa64a3fa8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd39d94231e93bbc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3908d68787e0152;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h417308197a59b43d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4a977c23e0ac742;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h680987dbf429b240;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ab92a998317b012;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99d914db987b2bcc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h681420c8533a5b7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha72d2740f2586340;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd135e1f79ebc787a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6be5349163db399;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h300f620ce9a7abdf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80dda5f7bb6232c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed5aa02a3c36b596;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2692814bd87d970a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb50dd28d5345c135;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fd0c519619f0c2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdff4d9a2085445a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e824673a2cbbd3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha17ffa7cbf2c1043;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6176aa805b3f971;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73f01021106f3822;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38fa1d64168726c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ddf81010d4a394a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ec0140cec83f1c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aa1fdf3d065225c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h406473474e7f083c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde44ab029a3ec7bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb44b6a78e3229b9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99695fd65847be6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bb5c844a49587a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h217795e25a60b525;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1189d756e013e64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69fb62393d432dca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he55388d73e701fb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57190229b9ec38cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe46d0c2af016a39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc784379a31e2344;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb42eccbb2232164f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf26894e392857d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f108db7411fffc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1fd670d45328824;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb73f2e83d9599d80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16034b93383e76e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7140f9397252c9af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb19553956556a8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5079dcd1b7de779;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50b9388b2b29268a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h331992782597179;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h787dad41887d9021;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaa165c195fd1b8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93008f0fdb2d7f05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92d3a204c08ea45f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45a0bf66ad5037d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43ea92bc8808d35f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4e7e650d806bbea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b1c5ebbff9fcb59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5d69d3ebd84556e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63a07bc39e27672f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h418e9eb7704fd771;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb23b7935702db232;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e63bf27ebe514d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b0f32880f6b1551;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h519cb95b6a201bf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7b8334fa9369e31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcde3ae28c42ca467;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42b66507fb998dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99d06f00219f1bf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h255ebe6adefc582d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2529a85f564a9dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf18b631f2d1542ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dc51e27ff6387c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfde01b9585af894;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha78d52e192d72aaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3bb18336ece7c79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fdd38caee3a1732;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha104841187118898;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4e8859188e35c7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2ca4ebb92c1b466;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45d5355bf1618c71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heab37ed10573b71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb13390af2c96db45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae331eb585aebda1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcee389d21f9a6d38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7741cc795e255bdf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16a1fbf7eaa800b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e515b15121c8dda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fb2709df8eb884c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80359f7fa8af4400;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h774d0ebaf8b15c32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfce8fe845ffb73d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62639def819c8513;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h869d0773d0c738cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4199bd857289797;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74c5b31e451e657d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f22286466a34df8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6257100786fe09f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h368707ed071886f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaea7f1ffe6b2a53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dcf5cc7aa436b58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105d9c2187152557;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdac4e74ab8dc481;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75358f1a186f0652;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h493440d561e42d8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ae111dac87cf534;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb234b5817227f33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef339ec657507da4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d6bd870d209b908;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h654558b1e9453cc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23145f0d4cc0ce9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb683372daad6ff5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39e28cbccf00c08e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4eb8b819d904878;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ecad497ae5d6282;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58053d46a2212023;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fe4e8a481c22c19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc56afe086cda8d55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d171d4fc2bf490;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f4c6f3558c8bdf1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac4554729ac90485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7ded799e08623f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6abfd69275ab49d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33e2336c8672c932;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee98359e714c5c8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cab237eb992acc2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5c8e11912f48972;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56f10d83838fae74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf252c091f256341f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1a16502f3f7ecbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c2c087a81b4c1ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h414819684612d2e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a324ef8dbb4fdf0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56f1233741d75b92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc60bf6baedfe5bd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b88ddaa9b5a312;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2ee5131821f4145;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96ca377f709a53ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ded6fddf929d6f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he75d9b447156bd01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4dad1789dd3313d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cd9209c0d031c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fe9ffd8e9f66a45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfea3d2c77f953fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4631ba538f09915;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aa53ce3998293b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdf114e62ae3dc8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4d01002bb9b7ad5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11ebc94cbec0b877;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha91c16cb36cfe090;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d945a91539244b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62ab76df94179cbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf400dac5cfc1124;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7114ed96922645e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28f8e45929e748b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab923f7c1124d9a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecf6bc2869446a1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dccff34d489593f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c6cc9b018a596f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17b485b70929f4d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h222943c13c7d6bec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0386481231b4159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa7e72731622959;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c9c033edca5c470;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ea7345b9e058058;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h313785b199f552bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cea6ab55df9287e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53239c7cae18482e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4646fbe8f81cdc9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ed9eac386672b32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e4333586c4b52f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6dfa121391da1229;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e39f484f32aec26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59d2d4e13bab4beb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfee5f5a91d5a8fc6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3c9c22c181b9e8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7bfa1b765cc9dda8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95840708bfc70fba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb652f673f70dea26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f74fc8e326f3fab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb062bbef23ff7287;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb56c2a4432318a26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e0c2f1c44da43c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8a08ac7f61811ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e496f641c877897;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe2638fae6dfdbc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa55f46631e52dd9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8afd947fa1ca9889;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac3a0724306ccb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4750a88d8be47834;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4857e3c80d19fe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd57d433ea4bd409;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf499d3beda071879;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8976b8d4e9523fbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5671172c09457ade;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha29d8e85e3f2d164;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7248b2f4dc985305;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc73b8097f6ff8267;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cb1c0a621d5332d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec297e75fca925fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0b671fe5912b8ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccc1a809f9a79406;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h962a6ec6a8a6ce5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he347e3c300412330;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he23bb262dcc4edc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde15e61de79bad13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2610f5f2561c6820;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6766c17e3f07bd86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habfdef0fc193336a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d146a3aabc8d77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8d8c32021847f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6fdeaca1a232299;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he74c229d51f0c61a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d7d0318d3b490d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6d0e71d62f6371e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa06b3703157150f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57ee8d6bc2196ed6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15f0002c592d2ed0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96ddc92dc96387d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f633253d996767d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a63fd34820a847a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb3e400d7777137d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb76b203d1ac070a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h455152813205f51f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ea56d41fccdad96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29d15f83772187c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc789d398f4b6e51b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaab37e01a690b8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77e8a8239de07b11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15922670fc899b0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f6339be186e4eae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d92a47288a58d82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb38e191af747a1ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a2761c817bc7f51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd9980790614fdc1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd31a6124629125a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb13fd0884ee5cd6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c7636f41903d25b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebc60c9d569320ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12f7b5539903a9c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70479586965754d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8fa5dd4067a9c07;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h372aa996ec0f7b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d78879d867782c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha986f741af6dda34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h107b82e65b4c25b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h988bce2b6304e344;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38e6bdc19e88a612;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66910b3288b868fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadb8adfa4751e728;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3a3d0bd4a2ba06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he76504ffcb3d0a4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h966902399b4b8714;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35191b461cb278d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9203231b2e2f15b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf76f1c176d544ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfe63f7c18155358;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56d44bf4dccbdf3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h912f7b312a5d84b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86a4d19905c674e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2191a8daeaa6f2d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24c538e5dc6ac733;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb98e096810256445;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85fa24eefa294c40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6ed9655eada1ec4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4cd963f0d59588e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55b2a5432cc4a45c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6295b511eed6b4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h598298aac40b5331;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6262beac8411902;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7bf9ca7c28bf0bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h110c517e7e779f65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba0a0467a18a510;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0ee1ff700f9864f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h652c2301a6955a03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb1d5236d92eaa39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27ec58e8cb26126;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79bbcaa3c5396311;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42e1ed3ef1a81290;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7278bdf9073070c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95073f962efa4389;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d51f017dd0946f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9219c553b1577b16;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfd82d57071440e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he20f7a0a0cc97610;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28a8e08f8bfbe1dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h869ae566a024ade1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44b57fbfc853c39a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30c48fbe5ffd326b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74f04746cba87ac0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h659af2456e89d032;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92f0b6e2cb142429;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc458f81105355001;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h138b7f0ffa891191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedb865675af58fed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16e5eeff293fc7de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0c38c84e1ddbee1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2be9208f3278364;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a4cb35887533b99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha306c6fbdf4be64d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f1e162481601ed2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd2ab309ccd19b67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd04c0f0b5123aced;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb84ca38bb94fde55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e8e4d5ea714c0a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9a8de3c3f675e7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5dcabdc31f4bc11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ba0711e6197a513;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8394acaf8a706764;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcfb93d636220e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb095a02343bddc2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32740315b3250bee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c534aa84e4730b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3675fe269706539e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79849f43a0eb6587;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h950361e2ddcef1cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3493e969755ed03e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haefab9400fdbd3f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb9c5bcea7a06f22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd0580d2f6d2baff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59d28abaaec9e927;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb301f4f025ccc45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h167f5fb012b562b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf702b2e981b5721f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h165785e7d9ba5bd1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0aec14e0128fd85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd456407538a43f55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb85c906d390dbf9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heee89c9f54f55c03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfa882129a032f6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38449372468f3a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h630948191efe3229;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd855e37758becc70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7045346c7b2a0d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd44c32616cea7df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe184b7d1688d8ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he83bf23c5eba06bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2a5ed0c9c75f90f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63c963c5d981cf7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b048429c6f493a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bb1ca4b3d990100;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a7be40c621c6918;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7816db03dc0b4ba5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h519da34538b9cbfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53e68b78cfe1c60e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c1f2a7ddeeff753;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99c47f9e327fbce9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd6f1d258b367cb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h945e4788acff1ce8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f7818f400cbfec2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93ff6cebed735240;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4842265d710693ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c2623e713375af9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d05f31062bfdc18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dc7bf67490111e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95f3f2c9e669c36c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4186805e3508a6e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a6db6b65c961af2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habca9c173813df33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9697d31be9132b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a2c2a9bf6d39e19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14478a21c4f381d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60419fe5bea46f46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc37e6e50a73590ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1e43ea44ac41b2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h340d693fc6d7d9e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55a484e9336e925b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h576b898d6ce7b163;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb324394e5e004c89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12b20b5a27234cee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dcca50fb9232ad8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6728bf5324ef12c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73c84337464313c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb86db3a3a05bae08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c5079fe7890ffb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd827139cc2afb0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e749a6e75ce5ffc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb9ddf94a7b4b9bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf1cffc511fa3c31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbedebcedc5da73e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1edf8219ce19555;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6317fc31cc7b5e44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4db32edfbb5c1897;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4772ca0abbaedc12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72587c11d327f2d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf75863390c364270;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h376fec0d4c04519e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he464d2105f3bd908;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24717b62e3f4e787;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a5259b883a8995e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24b5e4ca564ae59a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6aec8dd314c761ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a2d51f46ae6c50a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a25883b66eb3f6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h617273b3936ea7ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34377eadd9f3cc98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd5263694c8271c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54b09f089dc66e85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6ab6346e12329d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25f6e2031a8149a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66907aa4af6aa5f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h851d2de9c99677ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b0fe6d83c28be4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa4d7b46037c1958;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9efeacfa6ecb0052;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fd11e7271501dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7e738b7e240adb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h604f371ede8bbb73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc67bdbe5bde93acb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6712d4b5bae4641d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb30b32d2e8a23ff5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2af7f1cb30cb8fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14d1a49b435b2edf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6e7f5bab1293fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dc1b80c2fb8d2d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec3e9c2123df1179;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba0781b26b12b3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3debbd9c541d46da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacc843b1d16a8c4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48d1a37a3730c4e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb89d09285595abb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3555df657c17f20e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64bb6c6a0ed76c03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b8aaf9e5471ee3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf692ed4592507e70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c7733ac9f1e086;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9a54f4d7953c9e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85d2c178456fcc58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e654b9542657a78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96ecb6d10bccda8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h758322a2434800ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84a7e89662fb413a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dce79b680f8cf21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h336da1f775468228;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80eaf9cf74176abc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93bd863b2f09d663;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1c4a2370074fea1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd2874f8c772cbd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5deea7296892c32a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9576146110ec6bdb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3085f9def0c93cd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22b7f94c375e1561;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78e42c3d22d3d30e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3a0a7f65b986bde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h786964338daec1e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f06e5f6ce645f6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h265ac1ed11bbb5f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca72e7d38fed2fb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb69e9f2162a31470;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8020202f58c1792c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94a4f90b6e930368;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb8467ed63dcd543;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf873a822a912643a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heed55cc94cff2dca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0fcea0d5c87554e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeb216ad52385d67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdb6c801c52ef928;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbf2c242e6fff06f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0c598223d2ea36f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72b3c694b2bd1fe2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h364ddcaa297596ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc73090ce50653459;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f4262bebea50c5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6acd6cdf2f55dae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1406c81ab06c1d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h489156a6c181a4b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he47be4e32392dc62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5b99bc22531f775;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7842c0628c0e10bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h387842111e0c7c7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h727eac13718c1695;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e77cce6a7eb8cf1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e85d485326ac7f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8eadd680d30c8a5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b9e9058bd505ac1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h659e82f83196d29a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce2a61d7a5dde44e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h160e802a2d1145ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a723a430e417a31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf04218f1e434a97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36ebb271778e540f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he28e7acfb8a4a6e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e5a303f2da295bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd16f29c373ef794;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6869d3196d725191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha07b0a790b6940eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9235be4756021bb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91c8273797e92368;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb724e64f60d1a604;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfc71ebd89cd80a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ac7c0a8abe5538f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc81c1d4520f5c8a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc48794ab9bf50dd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h397fc1d09590a694;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4db833e6d106353;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda0ce534e9d1a6bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h141097f1f9182d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec7d21324faac846;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd60648f93e7a098d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa1e46917e5cb1b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87fbdc9a54fb2704;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h379d19389513f82c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc2c032c52a408b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb2e05cd3bae2a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h645fe3d93e79b1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8cdf6bcc98b390a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3722f69859a269e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f2ae29bfc759a87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aa7fa3301ee861d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf45a66e3034d0b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74a158a71f8212eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77af8ea678bda5e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1520c1df91d7d8e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca8f33d01909bb35;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ebe3bb85aa66c17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7d6308ceafa4a05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85d43b78251c8e91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha378db0bd7a0f7a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb346a5db28e90643;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53c7093764852c0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe204855c4ef4d1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b97ed83d2d3bbe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f9ea95cc362dd86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2542801fac92acfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0e4c3d7a8376fe5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21f15ef5640082b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d450bb2fcb66e57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1abae57321532728;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf50b716ddcdb5fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab943389eae1989b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h257b5e4298b1da3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43ad181b4b7c38a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6773a046cd29c80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he57a9ae42f0fa7d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ebede76379a81e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h126abc87563da1f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6ec0376f3555eb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78aa9bb6412d64b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he97258e189f63187;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4390d2bc6ae0793;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc33298cd283a6115;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h837edffbfa08fbda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a97771d87ea869b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64f1be87c5ce8c73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h947d7546720c4d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97a3ba01cb0c33a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ac01cd260c1fbee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfee3d03a69ddbb8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d995bc730a3947b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c535959a803a26a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99b187457c030ca5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he052aa3c9bb415b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c2e073bcd045847;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5e9b1330bbe8a24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2332f89f22a352b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3199c73a0e425d7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5f8f590056a23ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48fd1a549112b290;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h824b3b107845bbe8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49af8dba3c21c4d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb98ee2dfb439efcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71833305539610d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe82b311f2a911fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf04ff357bfbc820;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4430a65e27597501;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h833b49eaf1ea639a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a0ab7cb4b3d1eba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8edfa2e3d23e455;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda304ad828a0025e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3693ec37e20caee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43e192e1f95df780;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83f368131c3e736a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58a592f37318f919;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8e375d56835410;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5901c7c0e08be516;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f46e611b2c98779;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28906b85b11ca15c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fd9fe4dc15d8214;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71f5b6a805d3c2fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f267e800e805b36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h996ec29337d7dbf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6839f8ae19e27f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba817fe12abff2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e99820c1299de86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8b0bbfe12954a24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9ea5a2e24897a03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e2bcd1fab650457;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7f18eab8e0f9dc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6f4d83a6015174d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3873a10d864f3f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe4b0ee4d4c6dbf4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86eb57eac5c3693f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6627b0de2f5d61b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f9eef1ad54d99b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd89b9ce647d3134;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58dd2381ea95e37b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cfbcfb62692d857;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf23fb50b8a9e3c25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he678d843f839ced4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73211f7cda45cc3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8edd21d7a8e392fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14edc423e2875786;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88dab713302cb4bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha111821d52d6394a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h181a0173d3384b1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3286ab214194349;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfea577e10d56874e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7ef8c3d3554e420;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0cf43e1f049cf43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h731daa880e2c82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h478c76fc66417157;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1d64e8946c9765a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb84bbf9f634e4829;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe5261ce57e857ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h891f8cd0c92a87ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aba7c8fa5ffb9df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5cf3c295015084e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51ee6f8b67a4d956;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h299f4f804cd1901d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ddf5ed7fa319b59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fb9e35987dd7b0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0502b8e9b139220;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba7d611b101854c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31c52fe1eaa26493;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf06de031abbe07bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b4d79b9751551da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha730b004b87d21c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha713a9cdafb6f5db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57f7920281e5a4e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94a13033a781e3ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25e78998f22dd970;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd1affea48f754cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa3aa6c9be8e99c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c12f7039c9065b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ce352c13619c18c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf17317488d7b2ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2417f271d14f967b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a3b69596afecf7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h902ccc99e2b35bc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d3f6a97af9726bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8456e62fee948d53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h707ae842acf6269a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb699343349549a91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haab3a47bb66d34a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he64be457222725c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52c77e0ed4cfb216;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f9534cb5250f4b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec2135c8e1d0b18e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h458bc9fb0530e8af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3bdd05a65af7e0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fd05d2a8e93e906;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h480ec4561b9b00ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e256df0b6183184;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef0337b3bbe08a59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27d3e6035453a097;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560a852d82519780;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha807fb1d5b31244a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79a65899d9a3df5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf84ef6804627b3c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e2dd82b0e50effe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd107b5069c9fbd6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36d31973db9259e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5a0b83f5c7ab9d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecb4b7ab39e1bbdb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9ce6080cf1bec14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc83242b31d032ad8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76cc6353d1df37c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h189e0c7c73f22d2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3e7f84d65448fb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h916c23ad13cd761a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h877c531a98239bd2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3db1c6acab8bcda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e7a53427973edcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7191105db77959f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h117d805774ff6beb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ae63179e795e4c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc6714016215ad79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16b74dd06035915e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9185746ee5637774;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30eda5955ed18e6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdff7fa1f72b2ca1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17d526e93b936a3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h559924dcc718d388;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2d9a98a852c9605;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6890e0c2735ca6b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddf1e693cd374d14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac2d8a3a96a6281a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h843f60c0168f60e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7249aebc73e1b73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97e31978756af79c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75a5f1911fbe07a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42f7de3fea3c0618;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae69cab48895b96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h337802a94a3f2507;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73fc99471b6417de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba5c061e548c17d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb05fe664a5edbd47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h513717d8b13935a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0d32ccaadfe89f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdf263f94f53bd64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h794356a94266d615;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b6aa877e37f2798;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc78f8521bd3d82aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h658d80ffda504b74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbcb334e7d9eefe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45b22729c41520b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h316e06876865d36e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0d2d9ed71ac3912;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc64e30dd8d301af2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b3764e163303188;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47888e5fa5ffff8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h638c0e566afc75df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29062d91f0a9d86e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdec8964c1f5c0cac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9279b5e40d2874;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a04ecb247088ad0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb6ad57b2f14e5dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h248cfe807501cb20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h931238b54e8bfeed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45400e69e4406096;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h108e461920cef411;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f555afafbfaf71d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1673953fa48f50c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2312ebc713bf113d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef6d9c692af682c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11651c4581bcd040;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79040a24b53d1827;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ffd1f04e57bddf4;
        #1
        $finish();
    end
endmodule
