module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    compressor_CLA512_16 compressor_CLA512_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA512_16(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [100:0] stage1_0;
   wire [179:0] stage1_1;
   wire [172:0] stage1_2;
   wire [245:0] stage1_3;
   wire [240:0] stage1_4;
   wire [217:0] stage1_5;
   wire [206:0] stage1_6;
   wire [206:0] stage1_7;
   wire [217:0] stage1_8;
   wire [263:0] stage1_9;
   wire [209:0] stage1_10;
   wire [189:0] stage1_11;
   wire [221:0] stage1_12;
   wire [281:0] stage1_13;
   wire [244:0] stage1_14;
   wire [271:0] stage1_15;
   wire [126:0] stage1_16;
   wire [63:0] stage1_17;
   wire [22:0] stage2_0;
   wire [40:0] stage2_1;
   wire [59:0] stage2_2;
   wire [102:0] stage2_3;
   wire [116:0] stage2_4;
   wire [93:0] stage2_5;
   wire [103:0] stage2_6;
   wire [84:0] stage2_7;
   wire [86:0] stage2_8;
   wire [137:0] stage2_9;
   wire [85:0] stage2_10;
   wire [143:0] stage2_11;
   wire [84:0] stage2_12;
   wire [140:0] stage2_13;
   wire [124:0] stage2_14;
   wire [84:0] stage2_15;
   wire [104:0] stage2_16;
   wire [61:0] stage2_17;
   wire [25:0] stage2_18;
   wire [10:0] stage2_19;
   wire [5:0] stage3_0;
   wire [11:0] stage3_1;
   wire [16:0] stage3_2;
   wire [28:0] stage3_3;
   wire [39:0] stage3_4;
   wire [47:0] stage3_5;
   wire [37:0] stage3_6;
   wire [45:0] stage3_7;
   wire [40:0] stage3_8;
   wire [51:0] stage3_9;
   wire [63:0] stage3_10;
   wire [60:0] stage3_11;
   wire [52:0] stage3_12;
   wire [41:0] stage3_13;
   wire [57:0] stage3_14;
   wire [56:0] stage3_15;
   wire [49:0] stage3_16;
   wire [31:0] stage3_17;
   wire [25:0] stage3_18;
   wire [13:0] stage3_19;
   wire [5:0] stage3_20;
   wire [1:0] stage3_21;
   wire [5:0] stage4_0;
   wire [1:0] stage4_1;
   wire [10:0] stage4_2;
   wire [10:0] stage4_3;
   wire [26:0] stage4_4;
   wire [14:0] stage4_5;
   wire [21:0] stage4_6;
   wire [16:0] stage4_7;
   wire [25:0] stage4_8;
   wire [24:0] stage4_9;
   wire [37:0] stage4_10;
   wire [21:0] stage4_11;
   wire [23:0] stage4_12;
   wire [25:0] stage4_13;
   wire [18:0] stage4_14;
   wire [21:0] stage4_15;
   wire [30:0] stage4_16;
   wire [21:0] stage4_17;
   wire [12:0] stage4_18;
   wire [10:0] stage4_19;
   wire [11:0] stage4_20;
   wire [3:0] stage4_21;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [6:0] stage5_2;
   wire [5:0] stage5_3;
   wire [12:0] stage5_4;
   wire [7:0] stage5_5;
   wire [16:0] stage5_6;
   wire [5:0] stage5_7;
   wire [9:0] stage5_8;
   wire [8:0] stage5_9;
   wire [14:0] stage5_10;
   wire [12:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [11:0] stage5_14;
   wire [14:0] stage5_15;
   wire [16:0] stage5_16;
   wire [6:0] stage5_17;
   wire [8:0] stage5_18;
   wire [8:0] stage5_19;
   wire [5:0] stage5_20;
   wire [3:0] stage5_21;
   wire [1:0] stage5_22;
   wire [0:0] stage5_23;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [6:0] stage6_4;
   wire [2:0] stage6_5;
   wire [5:0] stage6_6;
   wire [4:0] stage6_7;
   wire [3:0] stage6_8;
   wire [8:0] stage6_9;
   wire [9:0] stage6_10;
   wire [2:0] stage6_11;
   wire [3:0] stage6_12;
   wire [7:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [7:0] stage6_20;
   wire [4:0] stage6_21;
   wire [1:0] stage6_22;
   wire [0:0] stage6_23;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [2:0] stage7_5;
   wire [0:0] stage7_6;
   wire [5:0] stage7_7;
   wire [0:0] stage7_8;
   wire [2:0] stage7_9;
   wire [6:0] stage7_10;
   wire [2:0] stage7_11;
   wire [1:0] stage7_12;
   wire [2:0] stage7_13;
   wire [4:0] stage7_14;
   wire [3:0] stage7_15;
   wire [1:0] stage7_16;
   wire [6:0] stage7_17;
   wire [2:0] stage7_18;
   wire [1:0] stage7_19;
   wire [3:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [0:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [0:0] stage8_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_1[13]},
      {stage0_2[13]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[14]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[15]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[16]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[17]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[110], stage0_0[111], stage0_0[112]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[18]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[19]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[20]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[21]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[22]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[23]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[128], stage0_0[129], stage0_0[130]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[24]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[25]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[134], stage0_0[135], stage0_0[136]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[26]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[137], stage0_0[138], stage0_0[139]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[27]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[140], stage0_0[141], stage0_0[142]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[28]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[143], stage0_0[144], stage0_0[145]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[29]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[30]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[31]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[32]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[155], stage0_0[156], stage0_0[157]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[33]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[158], stage0_0[159], stage0_0[160]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[34]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[161], stage0_0[162], stage0_0[163]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[35]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[164], stage0_0[165], stage0_0[166]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[36]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[167], stage0_0[168], stage0_0[169]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[37]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[170], stage0_0[171], stage0_0[172]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[38]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[173], stage0_0[174], stage0_0[175]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[39]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[176], stage0_0[177], stage0_0[178]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[40]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[179], stage0_0[180], stage0_0[181]},
      {stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181]},
      {stage0_2[41]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[182], stage0_0[183], stage0_0[184]},
      {stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187]},
      {stage0_2[42]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[185], stage0_0[186], stage0_0[187]},
      {stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193]},
      {stage0_2[43]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[188], stage0_0[189], stage0_0[190]},
      {stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199]},
      {stage0_2[44]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[31],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[32],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[33],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[34],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[35],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[36],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[37],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[38],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[39],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[40],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[41],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[42],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[43],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[44],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[45],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[46],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[47],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[48],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[49],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[50],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[51],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[52],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[53],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[54],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[55],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[56],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[57],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[58],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[59],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[60],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[61],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[62],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[63],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[64],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[65],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[66],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[67],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[68],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[69],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[70],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[71],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[72],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[73],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[74],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[75],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[76],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[77],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[78],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[79],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489], stage0_0[490]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[80],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[81],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[82],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507], stage0_0[508]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[83],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[0],stage1_4[84],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[1],stage1_4[85],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[2],stage1_4[86],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[3],stage1_4[87],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[4],stage1_4[88],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[5],stage1_4[89],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[6],stage1_4[90],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[7],stage1_4[91],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[8],stage1_4[92],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[9],stage1_4[93],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[10],stage1_4[94],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[11],stage1_4[95],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[12],stage1_4[96],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[13],stage1_4[97],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[14],stage1_4[98],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[15],stage1_4[99],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[16],stage1_4[100],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[17],stage1_4[101],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[18],stage1_4[102],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[19],stage1_4[103],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[20],stage1_4[104],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[21],stage1_4[105],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[22],stage1_4[106],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[23],stage1_4[107],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[24],stage1_4[108],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[25],stage1_4[109],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[26],stage1_4[110],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[27],stage1_4[111],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[28],stage1_4[112],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[29],stage1_4[113],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[30],stage1_4[114],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[31],stage1_4[115],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[32],stage1_4[116],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[33],stage1_4[117],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[34],stage1_4[118],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[35],stage1_4[119],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[36],stage1_4[120],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[37],stage1_4[121],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[38],stage1_4[122],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[39],stage1_4[123],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[40],stage1_4[124],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[41],stage1_4[125],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[42],stage1_4[126],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[43],stage1_4[127],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[44],stage1_4[128],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[45],stage1_4[129],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[46],stage1_4[130],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[47],stage1_4[131],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[48],stage1_4[132],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[49],stage1_4[133],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[50],stage1_4[134],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397]},
      {stage0_3[307]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[51],stage1_4[135],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage0_3[308]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[52],stage1_4[136],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_3[309]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[53],stage1_4[137],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412]},
      {stage0_3[310]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[54],stage1_4[138],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417]},
      {stage0_3[311]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[55],stage1_4[139],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage0_3[312]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[56],stage1_4[140],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427]},
      {stage0_3[313]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[57],stage1_4[141],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432]},
      {stage0_3[314]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[58],stage1_4[142],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_3[315]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[59],stage1_4[143],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442]},
      {stage0_3[316]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[60],stage1_4[144],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447]},
      {stage0_3[317]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[61],stage1_4[145],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[448], stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452]},
      {stage0_3[318]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[62],stage1_4[146],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[453], stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457]},
      {stage0_3[319]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[63],stage1_4[147],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462]},
      {stage0_3[320]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[64],stage1_4[148],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_3[321]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[65],stage1_4[149],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472]},
      {stage0_3[322]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[66],stage1_4[150],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[473], stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477]},
      {stage0_3[323]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[67],stage1_4[151],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_2[478], stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482]},
      {stage0_3[324]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[68],stage1_4[152],stage1_3[166],stage1_2[166]}
   );
   gpc615_5 gpc167 (
      {stage0_2[483], stage0_2[484], stage0_2[485], stage0_2[486], stage0_2[487]},
      {stage0_3[325]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[69],stage1_4[153],stage1_3[167],stage1_2[167]}
   );
   gpc615_5 gpc168 (
      {stage0_2[488], stage0_2[489], stage0_2[490], stage0_2[491], stage0_2[492]},
      {stage0_3[326]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[70],stage1_4[154],stage1_3[168],stage1_2[168]}
   );
   gpc615_5 gpc169 (
      {stage0_2[493], stage0_2[494], stage0_2[495], stage0_2[496], stage0_2[497]},
      {stage0_3[327]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[71],stage1_4[155],stage1_3[169],stage1_2[169]}
   );
   gpc615_5 gpc170 (
      {stage0_2[498], stage0_2[499], stage0_2[500], stage0_2[501], stage0_2[502]},
      {stage0_3[328]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[72],stage1_4[156],stage1_3[170],stage1_2[170]}
   );
   gpc615_5 gpc171 (
      {stage0_2[503], stage0_2[504], stage0_2[505], stage0_2[506], stage0_2[507]},
      {stage0_3[329]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[73],stage1_4[157],stage1_3[171],stage1_2[171]}
   );
   gpc615_5 gpc172 (
      {stage0_2[508], stage0_2[509], stage0_2[510], stage0_2[511], 1'b0},
      {stage0_3[330]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[74],stage1_4[158],stage1_3[172],stage1_2[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[75],stage1_4[159],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[76],stage1_4[160],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[77],stage1_4[161],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[78],stage1_4[162],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[79],stage1_4[163],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[80],stage1_4[164],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[81],stage1_4[165],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[82],stage1_4[166],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[83],stage1_4[167],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[84],stage1_4[168],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[85],stage1_4[169],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[86],stage1_4[170],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[87],stage1_4[171],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[88],stage1_4[172],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[89],stage1_4[173],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[90],stage1_4[174],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[91],stage1_4[175],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[92],stage1_4[176],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[93],stage1_4[177],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[94],stage1_4[178],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[95],stage1_4[179],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[96],stage1_4[180],stage1_3[194]}
   );
   gpc615_5 gpc195 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[97],stage1_4[181],stage1_3[195]}
   );
   gpc615_5 gpc196 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[98],stage1_4[182],stage1_3[196]}
   );
   gpc615_5 gpc197 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[99],stage1_4[183],stage1_3[197]}
   );
   gpc615_5 gpc198 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[100],stage1_4[184],stage1_3[198]}
   );
   gpc615_5 gpc199 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[101],stage1_4[185],stage1_3[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[27],stage1_6[56],stage1_5[102],stage1_4[186]}
   );
   gpc606_5 gpc201 (
      {stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[28],stage1_6[57],stage1_5[103],stage1_4[187]}
   );
   gpc606_5 gpc202 (
      {stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[29],stage1_6[58],stage1_5[104],stage1_4[188]}
   );
   gpc606_5 gpc203 (
      {stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[30],stage1_6[59],stage1_5[105],stage1_4[189]}
   );
   gpc606_5 gpc204 (
      {stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[31],stage1_6[60],stage1_5[106],stage1_4[190]}
   );
   gpc606_5 gpc205 (
      {stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[32],stage1_6[61],stage1_5[107],stage1_4[191]}
   );
   gpc606_5 gpc206 (
      {stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[33],stage1_6[62],stage1_5[108],stage1_4[192]}
   );
   gpc606_5 gpc207 (
      {stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[34],stage1_6[63],stage1_5[109],stage1_4[193]}
   );
   gpc606_5 gpc208 (
      {stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[35],stage1_6[64],stage1_5[110],stage1_4[194]}
   );
   gpc606_5 gpc209 (
      {stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[36],stage1_6[65],stage1_5[111],stage1_4[195]}
   );
   gpc606_5 gpc210 (
      {stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[37],stage1_6[66],stage1_5[112],stage1_4[196]}
   );
   gpc606_5 gpc211 (
      {stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[38],stage1_6[67],stage1_5[113],stage1_4[197]}
   );
   gpc606_5 gpc212 (
      {stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[39],stage1_6[68],stage1_5[114],stage1_4[198]}
   );
   gpc606_5 gpc213 (
      {stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[40],stage1_6[69],stage1_5[115],stage1_4[199]}
   );
   gpc606_5 gpc214 (
      {stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[41],stage1_6[70],stage1_5[116],stage1_4[200]}
   );
   gpc606_5 gpc215 (
      {stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[42],stage1_6[71],stage1_5[117],stage1_4[201]}
   );
   gpc606_5 gpc216 (
      {stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[43],stage1_6[72],stage1_5[118],stage1_4[202]}
   );
   gpc606_5 gpc217 (
      {stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[44],stage1_6[73],stage1_5[119],stage1_4[203]}
   );
   gpc606_5 gpc218 (
      {stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[45],stage1_6[74],stage1_5[120],stage1_4[204]}
   );
   gpc606_5 gpc219 (
      {stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[46],stage1_6[75],stage1_5[121],stage1_4[205]}
   );
   gpc606_5 gpc220 (
      {stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[47],stage1_6[76],stage1_5[122],stage1_4[206]}
   );
   gpc606_5 gpc221 (
      {stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[48],stage1_6[77],stage1_5[123],stage1_4[207]}
   );
   gpc606_5 gpc222 (
      {stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[49],stage1_6[78],stage1_5[124],stage1_4[208]}
   );
   gpc606_5 gpc223 (
      {stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[50],stage1_6[79],stage1_5[125],stage1_4[209]}
   );
   gpc606_5 gpc224 (
      {stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[51],stage1_6[80],stage1_5[126],stage1_4[210]}
   );
   gpc606_5 gpc225 (
      {stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[52],stage1_6[81],stage1_5[127],stage1_4[211]}
   );
   gpc606_5 gpc226 (
      {stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[53],stage1_6[82],stage1_5[128],stage1_4[212]}
   );
   gpc606_5 gpc227 (
      {stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[54],stage1_6[83],stage1_5[129],stage1_4[213]}
   );
   gpc606_5 gpc228 (
      {stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[55],stage1_6[84],stage1_5[130],stage1_4[214]}
   );
   gpc606_5 gpc229 (
      {stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[56],stage1_6[85],stage1_5[131],stage1_4[215]}
   );
   gpc606_5 gpc230 (
      {stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[57],stage1_6[86],stage1_5[132],stage1_4[216]}
   );
   gpc606_5 gpc231 (
      {stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[58],stage1_6[87],stage1_5[133],stage1_4[217]}
   );
   gpc606_5 gpc232 (
      {stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[59],stage1_6[88],stage1_5[134],stage1_4[218]}
   );
   gpc606_5 gpc233 (
      {stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[60],stage1_6[89],stage1_5[135],stage1_4[219]}
   );
   gpc606_5 gpc234 (
      {stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[61],stage1_6[90],stage1_5[136],stage1_4[220]}
   );
   gpc606_5 gpc235 (
      {stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[62],stage1_6[91],stage1_5[137],stage1_4[221]}
   );
   gpc615_5 gpc236 (
      {stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_5[162]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[63],stage1_6[92],stage1_5[138],stage1_4[222]}
   );
   gpc615_5 gpc237 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_5[163]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[64],stage1_6[93],stage1_5[139],stage1_4[223]}
   );
   gpc615_5 gpc238 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431]},
      {stage0_5[164]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[65],stage1_6[94],stage1_5[140],stage1_4[224]}
   );
   gpc615_5 gpc239 (
      {stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_5[165]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[66],stage1_6[95],stage1_5[141],stage1_4[225]}
   );
   gpc615_5 gpc240 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_5[166]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[67],stage1_6[96],stage1_5[142],stage1_4[226]}
   );
   gpc615_5 gpc241 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446]},
      {stage0_5[167]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[68],stage1_6[97],stage1_5[143],stage1_4[227]}
   );
   gpc615_5 gpc242 (
      {stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_5[168]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[69],stage1_6[98],stage1_5[144],stage1_4[228]}
   );
   gpc615_5 gpc243 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_5[169]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[70],stage1_6[99],stage1_5[145],stage1_4[229]}
   );
   gpc615_5 gpc244 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461]},
      {stage0_5[170]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[71],stage1_6[100],stage1_5[146],stage1_4[230]}
   );
   gpc615_5 gpc245 (
      {stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_5[171]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[72],stage1_6[101],stage1_5[147],stage1_4[231]}
   );
   gpc615_5 gpc246 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_5[172]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[73],stage1_6[102],stage1_5[148],stage1_4[232]}
   );
   gpc615_5 gpc247 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[173]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[74],stage1_6[103],stage1_5[149],stage1_4[233]}
   );
   gpc615_5 gpc248 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[174]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[75],stage1_6[104],stage1_5[150],stage1_4[234]}
   );
   gpc615_5 gpc249 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[175]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[76],stage1_6[105],stage1_5[151],stage1_4[235]}
   );
   gpc615_5 gpc250 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[176]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[77],stage1_6[106],stage1_5[152],stage1_4[236]}
   );
   gpc615_5 gpc251 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[177]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[78],stage1_6[107],stage1_5[153],stage1_4[237]}
   );
   gpc615_5 gpc252 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[178]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[79],stage1_6[108],stage1_5[154],stage1_4[238]}
   );
   gpc615_5 gpc253 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[179]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[80],stage1_6[109],stage1_5[155],stage1_4[239]}
   );
   gpc615_5 gpc254 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[180]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[81],stage1_6[110],stage1_5[156],stage1_4[240]}
   );
   gpc606_5 gpc255 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[82],stage1_6[111],stage1_5[157]}
   );
   gpc606_5 gpc256 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[83],stage1_6[112],stage1_5[158]}
   );
   gpc606_5 gpc257 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[84],stage1_6[113],stage1_5[159]}
   );
   gpc606_5 gpc258 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[85],stage1_6[114],stage1_5[160]}
   );
   gpc606_5 gpc259 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[86],stage1_6[115],stage1_5[161]}
   );
   gpc606_5 gpc260 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[87],stage1_6[116],stage1_5[162]}
   );
   gpc606_5 gpc261 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[88],stage1_6[117],stage1_5[163]}
   );
   gpc606_5 gpc262 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[89],stage1_6[118],stage1_5[164]}
   );
   gpc606_5 gpc263 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[90],stage1_6[119],stage1_5[165]}
   );
   gpc606_5 gpc264 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[91],stage1_6[120],stage1_5[166]}
   );
   gpc606_5 gpc265 (
      {stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[92],stage1_6[121],stage1_5[167]}
   );
   gpc606_5 gpc266 (
      {stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[93],stage1_6[122],stage1_5[168]}
   );
   gpc606_5 gpc267 (
      {stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[94],stage1_6[123],stage1_5[169]}
   );
   gpc606_5 gpc268 (
      {stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[95],stage1_6[124],stage1_5[170]}
   );
   gpc606_5 gpc269 (
      {stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[96],stage1_6[125],stage1_5[171]}
   );
   gpc606_5 gpc270 (
      {stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[97],stage1_6[126],stage1_5[172]}
   );
   gpc606_5 gpc271 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[98],stage1_6[127],stage1_5[173]}
   );
   gpc606_5 gpc272 (
      {stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[99],stage1_6[128],stage1_5[174]}
   );
   gpc606_5 gpc273 (
      {stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[100],stage1_6[129],stage1_5[175]}
   );
   gpc606_5 gpc274 (
      {stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[101],stage1_6[130],stage1_5[176]}
   );
   gpc606_5 gpc275 (
      {stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[102],stage1_6[131],stage1_5[177]}
   );
   gpc606_5 gpc276 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[103],stage1_6[132],stage1_5[178]}
   );
   gpc606_5 gpc277 (
      {stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[104],stage1_6[133],stage1_5[179]}
   );
   gpc606_5 gpc278 (
      {stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[105],stage1_6[134],stage1_5[180]}
   );
   gpc606_5 gpc279 (
      {stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[106],stage1_6[135],stage1_5[181]}
   );
   gpc606_5 gpc280 (
      {stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[107],stage1_6[136],stage1_5[182]}
   );
   gpc606_5 gpc281 (
      {stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[108],stage1_6[137],stage1_5[183]}
   );
   gpc606_5 gpc282 (
      {stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[109],stage1_6[138],stage1_5[184]}
   );
   gpc606_5 gpc283 (
      {stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[110],stage1_6[139],stage1_5[185]}
   );
   gpc606_5 gpc284 (
      {stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[111],stage1_6[140],stage1_5[186]}
   );
   gpc606_5 gpc285 (
      {stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[112],stage1_6[141],stage1_5[187]}
   );
   gpc606_5 gpc286 (
      {stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[113],stage1_6[142],stage1_5[188]}
   );
   gpc606_5 gpc287 (
      {stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[114],stage1_6[143],stage1_5[189]}
   );
   gpc606_5 gpc288 (
      {stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[115],stage1_6[144],stage1_5[190]}
   );
   gpc606_5 gpc289 (
      {stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[116],stage1_6[145],stage1_5[191]}
   );
   gpc606_5 gpc290 (
      {stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[117],stage1_6[146],stage1_5[192]}
   );
   gpc606_5 gpc291 (
      {stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[118],stage1_6[147],stage1_5[193]}
   );
   gpc606_5 gpc292 (
      {stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[119],stage1_6[148],stage1_5[194]}
   );
   gpc606_5 gpc293 (
      {stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[120],stage1_6[149],stage1_5[195]}
   );
   gpc606_5 gpc294 (
      {stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[121],stage1_6[150],stage1_5[196]}
   );
   gpc606_5 gpc295 (
      {stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[122],stage1_6[151],stage1_5[197]}
   );
   gpc606_5 gpc296 (
      {stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[123],stage1_6[152],stage1_5[198]}
   );
   gpc606_5 gpc297 (
      {stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[124],stage1_6[153],stage1_5[199]}
   );
   gpc606_5 gpc298 (
      {stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[125],stage1_6[154],stage1_5[200]}
   );
   gpc606_5 gpc299 (
      {stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[126],stage1_6[155],stage1_5[201]}
   );
   gpc606_5 gpc300 (
      {stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[127],stage1_6[156],stage1_5[202]}
   );
   gpc606_5 gpc301 (
      {stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[128],stage1_6[157],stage1_5[203]}
   );
   gpc606_5 gpc302 (
      {stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[129],stage1_6[158],stage1_5[204]}
   );
   gpc606_5 gpc303 (
      {stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[130],stage1_6[159],stage1_5[205]}
   );
   gpc606_5 gpc304 (
      {stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[131],stage1_6[160],stage1_5[206]}
   );
   gpc606_5 gpc305 (
      {stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[105],stage1_7[132],stage1_6[161],stage1_5[207]}
   );
   gpc606_5 gpc306 (
      {stage0_5[487], stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[106],stage1_7[133],stage1_6[162],stage1_5[208]}
   );
   gpc606_5 gpc307 (
      {stage0_5[493], stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[107],stage1_7[134],stage1_6[163],stage1_5[209]}
   );
   gpc606_5 gpc308 (
      {stage0_5[499], stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[108],stage1_7[135],stage1_6[164],stage1_5[210]}
   );
   gpc615_5 gpc309 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[324]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[54],stage1_8[109],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc310 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[325]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[55],stage1_8[110],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc311 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[326]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[56],stage1_8[111],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc312 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[327]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[57],stage1_8[112],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc313 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[328]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[58],stage1_8[113],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc314 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[329]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[59],stage1_8[114],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc315 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[330]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[60],stage1_8[115],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc316 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[331]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[61],stage1_8[116],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc317 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[332]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[62],stage1_8[117],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc318 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[333]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[63],stage1_8[118],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc319 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[334]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[64],stage1_8[119],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc320 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[335]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[65],stage1_8[120],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc321 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[336]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[66],stage1_8[121],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc322 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[337]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[67],stage1_8[122],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc323 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[338]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[68],stage1_8[123],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc324 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[339]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[69],stage1_8[124],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc325 (
      {stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414]},
      {stage0_7[340]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[70],stage1_8[125],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc326 (
      {stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage0_7[341]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[71],stage1_8[126],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc327 (
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424]},
      {stage0_7[342]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[72],stage1_8[127],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc328 (
      {stage0_6[425], stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429]},
      {stage0_7[343]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[73],stage1_8[128],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc329 (
      {stage0_6[430], stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434]},
      {stage0_7[344]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[74],stage1_8[129],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc330 (
      {stage0_6[435], stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439]},
      {stage0_7[345]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[75],stage1_8[130],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc331 (
      {stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444]},
      {stage0_7[346]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[76],stage1_8[131],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc332 (
      {stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage0_7[347]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[77],stage1_8[132],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc333 (
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454]},
      {stage0_7[348]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[78],stage1_8[133],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc334 (
      {stage0_6[455], stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459]},
      {stage0_7[349]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[79],stage1_8[134],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc335 (
      {stage0_6[460], stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464]},
      {stage0_7[350]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[80],stage1_8[135],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc336 (
      {stage0_6[465], stage0_6[466], stage0_6[467], stage0_6[468], stage0_6[469]},
      {stage0_7[351]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[81],stage1_8[136],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc337 (
      {stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473], stage0_6[474]},
      {stage0_7[352]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[82],stage1_8[137],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc338 (
      {stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_7[353]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[83],stage1_8[138],stage1_7[165],stage1_6[194]}
   );
   gpc615_5 gpc339 (
      {stage0_6[480], stage0_6[481], stage0_6[482], stage0_6[483], stage0_6[484]},
      {stage0_7[354]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[84],stage1_8[139],stage1_7[166],stage1_6[195]}
   );
   gpc615_5 gpc340 (
      {stage0_6[485], stage0_6[486], stage0_6[487], stage0_6[488], stage0_6[489]},
      {stage0_7[355]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[85],stage1_8[140],stage1_7[167],stage1_6[196]}
   );
   gpc615_5 gpc341 (
      {stage0_6[490], stage0_6[491], stage0_6[492], stage0_6[493], stage0_6[494]},
      {stage0_7[356]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[86],stage1_8[141],stage1_7[168],stage1_6[197]}
   );
   gpc615_5 gpc342 (
      {stage0_6[495], stage0_6[496], stage0_6[497], stage0_6[498], stage0_6[499]},
      {stage0_7[357]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[87],stage1_8[142],stage1_7[169],stage1_6[198]}
   );
   gpc615_5 gpc343 (
      {stage0_6[500], stage0_6[501], stage0_6[502], stage0_6[503], stage0_6[504]},
      {stage0_7[358]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[88],stage1_8[143],stage1_7[170],stage1_6[199]}
   );
   gpc606_5 gpc344 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[35],stage1_9[89],stage1_8[144],stage1_7[171]}
   );
   gpc606_5 gpc345 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[36],stage1_9[90],stage1_8[145],stage1_7[172]}
   );
   gpc606_5 gpc346 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[37],stage1_9[91],stage1_8[146],stage1_7[173]}
   );
   gpc606_5 gpc347 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[38],stage1_9[92],stage1_8[147],stage1_7[174]}
   );
   gpc606_5 gpc348 (
      {stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[39],stage1_9[93],stage1_8[148],stage1_7[175]}
   );
   gpc606_5 gpc349 (
      {stage0_7[389], stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[40],stage1_9[94],stage1_8[149],stage1_7[176]}
   );
   gpc606_5 gpc350 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[41],stage1_9[95],stage1_8[150],stage1_7[177]}
   );
   gpc606_5 gpc351 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[42],stage1_9[96],stage1_8[151],stage1_7[178]}
   );
   gpc606_5 gpc352 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[43],stage1_9[97],stage1_8[152],stage1_7[179]}
   );
   gpc606_5 gpc353 (
      {stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[44],stage1_9[98],stage1_8[153],stage1_7[180]}
   );
   gpc606_5 gpc354 (
      {stage0_7[419], stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[45],stage1_9[99],stage1_8[154],stage1_7[181]}
   );
   gpc606_5 gpc355 (
      {stage0_7[425], stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[46],stage1_9[100],stage1_8[155],stage1_7[182]}
   );
   gpc606_5 gpc356 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[47],stage1_9[101],stage1_8[156],stage1_7[183]}
   );
   gpc606_5 gpc357 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[48],stage1_9[102],stage1_8[157],stage1_7[184]}
   );
   gpc606_5 gpc358 (
      {stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[49],stage1_9[103],stage1_8[158],stage1_7[185]}
   );
   gpc606_5 gpc359 (
      {stage0_7[449], stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[50],stage1_9[104],stage1_8[159],stage1_7[186]}
   );
   gpc606_5 gpc360 (
      {stage0_7[455], stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[51],stage1_9[105],stage1_8[160],stage1_7[187]}
   );
   gpc615_5 gpc361 (
      {stage0_7[461], stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465]},
      {stage0_8[210]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[52],stage1_9[106],stage1_8[161],stage1_7[188]}
   );
   gpc615_5 gpc362 (
      {stage0_7[466], stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470]},
      {stage0_8[211]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[53],stage1_9[107],stage1_8[162],stage1_7[189]}
   );
   gpc615_5 gpc363 (
      {stage0_7[471], stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475]},
      {stage0_8[212]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[54],stage1_9[108],stage1_8[163],stage1_7[190]}
   );
   gpc615_5 gpc364 (
      {stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480]},
      {stage0_8[213]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[55],stage1_9[109],stage1_8[164],stage1_7[191]}
   );
   gpc615_5 gpc365 (
      {stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_8[214]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[56],stage1_9[110],stage1_8[165],stage1_7[192]}
   );
   gpc615_5 gpc366 (
      {stage0_7[486], stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490]},
      {stage0_8[215]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[57],stage1_9[111],stage1_8[166],stage1_7[193]}
   );
   gpc615_5 gpc367 (
      {stage0_7[491], stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495]},
      {stage0_8[216]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[58],stage1_9[112],stage1_8[167],stage1_7[194]}
   );
   gpc615_5 gpc368 (
      {stage0_7[496], stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500]},
      {stage0_8[217]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[59],stage1_9[113],stage1_8[168],stage1_7[195]}
   );
   gpc606_5 gpc369 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[25],stage1_10[60],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc370 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[26],stage1_10[61],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc371 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[27],stage1_10[62],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc372 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[28],stage1_10[63],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc373 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[29],stage1_10[64],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc374 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[30],stage1_10[65],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc375 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[31],stage1_10[66],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc376 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[32],stage1_10[67],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc377 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[33],stage1_10[68],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc378 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[34],stage1_10[69],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc379 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[35],stage1_10[70],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc380 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[36],stage1_10[71],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc381 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[37],stage1_10[72],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc382 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[38],stage1_10[73],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc383 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[39],stage1_10[74],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc384 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[40],stage1_10[75],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc385 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[41],stage1_10[76],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc386 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[42],stage1_10[77],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc387 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[43],stage1_10[78],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc388 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[44],stage1_10[79],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc389 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[45],stage1_10[80],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc390 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[46],stage1_10[81],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc391 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[47],stage1_10[82],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc392 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[48],stage1_10[83],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc393 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[49],stage1_10[84],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc394 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[50],stage1_10[85],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc395 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[51],stage1_10[86],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc396 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[52],stage1_10[87],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc397 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[53],stage1_10[88],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc398 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[54],stage1_10[89],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc399 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[55],stage1_10[90],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc400 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[56],stage1_10[91],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc401 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[57],stage1_10[92],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc402 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[58],stage1_10[93],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc403 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[59],stage1_10[94],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc404 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[60],stage1_10[95],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc405 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[61],stage1_10[96],stage1_9[150],stage1_8[205]}
   );
   gpc606_5 gpc406 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[62],stage1_10[97],stage1_9[151],stage1_8[206]}
   );
   gpc606_5 gpc407 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[63],stage1_10[98],stage1_9[152],stage1_8[207]}
   );
   gpc606_5 gpc408 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[64],stage1_10[99],stage1_9[153],stage1_8[208]}
   );
   gpc606_5 gpc409 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[65],stage1_10[100],stage1_9[154],stage1_8[209]}
   );
   gpc606_5 gpc410 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[66],stage1_10[101],stage1_9[155],stage1_8[210]}
   );
   gpc606_5 gpc411 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[67],stage1_10[102],stage1_9[156],stage1_8[211]}
   );
   gpc606_5 gpc412 (
      {stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480], stage0_8[481]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[68],stage1_10[103],stage1_9[157],stage1_8[212]}
   );
   gpc606_5 gpc413 (
      {stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486], stage0_8[487]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[69],stage1_10[104],stage1_9[158],stage1_8[213]}
   );
   gpc606_5 gpc414 (
      {stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492], stage0_8[493]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[70],stage1_10[105],stage1_9[159],stage1_8[214]}
   );
   gpc606_5 gpc415 (
      {stage0_8[494], stage0_8[495], stage0_8[496], stage0_8[497], stage0_8[498], stage0_8[499]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[71],stage1_10[106],stage1_9[160],stage1_8[215]}
   );
   gpc606_5 gpc416 (
      {stage0_8[500], stage0_8[501], stage0_8[502], stage0_8[503], stage0_8[504], stage0_8[505]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[72],stage1_10[107],stage1_9[161],stage1_8[216]}
   );
   gpc606_5 gpc417 (
      {stage0_8[506], stage0_8[507], stage0_8[508], stage0_8[509], stage0_8[510], stage0_8[511]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[73],stage1_10[108],stage1_9[162],stage1_8[217]}
   );
   gpc606_5 gpc418 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[49],stage1_11[74],stage1_10[109],stage1_9[163]}
   );
   gpc615_5 gpc419 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[294]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[50],stage1_11[75],stage1_10[110],stage1_9[164]}
   );
   gpc615_5 gpc420 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[295]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[51],stage1_11[76],stage1_10[111],stage1_9[165]}
   );
   gpc615_5 gpc421 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[296]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[52],stage1_11[77],stage1_10[112],stage1_9[166]}
   );
   gpc615_5 gpc422 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[297]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[53],stage1_11[78],stage1_10[113],stage1_9[167]}
   );
   gpc615_5 gpc423 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[298]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[54],stage1_11[79],stage1_10[114],stage1_9[168]}
   );
   gpc615_5 gpc424 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[299]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[55],stage1_11[80],stage1_10[115],stage1_9[169]}
   );
   gpc615_5 gpc425 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[300]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[56],stage1_11[81],stage1_10[116],stage1_9[170]}
   );
   gpc615_5 gpc426 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[301]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[57],stage1_11[82],stage1_10[117],stage1_9[171]}
   );
   gpc615_5 gpc427 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[302]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[58],stage1_11[83],stage1_10[118],stage1_9[172]}
   );
   gpc615_5 gpc428 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[303]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[59],stage1_11[84],stage1_10[119],stage1_9[173]}
   );
   gpc615_5 gpc429 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[304]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[60],stage1_11[85],stage1_10[120],stage1_9[174]}
   );
   gpc615_5 gpc430 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[305]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[61],stage1_11[86],stage1_10[121],stage1_9[175]}
   );
   gpc615_5 gpc431 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[306]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[62],stage1_11[87],stage1_10[122],stage1_9[176]}
   );
   gpc615_5 gpc432 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[307]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[63],stage1_11[88],stage1_10[123],stage1_9[177]}
   );
   gpc615_5 gpc433 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[308]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[64],stage1_11[89],stage1_10[124],stage1_9[178]}
   );
   gpc615_5 gpc434 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[309]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[65],stage1_11[90],stage1_10[125],stage1_9[179]}
   );
   gpc615_5 gpc435 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[310]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[66],stage1_11[91],stage1_10[126],stage1_9[180]}
   );
   gpc615_5 gpc436 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[311]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[67],stage1_11[92],stage1_10[127],stage1_9[181]}
   );
   gpc615_5 gpc437 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[312]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[68],stage1_11[93],stage1_10[128],stage1_9[182]}
   );
   gpc615_5 gpc438 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[313]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[69],stage1_11[94],stage1_10[129],stage1_9[183]}
   );
   gpc615_5 gpc439 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_10[314]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[70],stage1_11[95],stage1_10[130],stage1_9[184]}
   );
   gpc615_5 gpc440 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265]},
      {stage0_10[315]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[71],stage1_11[96],stage1_10[131],stage1_9[185]}
   );
   gpc615_5 gpc441 (
      {stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_10[316]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[72],stage1_11[97],stage1_10[132],stage1_9[186]}
   );
   gpc615_5 gpc442 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_10[317]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[73],stage1_11[98],stage1_10[133],stage1_9[187]}
   );
   gpc615_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280]},
      {stage0_10[318]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[74],stage1_11[99],stage1_10[134],stage1_9[188]}
   );
   gpc615_5 gpc444 (
      {stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_10[319]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[75],stage1_11[100],stage1_10[135],stage1_9[189]}
   );
   gpc615_5 gpc445 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_10[320]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[76],stage1_11[101],stage1_10[136],stage1_9[190]}
   );
   gpc615_5 gpc446 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295]},
      {stage0_10[321]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[77],stage1_11[102],stage1_10[137],stage1_9[191]}
   );
   gpc615_5 gpc447 (
      {stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_10[322]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[78],stage1_11[103],stage1_10[138],stage1_9[192]}
   );
   gpc615_5 gpc448 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_10[323]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[79],stage1_11[104],stage1_10[139],stage1_9[193]}
   );
   gpc615_5 gpc449 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310]},
      {stage0_10[324]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[80],stage1_11[105],stage1_10[140],stage1_9[194]}
   );
   gpc615_5 gpc450 (
      {stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_10[325]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[81],stage1_11[106],stage1_10[141],stage1_9[195]}
   );
   gpc615_5 gpc451 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_10[326]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[82],stage1_11[107],stage1_10[142],stage1_9[196]}
   );
   gpc615_5 gpc452 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325]},
      {stage0_10[327]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[83],stage1_11[108],stage1_10[143],stage1_9[197]}
   );
   gpc615_5 gpc453 (
      {stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_10[328]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[84],stage1_11[109],stage1_10[144],stage1_9[198]}
   );
   gpc615_5 gpc454 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_10[329]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[85],stage1_11[110],stage1_10[145],stage1_9[199]}
   );
   gpc615_5 gpc455 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340]},
      {stage0_10[330]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[86],stage1_11[111],stage1_10[146],stage1_9[200]}
   );
   gpc615_5 gpc456 (
      {stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_10[331]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[87],stage1_11[112],stage1_10[147],stage1_9[201]}
   );
   gpc615_5 gpc457 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_10[332]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[88],stage1_11[113],stage1_10[148],stage1_9[202]}
   );
   gpc615_5 gpc458 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355]},
      {stage0_10[333]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[89],stage1_11[114],stage1_10[149],stage1_9[203]}
   );
   gpc615_5 gpc459 (
      {stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_10[334]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[90],stage1_11[115],stage1_10[150],stage1_9[204]}
   );
   gpc615_5 gpc460 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_10[335]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[91],stage1_11[116],stage1_10[151],stage1_9[205]}
   );
   gpc615_5 gpc461 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370]},
      {stage0_10[336]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[92],stage1_11[117],stage1_10[152],stage1_9[206]}
   );
   gpc615_5 gpc462 (
      {stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_10[337]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[93],stage1_11[118],stage1_10[153],stage1_9[207]}
   );
   gpc615_5 gpc463 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_10[338]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[94],stage1_11[119],stage1_10[154],stage1_9[208]}
   );
   gpc615_5 gpc464 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385]},
      {stage0_10[339]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[95],stage1_11[120],stage1_10[155],stage1_9[209]}
   );
   gpc615_5 gpc465 (
      {stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_10[340]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[96],stage1_11[121],stage1_10[156],stage1_9[210]}
   );
   gpc615_5 gpc466 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_10[341]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[97],stage1_11[122],stage1_10[157],stage1_9[211]}
   );
   gpc615_5 gpc467 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400]},
      {stage0_10[342]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[98],stage1_11[123],stage1_10[158],stage1_9[212]}
   );
   gpc615_5 gpc468 (
      {stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_10[343]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[99],stage1_11[124],stage1_10[159],stage1_9[213]}
   );
   gpc615_5 gpc469 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410]},
      {stage0_10[344]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[100],stage1_11[125],stage1_10[160],stage1_9[214]}
   );
   gpc615_5 gpc470 (
      {stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415]},
      {stage0_10[345]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[101],stage1_11[126],stage1_10[161],stage1_9[215]}
   );
   gpc615_5 gpc471 (
      {stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_10[346]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[102],stage1_11[127],stage1_10[162],stage1_9[216]}
   );
   gpc615_5 gpc472 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[347]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[103],stage1_11[128],stage1_10[163],stage1_9[217]}
   );
   gpc615_5 gpc473 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[348]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[104],stage1_11[129],stage1_10[164],stage1_9[218]}
   );
   gpc615_5 gpc474 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[349]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[105],stage1_11[130],stage1_10[165],stage1_9[219]}
   );
   gpc615_5 gpc475 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[350]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[106],stage1_11[131],stage1_10[166],stage1_9[220]}
   );
   gpc615_5 gpc476 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[351]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[107],stage1_11[132],stage1_10[167],stage1_9[221]}
   );
   gpc615_5 gpc477 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[352]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[108],stage1_11[133],stage1_10[168],stage1_9[222]}
   );
   gpc615_5 gpc478 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[353]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[109],stage1_11[134],stage1_10[169],stage1_9[223]}
   );
   gpc615_5 gpc479 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[354]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[110],stage1_11[135],stage1_10[170],stage1_9[224]}
   );
   gpc615_5 gpc480 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[355]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[111],stage1_11[136],stage1_10[171],stage1_9[225]}
   );
   gpc615_5 gpc481 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[356]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[112],stage1_11[137],stage1_10[172],stage1_9[226]}
   );
   gpc615_5 gpc482 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[357]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[113],stage1_11[138],stage1_10[173],stage1_9[227]}
   );
   gpc606_5 gpc483 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[65],stage1_12[114],stage1_11[139],stage1_10[174]}
   );
   gpc606_5 gpc484 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[66],stage1_12[115],stage1_11[140],stage1_10[175]}
   );
   gpc606_5 gpc485 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[67],stage1_12[116],stage1_11[141],stage1_10[176]}
   );
   gpc606_5 gpc486 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[68],stage1_12[117],stage1_11[142],stage1_10[177]}
   );
   gpc606_5 gpc487 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[69],stage1_12[118],stage1_11[143],stage1_10[178]}
   );
   gpc606_5 gpc488 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[70],stage1_12[119],stage1_11[144],stage1_10[179]}
   );
   gpc615_5 gpc489 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[71],stage1_12[120],stage1_11[145],stage1_10[180]}
   );
   gpc615_5 gpc490 (
      {stage0_10[399], stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[72],stage1_12[121],stage1_11[146],stage1_10[181]}
   );
   gpc615_5 gpc491 (
      {stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[73],stage1_12[122],stage1_11[147],stage1_10[182]}
   );
   gpc615_5 gpc492 (
      {stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[74],stage1_12[123],stage1_11[148],stage1_10[183]}
   );
   gpc615_5 gpc493 (
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[75],stage1_12[124],stage1_11[149],stage1_10[184]}
   );
   gpc615_5 gpc494 (
      {stage0_10[419], stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[76],stage1_12[125],stage1_11[150],stage1_10[185]}
   );
   gpc615_5 gpc495 (
      {stage0_10[424], stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[77],stage1_12[126],stage1_11[151],stage1_10[186]}
   );
   gpc615_5 gpc496 (
      {stage0_10[429], stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[78],stage1_12[127],stage1_11[152],stage1_10[187]}
   );
   gpc615_5 gpc497 (
      {stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[79],stage1_12[128],stage1_11[153],stage1_10[188]}
   );
   gpc615_5 gpc498 (
      {stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[80],stage1_12[129],stage1_11[154],stage1_10[189]}
   );
   gpc615_5 gpc499 (
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448]},
      {stage0_11[400]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[81],stage1_12[130],stage1_11[155],stage1_10[190]}
   );
   gpc615_5 gpc500 (
      {stage0_10[449], stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453]},
      {stage0_11[401]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[82],stage1_12[131],stage1_11[156],stage1_10[191]}
   );
   gpc615_5 gpc501 (
      {stage0_10[454], stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458]},
      {stage0_11[402]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[83],stage1_12[132],stage1_11[157],stage1_10[192]}
   );
   gpc615_5 gpc502 (
      {stage0_10[459], stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463]},
      {stage0_11[403]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[84],stage1_12[133],stage1_11[158],stage1_10[193]}
   );
   gpc615_5 gpc503 (
      {stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468]},
      {stage0_11[404]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[85],stage1_12[134],stage1_11[159],stage1_10[194]}
   );
   gpc615_5 gpc504 (
      {stage0_10[469], stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473]},
      {stage0_11[405]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[86],stage1_12[135],stage1_11[160],stage1_10[195]}
   );
   gpc615_5 gpc505 (
      {stage0_10[474], stage0_10[475], stage0_10[476], stage0_10[477], stage0_10[478]},
      {stage0_11[406]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[87],stage1_12[136],stage1_11[161],stage1_10[196]}
   );
   gpc615_5 gpc506 (
      {stage0_10[479], stage0_10[480], stage0_10[481], stage0_10[482], stage0_10[483]},
      {stage0_11[407]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[88],stage1_12[137],stage1_11[162],stage1_10[197]}
   );
   gpc615_5 gpc507 (
      {stage0_10[484], stage0_10[485], stage0_10[486], stage0_10[487], stage0_10[488]},
      {stage0_11[408]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[89],stage1_12[138],stage1_11[163],stage1_10[198]}
   );
   gpc615_5 gpc508 (
      {stage0_10[489], stage0_10[490], stage0_10[491], stage0_10[492], stage0_10[493]},
      {stage0_11[409]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[90],stage1_12[139],stage1_11[164],stage1_10[199]}
   );
   gpc615_5 gpc509 (
      {stage0_10[494], stage0_10[495], stage0_10[496], stage0_10[497], stage0_10[498]},
      {stage0_11[410]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[91],stage1_12[140],stage1_11[165],stage1_10[200]}
   );
   gpc615_5 gpc510 (
      {stage0_10[499], stage0_10[500], stage0_10[501], stage0_10[502], stage0_10[503]},
      {stage0_11[411]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[92],stage1_12[141],stage1_11[166],stage1_10[201]}
   );
   gpc606_5 gpc511 (
      {stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[28],stage1_13[93],stage1_12[142],stage1_11[167]}
   );
   gpc606_5 gpc512 (
      {stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[29],stage1_13[94],stage1_12[143],stage1_11[168]}
   );
   gpc606_5 gpc513 (
      {stage0_11[424], stage0_11[425], stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[30],stage1_13[95],stage1_12[144],stage1_11[169]}
   );
   gpc606_5 gpc514 (
      {stage0_11[430], stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[31],stage1_13[96],stage1_12[145],stage1_11[170]}
   );
   gpc606_5 gpc515 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[32],stage1_13[97],stage1_12[146],stage1_11[171]}
   );
   gpc606_5 gpc516 (
      {stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[33],stage1_13[98],stage1_12[147],stage1_11[172]}
   );
   gpc606_5 gpc517 (
      {stage0_11[448], stage0_11[449], stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[34],stage1_13[99],stage1_12[148],stage1_11[173]}
   );
   gpc606_5 gpc518 (
      {stage0_11[454], stage0_11[455], stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[35],stage1_13[100],stage1_12[149],stage1_11[174]}
   );
   gpc606_5 gpc519 (
      {stage0_11[460], stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[36],stage1_13[101],stage1_12[150],stage1_11[175]}
   );
   gpc615_5 gpc520 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[168]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[37],stage1_13[102],stage1_12[151],stage1_11[176]}
   );
   gpc615_5 gpc521 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[169]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[38],stage1_13[103],stage1_12[152],stage1_11[177]}
   );
   gpc615_5 gpc522 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[170]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[39],stage1_13[104],stage1_12[153],stage1_11[178]}
   );
   gpc615_5 gpc523 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[171]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[40],stage1_13[105],stage1_12[154],stage1_11[179]}
   );
   gpc615_5 gpc524 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[172]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[41],stage1_13[106],stage1_12[155],stage1_11[180]}
   );
   gpc615_5 gpc525 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[173]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[42],stage1_13[107],stage1_12[156],stage1_11[181]}
   );
   gpc615_5 gpc526 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[174]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[43],stage1_13[108],stage1_12[157],stage1_11[182]}
   );
   gpc615_5 gpc527 (
      {stage0_11[501], stage0_11[502], stage0_11[503], stage0_11[504], stage0_11[505]},
      {stage0_12[175]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[44],stage1_13[109],stage1_12[158],stage1_11[183]}
   );
   gpc606_5 gpc528 (
      {stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[17],stage1_14[45],stage1_13[110],stage1_12[159]}
   );
   gpc606_5 gpc529 (
      {stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[18],stage1_14[46],stage1_13[111],stage1_12[160]}
   );
   gpc606_5 gpc530 (
      {stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[19],stage1_14[47],stage1_13[112],stage1_12[161]}
   );
   gpc606_5 gpc531 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[20],stage1_14[48],stage1_13[113],stage1_12[162]}
   );
   gpc606_5 gpc532 (
      {stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[21],stage1_14[49],stage1_13[114],stage1_12[163]}
   );
   gpc606_5 gpc533 (
      {stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[22],stage1_14[50],stage1_13[115],stage1_12[164]}
   );
   gpc606_5 gpc534 (
      {stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[23],stage1_14[51],stage1_13[116],stage1_12[165]}
   );
   gpc606_5 gpc535 (
      {stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[24],stage1_14[52],stage1_13[117],stage1_12[166]}
   );
   gpc606_5 gpc536 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[25],stage1_14[53],stage1_13[118],stage1_12[167]}
   );
   gpc606_5 gpc537 (
      {stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[26],stage1_14[54],stage1_13[119],stage1_12[168]}
   );
   gpc606_5 gpc538 (
      {stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[27],stage1_14[55],stage1_13[120],stage1_12[169]}
   );
   gpc606_5 gpc539 (
      {stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[28],stage1_14[56],stage1_13[121],stage1_12[170]}
   );
   gpc606_5 gpc540 (
      {stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[29],stage1_14[57],stage1_13[122],stage1_12[171]}
   );
   gpc606_5 gpc541 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[30],stage1_14[58],stage1_13[123],stage1_12[172]}
   );
   gpc606_5 gpc542 (
      {stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[31],stage1_14[59],stage1_13[124],stage1_12[173]}
   );
   gpc606_5 gpc543 (
      {stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[32],stage1_14[60],stage1_13[125],stage1_12[174]}
   );
   gpc606_5 gpc544 (
      {stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[33],stage1_14[61],stage1_13[126],stage1_12[175]}
   );
   gpc606_5 gpc545 (
      {stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[34],stage1_14[62],stage1_13[127],stage1_12[176]}
   );
   gpc606_5 gpc546 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[35],stage1_14[63],stage1_13[128],stage1_12[177]}
   );
   gpc606_5 gpc547 (
      {stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[36],stage1_14[64],stage1_13[129],stage1_12[178]}
   );
   gpc606_5 gpc548 (
      {stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[37],stage1_14[65],stage1_13[130],stage1_12[179]}
   );
   gpc615_5 gpc549 (
      {stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306]},
      {stage0_13[102]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[38],stage1_14[66],stage1_13[131],stage1_12[180]}
   );
   gpc615_5 gpc550 (
      {stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_13[103]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[39],stage1_14[67],stage1_13[132],stage1_12[181]}
   );
   gpc615_5 gpc551 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_13[104]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[40],stage1_14[68],stage1_13[133],stage1_12[182]}
   );
   gpc615_5 gpc552 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[105]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[41],stage1_14[69],stage1_13[134],stage1_12[183]}
   );
   gpc615_5 gpc553 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[106]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[42],stage1_14[70],stage1_13[135],stage1_12[184]}
   );
   gpc615_5 gpc554 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[107]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[43],stage1_14[71],stage1_13[136],stage1_12[185]}
   );
   gpc615_5 gpc555 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[108]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[44],stage1_14[72],stage1_13[137],stage1_12[186]}
   );
   gpc615_5 gpc556 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[109]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[45],stage1_14[73],stage1_13[138],stage1_12[187]}
   );
   gpc615_5 gpc557 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[110]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[46],stage1_14[74],stage1_13[139],stage1_12[188]}
   );
   gpc615_5 gpc558 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[111]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[47],stage1_14[75],stage1_13[140],stage1_12[189]}
   );
   gpc615_5 gpc559 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[112]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[48],stage1_14[76],stage1_13[141],stage1_12[190]}
   );
   gpc615_5 gpc560 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[113]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[49],stage1_14[77],stage1_13[142],stage1_12[191]}
   );
   gpc615_5 gpc561 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[114]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[50],stage1_14[78],stage1_13[143],stage1_12[192]}
   );
   gpc615_5 gpc562 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[115]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[51],stage1_14[79],stage1_13[144],stage1_12[193]}
   );
   gpc615_5 gpc563 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[116]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[52],stage1_14[80],stage1_13[145],stage1_12[194]}
   );
   gpc615_5 gpc564 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[117]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[53],stage1_14[81],stage1_13[146],stage1_12[195]}
   );
   gpc615_5 gpc565 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[118]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[54],stage1_14[82],stage1_13[147],stage1_12[196]}
   );
   gpc615_5 gpc566 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[119]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[55],stage1_14[83],stage1_13[148],stage1_12[197]}
   );
   gpc615_5 gpc567 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[120]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[56],stage1_14[84],stage1_13[149],stage1_12[198]}
   );
   gpc615_5 gpc568 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[121]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[57],stage1_14[85],stage1_13[150],stage1_12[199]}
   );
   gpc615_5 gpc569 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[122]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[58],stage1_14[86],stage1_13[151],stage1_12[200]}
   );
   gpc615_5 gpc570 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[123]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[59],stage1_14[87],stage1_13[152],stage1_12[201]}
   );
   gpc615_5 gpc571 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[124]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[60],stage1_14[88],stage1_13[153],stage1_12[202]}
   );
   gpc615_5 gpc572 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[125]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[61],stage1_14[89],stage1_13[154],stage1_12[203]}
   );
   gpc615_5 gpc573 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[126]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[62],stage1_14[90],stage1_13[155],stage1_12[204]}
   );
   gpc615_5 gpc574 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[127]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[63],stage1_14[91],stage1_13[156],stage1_12[205]}
   );
   gpc615_5 gpc575 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[128]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[64],stage1_14[92],stage1_13[157],stage1_12[206]}
   );
   gpc615_5 gpc576 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[129]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[65],stage1_14[93],stage1_13[158],stage1_12[207]}
   );
   gpc615_5 gpc577 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[130]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[66],stage1_14[94],stage1_13[159],stage1_12[208]}
   );
   gpc615_5 gpc578 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[131]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[67],stage1_14[95],stage1_13[160],stage1_12[209]}
   );
   gpc615_5 gpc579 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[132]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[68],stage1_14[96],stage1_13[161],stage1_12[210]}
   );
   gpc615_5 gpc580 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[133]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[69],stage1_14[97],stage1_13[162],stage1_12[211]}
   );
   gpc615_5 gpc581 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[134]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[70],stage1_14[98],stage1_13[163],stage1_12[212]}
   );
   gpc615_5 gpc582 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[135]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[71],stage1_14[99],stage1_13[164],stage1_12[213]}
   );
   gpc615_5 gpc583 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[136]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[72],stage1_14[100],stage1_13[165],stage1_12[214]}
   );
   gpc615_5 gpc584 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[137]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[73],stage1_14[101],stage1_13[166],stage1_12[215]}
   );
   gpc615_5 gpc585 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[138]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[74],stage1_14[102],stage1_13[167],stage1_12[216]}
   );
   gpc615_5 gpc586 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[139]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[75],stage1_14[103],stage1_13[168],stage1_12[217]}
   );
   gpc615_5 gpc587 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[140]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[76],stage1_14[104],stage1_13[169],stage1_12[218]}
   );
   gpc615_5 gpc588 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[141]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[77],stage1_14[105],stage1_13[170],stage1_12[219]}
   );
   gpc615_5 gpc589 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[142]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[78],stage1_14[106],stage1_13[171],stage1_12[220]}
   );
   gpc615_5 gpc590 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[143]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[79],stage1_14[107],stage1_13[172],stage1_12[221]}
   );
   gpc606_5 gpc591 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[63],stage1_15[80],stage1_14[108],stage1_13[173]}
   );
   gpc606_5 gpc592 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[64],stage1_15[81],stage1_14[109],stage1_13[174]}
   );
   gpc606_5 gpc593 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[65],stage1_15[82],stage1_14[110],stage1_13[175]}
   );
   gpc615_5 gpc594 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166]},
      {stage0_14[378]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[66],stage1_15[83],stage1_14[111],stage1_13[176]}
   );
   gpc615_5 gpc595 (
      {stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_14[379]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[67],stage1_15[84],stage1_14[112],stage1_13[177]}
   );
   gpc615_5 gpc596 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_14[380]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[68],stage1_15[85],stage1_14[113],stage1_13[178]}
   );
   gpc615_5 gpc597 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181]},
      {stage0_14[381]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[69],stage1_15[86],stage1_14[114],stage1_13[179]}
   );
   gpc615_5 gpc598 (
      {stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186]},
      {stage0_14[382]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[70],stage1_15[87],stage1_14[115],stage1_13[180]}
   );
   gpc615_5 gpc599 (
      {stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_14[383]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[71],stage1_15[88],stage1_14[116],stage1_13[181]}
   );
   gpc615_5 gpc600 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196]},
      {stage0_14[384]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[72],stage1_15[89],stage1_14[117],stage1_13[182]}
   );
   gpc615_5 gpc601 (
      {stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_14[385]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[73],stage1_15[90],stage1_14[118],stage1_13[183]}
   );
   gpc615_5 gpc602 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_14[386]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[74],stage1_15[91],stage1_14[119],stage1_13[184]}
   );
   gpc615_5 gpc603 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211]},
      {stage0_14[387]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[75],stage1_15[92],stage1_14[120],stage1_13[185]}
   );
   gpc615_5 gpc604 (
      {stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216]},
      {stage0_14[388]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[76],stage1_15[93],stage1_14[121],stage1_13[186]}
   );
   gpc615_5 gpc605 (
      {stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_14[389]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[77],stage1_15[94],stage1_14[122],stage1_13[187]}
   );
   gpc615_5 gpc606 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226]},
      {stage0_14[390]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[78],stage1_15[95],stage1_14[123],stage1_13[188]}
   );
   gpc615_5 gpc607 (
      {stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231]},
      {stage0_14[391]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[79],stage1_15[96],stage1_14[124],stage1_13[189]}
   );
   gpc615_5 gpc608 (
      {stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_14[392]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[80],stage1_15[97],stage1_14[125],stage1_13[190]}
   );
   gpc615_5 gpc609 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241]},
      {stage0_14[393]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[81],stage1_15[98],stage1_14[126],stage1_13[191]}
   );
   gpc615_5 gpc610 (
      {stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246]},
      {stage0_14[394]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[82],stage1_15[99],stage1_14[127],stage1_13[192]}
   );
   gpc615_5 gpc611 (
      {stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_14[395]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[83],stage1_15[100],stage1_14[128],stage1_13[193]}
   );
   gpc615_5 gpc612 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256]},
      {stage0_14[396]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[84],stage1_15[101],stage1_14[129],stage1_13[194]}
   );
   gpc615_5 gpc613 (
      {stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261]},
      {stage0_14[397]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[85],stage1_15[102],stage1_14[130],stage1_13[195]}
   );
   gpc615_5 gpc614 (
      {stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_14[398]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[86],stage1_15[103],stage1_14[131],stage1_13[196]}
   );
   gpc615_5 gpc615 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271]},
      {stage0_14[399]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[87],stage1_15[104],stage1_14[132],stage1_13[197]}
   );
   gpc615_5 gpc616 (
      {stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276]},
      {stage0_14[400]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[88],stage1_15[105],stage1_14[133],stage1_13[198]}
   );
   gpc615_5 gpc617 (
      {stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_14[401]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[89],stage1_15[106],stage1_14[134],stage1_13[199]}
   );
   gpc615_5 gpc618 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286]},
      {stage0_14[402]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[90],stage1_15[107],stage1_14[135],stage1_13[200]}
   );
   gpc615_5 gpc619 (
      {stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291]},
      {stage0_14[403]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[91],stage1_15[108],stage1_14[136],stage1_13[201]}
   );
   gpc615_5 gpc620 (
      {stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_14[404]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[92],stage1_15[109],stage1_14[137],stage1_13[202]}
   );
   gpc615_5 gpc621 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301]},
      {stage0_14[405]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[93],stage1_15[110],stage1_14[138],stage1_13[203]}
   );
   gpc615_5 gpc622 (
      {stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306]},
      {stage0_14[406]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[94],stage1_15[111],stage1_14[139],stage1_13[204]}
   );
   gpc615_5 gpc623 (
      {stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_14[407]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[95],stage1_15[112],stage1_14[140],stage1_13[205]}
   );
   gpc615_5 gpc624 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316]},
      {stage0_14[408]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[96],stage1_15[113],stage1_14[141],stage1_13[206]}
   );
   gpc615_5 gpc625 (
      {stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321]},
      {stage0_14[409]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[97],stage1_15[114],stage1_14[142],stage1_13[207]}
   );
   gpc615_5 gpc626 (
      {stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_14[410]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[98],stage1_15[115],stage1_14[143],stage1_13[208]}
   );
   gpc615_5 gpc627 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331]},
      {stage0_14[411]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[99],stage1_15[116],stage1_14[144],stage1_13[209]}
   );
   gpc615_5 gpc628 (
      {stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336]},
      {stage0_14[412]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[100],stage1_15[117],stage1_14[145],stage1_13[210]}
   );
   gpc615_5 gpc629 (
      {stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_14[413]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[101],stage1_15[118],stage1_14[146],stage1_13[211]}
   );
   gpc615_5 gpc630 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346]},
      {stage0_14[414]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[102],stage1_15[119],stage1_14[147],stage1_13[212]}
   );
   gpc615_5 gpc631 (
      {stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351]},
      {stage0_14[415]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[103],stage1_15[120],stage1_14[148],stage1_13[213]}
   );
   gpc615_5 gpc632 (
      {stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_14[416]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[104],stage1_15[121],stage1_14[149],stage1_13[214]}
   );
   gpc615_5 gpc633 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361]},
      {stage0_14[417]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[105],stage1_15[122],stage1_14[150],stage1_13[215]}
   );
   gpc615_5 gpc634 (
      {stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366]},
      {stage0_14[418]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[106],stage1_15[123],stage1_14[151],stage1_13[216]}
   );
   gpc615_5 gpc635 (
      {stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_14[419]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[107],stage1_15[124],stage1_14[152],stage1_13[217]}
   );
   gpc615_5 gpc636 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376]},
      {stage0_14[420]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[108],stage1_15[125],stage1_14[153],stage1_13[218]}
   );
   gpc615_5 gpc637 (
      {stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381]},
      {stage0_14[421]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[109],stage1_15[126],stage1_14[154],stage1_13[219]}
   );
   gpc615_5 gpc638 (
      {stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_14[422]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[110],stage1_15[127],stage1_14[155],stage1_13[220]}
   );
   gpc615_5 gpc639 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391]},
      {stage0_14[423]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[111],stage1_15[128],stage1_14[156],stage1_13[221]}
   );
   gpc615_5 gpc640 (
      {stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396]},
      {stage0_14[424]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[112],stage1_15[129],stage1_14[157],stage1_13[222]}
   );
   gpc615_5 gpc641 (
      {stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_14[425]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[113],stage1_15[130],stage1_14[158],stage1_13[223]}
   );
   gpc615_5 gpc642 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406]},
      {stage0_14[426]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[114],stage1_15[131],stage1_14[159],stage1_13[224]}
   );
   gpc615_5 gpc643 (
      {stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411]},
      {stage0_14[427]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[115],stage1_15[132],stage1_14[160],stage1_13[225]}
   );
   gpc615_5 gpc644 (
      {stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_14[428]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[116],stage1_15[133],stage1_14[161],stage1_13[226]}
   );
   gpc615_5 gpc645 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421]},
      {stage0_14[429]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[117],stage1_15[134],stage1_14[162],stage1_13[227]}
   );
   gpc615_5 gpc646 (
      {stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426]},
      {stage0_14[430]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[118],stage1_15[135],stage1_14[163],stage1_13[228]}
   );
   gpc615_5 gpc647 (
      {stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_14[431]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[119],stage1_15[136],stage1_14[164],stage1_13[229]}
   );
   gpc615_5 gpc648 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436]},
      {stage0_14[432]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[120],stage1_15[137],stage1_14[165],stage1_13[230]}
   );
   gpc615_5 gpc649 (
      {stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441]},
      {stage0_14[433]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[121],stage1_15[138],stage1_14[166],stage1_13[231]}
   );
   gpc615_5 gpc650 (
      {stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_14[434]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[122],stage1_15[139],stage1_14[167],stage1_13[232]}
   );
   gpc615_5 gpc651 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451]},
      {stage0_14[435]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[123],stage1_15[140],stage1_14[168],stage1_13[233]}
   );
   gpc615_5 gpc652 (
      {stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456]},
      {stage0_14[436]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[124],stage1_15[141],stage1_14[169],stage1_13[234]}
   );
   gpc615_5 gpc653 (
      {stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_14[437]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[125],stage1_15[142],stage1_14[170],stage1_13[235]}
   );
   gpc615_5 gpc654 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466]},
      {stage0_14[438]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[126],stage1_15[143],stage1_14[171],stage1_13[236]}
   );
   gpc1_1 gpc655 (
      {stage0_0[509]},
      {stage1_0[98]}
   );
   gpc1_1 gpc656 (
      {stage0_0[510]},
      {stage1_0[99]}
   );
   gpc1_1 gpc657 (
      {stage0_0[511]},
      {stage1_0[100]}
   );
   gpc1_1 gpc658 (
      {stage0_1[476]},
      {stage1_1[144]}
   );
   gpc1_1 gpc659 (
      {stage0_1[477]},
      {stage1_1[145]}
   );
   gpc1_1 gpc660 (
      {stage0_1[478]},
      {stage1_1[146]}
   );
   gpc1_1 gpc661 (
      {stage0_1[479]},
      {stage1_1[147]}
   );
   gpc1_1 gpc662 (
      {stage0_1[480]},
      {stage1_1[148]}
   );
   gpc1_1 gpc663 (
      {stage0_1[481]},
      {stage1_1[149]}
   );
   gpc1_1 gpc664 (
      {stage0_1[482]},
      {stage1_1[150]}
   );
   gpc1_1 gpc665 (
      {stage0_1[483]},
      {stage1_1[151]}
   );
   gpc1_1 gpc666 (
      {stage0_1[484]},
      {stage1_1[152]}
   );
   gpc1_1 gpc667 (
      {stage0_1[485]},
      {stage1_1[153]}
   );
   gpc1_1 gpc668 (
      {stage0_1[486]},
      {stage1_1[154]}
   );
   gpc1_1 gpc669 (
      {stage0_1[487]},
      {stage1_1[155]}
   );
   gpc1_1 gpc670 (
      {stage0_1[488]},
      {stage1_1[156]}
   );
   gpc1_1 gpc671 (
      {stage0_1[489]},
      {stage1_1[157]}
   );
   gpc1_1 gpc672 (
      {stage0_1[490]},
      {stage1_1[158]}
   );
   gpc1_1 gpc673 (
      {stage0_1[491]},
      {stage1_1[159]}
   );
   gpc1_1 gpc674 (
      {stage0_1[492]},
      {stage1_1[160]}
   );
   gpc1_1 gpc675 (
      {stage0_1[493]},
      {stage1_1[161]}
   );
   gpc1_1 gpc676 (
      {stage0_1[494]},
      {stage1_1[162]}
   );
   gpc1_1 gpc677 (
      {stage0_1[495]},
      {stage1_1[163]}
   );
   gpc1_1 gpc678 (
      {stage0_1[496]},
      {stage1_1[164]}
   );
   gpc1_1 gpc679 (
      {stage0_1[497]},
      {stage1_1[165]}
   );
   gpc1_1 gpc680 (
      {stage0_1[498]},
      {stage1_1[166]}
   );
   gpc1_1 gpc681 (
      {stage0_1[499]},
      {stage1_1[167]}
   );
   gpc1_1 gpc682 (
      {stage0_1[500]},
      {stage1_1[168]}
   );
   gpc1_1 gpc683 (
      {stage0_1[501]},
      {stage1_1[169]}
   );
   gpc1_1 gpc684 (
      {stage0_1[502]},
      {stage1_1[170]}
   );
   gpc1_1 gpc685 (
      {stage0_1[503]},
      {stage1_1[171]}
   );
   gpc1_1 gpc686 (
      {stage0_1[504]},
      {stage1_1[172]}
   );
   gpc1_1 gpc687 (
      {stage0_1[505]},
      {stage1_1[173]}
   );
   gpc1_1 gpc688 (
      {stage0_1[506]},
      {stage1_1[174]}
   );
   gpc1_1 gpc689 (
      {stage0_1[507]},
      {stage1_1[175]}
   );
   gpc1_1 gpc690 (
      {stage0_1[508]},
      {stage1_1[176]}
   );
   gpc1_1 gpc691 (
      {stage0_1[509]},
      {stage1_1[177]}
   );
   gpc1_1 gpc692 (
      {stage0_1[510]},
      {stage1_1[178]}
   );
   gpc1_1 gpc693 (
      {stage0_1[511]},
      {stage1_1[179]}
   );
   gpc1_1 gpc694 (
      {stage0_3[466]},
      {stage1_3[200]}
   );
   gpc1_1 gpc695 (
      {stage0_3[467]},
      {stage1_3[201]}
   );
   gpc1_1 gpc696 (
      {stage0_3[468]},
      {stage1_3[202]}
   );
   gpc1_1 gpc697 (
      {stage0_3[469]},
      {stage1_3[203]}
   );
   gpc1_1 gpc698 (
      {stage0_3[470]},
      {stage1_3[204]}
   );
   gpc1_1 gpc699 (
      {stage0_3[471]},
      {stage1_3[205]}
   );
   gpc1_1 gpc700 (
      {stage0_3[472]},
      {stage1_3[206]}
   );
   gpc1_1 gpc701 (
      {stage0_3[473]},
      {stage1_3[207]}
   );
   gpc1_1 gpc702 (
      {stage0_3[474]},
      {stage1_3[208]}
   );
   gpc1_1 gpc703 (
      {stage0_3[475]},
      {stage1_3[209]}
   );
   gpc1_1 gpc704 (
      {stage0_3[476]},
      {stage1_3[210]}
   );
   gpc1_1 gpc705 (
      {stage0_3[477]},
      {stage1_3[211]}
   );
   gpc1_1 gpc706 (
      {stage0_3[478]},
      {stage1_3[212]}
   );
   gpc1_1 gpc707 (
      {stage0_3[479]},
      {stage1_3[213]}
   );
   gpc1_1 gpc708 (
      {stage0_3[480]},
      {stage1_3[214]}
   );
   gpc1_1 gpc709 (
      {stage0_3[481]},
      {stage1_3[215]}
   );
   gpc1_1 gpc710 (
      {stage0_3[482]},
      {stage1_3[216]}
   );
   gpc1_1 gpc711 (
      {stage0_3[483]},
      {stage1_3[217]}
   );
   gpc1_1 gpc712 (
      {stage0_3[484]},
      {stage1_3[218]}
   );
   gpc1_1 gpc713 (
      {stage0_3[485]},
      {stage1_3[219]}
   );
   gpc1_1 gpc714 (
      {stage0_3[486]},
      {stage1_3[220]}
   );
   gpc1_1 gpc715 (
      {stage0_3[487]},
      {stage1_3[221]}
   );
   gpc1_1 gpc716 (
      {stage0_3[488]},
      {stage1_3[222]}
   );
   gpc1_1 gpc717 (
      {stage0_3[489]},
      {stage1_3[223]}
   );
   gpc1_1 gpc718 (
      {stage0_3[490]},
      {stage1_3[224]}
   );
   gpc1_1 gpc719 (
      {stage0_3[491]},
      {stage1_3[225]}
   );
   gpc1_1 gpc720 (
      {stage0_3[492]},
      {stage1_3[226]}
   );
   gpc1_1 gpc721 (
      {stage0_3[493]},
      {stage1_3[227]}
   );
   gpc1_1 gpc722 (
      {stage0_3[494]},
      {stage1_3[228]}
   );
   gpc1_1 gpc723 (
      {stage0_3[495]},
      {stage1_3[229]}
   );
   gpc1_1 gpc724 (
      {stage0_3[496]},
      {stage1_3[230]}
   );
   gpc1_1 gpc725 (
      {stage0_3[497]},
      {stage1_3[231]}
   );
   gpc1_1 gpc726 (
      {stage0_3[498]},
      {stage1_3[232]}
   );
   gpc1_1 gpc727 (
      {stage0_3[499]},
      {stage1_3[233]}
   );
   gpc1_1 gpc728 (
      {stage0_3[500]},
      {stage1_3[234]}
   );
   gpc1_1 gpc729 (
      {stage0_3[501]},
      {stage1_3[235]}
   );
   gpc1_1 gpc730 (
      {stage0_3[502]},
      {stage1_3[236]}
   );
   gpc1_1 gpc731 (
      {stage0_3[503]},
      {stage1_3[237]}
   );
   gpc1_1 gpc732 (
      {stage0_3[504]},
      {stage1_3[238]}
   );
   gpc1_1 gpc733 (
      {stage0_3[505]},
      {stage1_3[239]}
   );
   gpc1_1 gpc734 (
      {stage0_3[506]},
      {stage1_3[240]}
   );
   gpc1_1 gpc735 (
      {stage0_3[507]},
      {stage1_3[241]}
   );
   gpc1_1 gpc736 (
      {stage0_3[508]},
      {stage1_3[242]}
   );
   gpc1_1 gpc737 (
      {stage0_3[509]},
      {stage1_3[243]}
   );
   gpc1_1 gpc738 (
      {stage0_3[510]},
      {stage1_3[244]}
   );
   gpc1_1 gpc739 (
      {stage0_3[511]},
      {stage1_3[245]}
   );
   gpc1_1 gpc740 (
      {stage0_5[505]},
      {stage1_5[211]}
   );
   gpc1_1 gpc741 (
      {stage0_5[506]},
      {stage1_5[212]}
   );
   gpc1_1 gpc742 (
      {stage0_5[507]},
      {stage1_5[213]}
   );
   gpc1_1 gpc743 (
      {stage0_5[508]},
      {stage1_5[214]}
   );
   gpc1_1 gpc744 (
      {stage0_5[509]},
      {stage1_5[215]}
   );
   gpc1_1 gpc745 (
      {stage0_5[510]},
      {stage1_5[216]}
   );
   gpc1_1 gpc746 (
      {stage0_5[511]},
      {stage1_5[217]}
   );
   gpc1_1 gpc747 (
      {stage0_6[505]},
      {stage1_6[200]}
   );
   gpc1_1 gpc748 (
      {stage0_6[506]},
      {stage1_6[201]}
   );
   gpc1_1 gpc749 (
      {stage0_6[507]},
      {stage1_6[202]}
   );
   gpc1_1 gpc750 (
      {stage0_6[508]},
      {stage1_6[203]}
   );
   gpc1_1 gpc751 (
      {stage0_6[509]},
      {stage1_6[204]}
   );
   gpc1_1 gpc752 (
      {stage0_6[510]},
      {stage1_6[205]}
   );
   gpc1_1 gpc753 (
      {stage0_6[511]},
      {stage1_6[206]}
   );
   gpc1_1 gpc754 (
      {stage0_7[501]},
      {stage1_7[196]}
   );
   gpc1_1 gpc755 (
      {stage0_7[502]},
      {stage1_7[197]}
   );
   gpc1_1 gpc756 (
      {stage0_7[503]},
      {stage1_7[198]}
   );
   gpc1_1 gpc757 (
      {stage0_7[504]},
      {stage1_7[199]}
   );
   gpc1_1 gpc758 (
      {stage0_7[505]},
      {stage1_7[200]}
   );
   gpc1_1 gpc759 (
      {stage0_7[506]},
      {stage1_7[201]}
   );
   gpc1_1 gpc760 (
      {stage0_7[507]},
      {stage1_7[202]}
   );
   gpc1_1 gpc761 (
      {stage0_7[508]},
      {stage1_7[203]}
   );
   gpc1_1 gpc762 (
      {stage0_7[509]},
      {stage1_7[204]}
   );
   gpc1_1 gpc763 (
      {stage0_7[510]},
      {stage1_7[205]}
   );
   gpc1_1 gpc764 (
      {stage0_7[511]},
      {stage1_7[206]}
   );
   gpc1_1 gpc765 (
      {stage0_9[476]},
      {stage1_9[228]}
   );
   gpc1_1 gpc766 (
      {stage0_9[477]},
      {stage1_9[229]}
   );
   gpc1_1 gpc767 (
      {stage0_9[478]},
      {stage1_9[230]}
   );
   gpc1_1 gpc768 (
      {stage0_9[479]},
      {stage1_9[231]}
   );
   gpc1_1 gpc769 (
      {stage0_9[480]},
      {stage1_9[232]}
   );
   gpc1_1 gpc770 (
      {stage0_9[481]},
      {stage1_9[233]}
   );
   gpc1_1 gpc771 (
      {stage0_9[482]},
      {stage1_9[234]}
   );
   gpc1_1 gpc772 (
      {stage0_9[483]},
      {stage1_9[235]}
   );
   gpc1_1 gpc773 (
      {stage0_9[484]},
      {stage1_9[236]}
   );
   gpc1_1 gpc774 (
      {stage0_9[485]},
      {stage1_9[237]}
   );
   gpc1_1 gpc775 (
      {stage0_9[486]},
      {stage1_9[238]}
   );
   gpc1_1 gpc776 (
      {stage0_9[487]},
      {stage1_9[239]}
   );
   gpc1_1 gpc777 (
      {stage0_9[488]},
      {stage1_9[240]}
   );
   gpc1_1 gpc778 (
      {stage0_9[489]},
      {stage1_9[241]}
   );
   gpc1_1 gpc779 (
      {stage0_9[490]},
      {stage1_9[242]}
   );
   gpc1_1 gpc780 (
      {stage0_9[491]},
      {stage1_9[243]}
   );
   gpc1_1 gpc781 (
      {stage0_9[492]},
      {stage1_9[244]}
   );
   gpc1_1 gpc782 (
      {stage0_9[493]},
      {stage1_9[245]}
   );
   gpc1_1 gpc783 (
      {stage0_9[494]},
      {stage1_9[246]}
   );
   gpc1_1 gpc784 (
      {stage0_9[495]},
      {stage1_9[247]}
   );
   gpc1_1 gpc785 (
      {stage0_9[496]},
      {stage1_9[248]}
   );
   gpc1_1 gpc786 (
      {stage0_9[497]},
      {stage1_9[249]}
   );
   gpc1_1 gpc787 (
      {stage0_9[498]},
      {stage1_9[250]}
   );
   gpc1_1 gpc788 (
      {stage0_9[499]},
      {stage1_9[251]}
   );
   gpc1_1 gpc789 (
      {stage0_9[500]},
      {stage1_9[252]}
   );
   gpc1_1 gpc790 (
      {stage0_9[501]},
      {stage1_9[253]}
   );
   gpc1_1 gpc791 (
      {stage0_9[502]},
      {stage1_9[254]}
   );
   gpc1_1 gpc792 (
      {stage0_9[503]},
      {stage1_9[255]}
   );
   gpc1_1 gpc793 (
      {stage0_9[504]},
      {stage1_9[256]}
   );
   gpc1_1 gpc794 (
      {stage0_9[505]},
      {stage1_9[257]}
   );
   gpc1_1 gpc795 (
      {stage0_9[506]},
      {stage1_9[258]}
   );
   gpc1_1 gpc796 (
      {stage0_9[507]},
      {stage1_9[259]}
   );
   gpc1_1 gpc797 (
      {stage0_9[508]},
      {stage1_9[260]}
   );
   gpc1_1 gpc798 (
      {stage0_9[509]},
      {stage1_9[261]}
   );
   gpc1_1 gpc799 (
      {stage0_9[510]},
      {stage1_9[262]}
   );
   gpc1_1 gpc800 (
      {stage0_9[511]},
      {stage1_9[263]}
   );
   gpc1_1 gpc801 (
      {stage0_10[504]},
      {stage1_10[202]}
   );
   gpc1_1 gpc802 (
      {stage0_10[505]},
      {stage1_10[203]}
   );
   gpc1_1 gpc803 (
      {stage0_10[506]},
      {stage1_10[204]}
   );
   gpc1_1 gpc804 (
      {stage0_10[507]},
      {stage1_10[205]}
   );
   gpc1_1 gpc805 (
      {stage0_10[508]},
      {stage1_10[206]}
   );
   gpc1_1 gpc806 (
      {stage0_10[509]},
      {stage1_10[207]}
   );
   gpc1_1 gpc807 (
      {stage0_10[510]},
      {stage1_10[208]}
   );
   gpc1_1 gpc808 (
      {stage0_10[511]},
      {stage1_10[209]}
   );
   gpc1_1 gpc809 (
      {stage0_11[506]},
      {stage1_11[184]}
   );
   gpc1_1 gpc810 (
      {stage0_11[507]},
      {stage1_11[185]}
   );
   gpc1_1 gpc811 (
      {stage0_11[508]},
      {stage1_11[186]}
   );
   gpc1_1 gpc812 (
      {stage0_11[509]},
      {stage1_11[187]}
   );
   gpc1_1 gpc813 (
      {stage0_11[510]},
      {stage1_11[188]}
   );
   gpc1_1 gpc814 (
      {stage0_11[511]},
      {stage1_11[189]}
   );
   gpc1_1 gpc815 (
      {stage0_13[467]},
      {stage1_13[237]}
   );
   gpc1_1 gpc816 (
      {stage0_13[468]},
      {stage1_13[238]}
   );
   gpc1_1 gpc817 (
      {stage0_13[469]},
      {stage1_13[239]}
   );
   gpc1_1 gpc818 (
      {stage0_13[470]},
      {stage1_13[240]}
   );
   gpc1_1 gpc819 (
      {stage0_13[471]},
      {stage1_13[241]}
   );
   gpc1_1 gpc820 (
      {stage0_13[472]},
      {stage1_13[242]}
   );
   gpc1_1 gpc821 (
      {stage0_13[473]},
      {stage1_13[243]}
   );
   gpc1_1 gpc822 (
      {stage0_13[474]},
      {stage1_13[244]}
   );
   gpc1_1 gpc823 (
      {stage0_13[475]},
      {stage1_13[245]}
   );
   gpc1_1 gpc824 (
      {stage0_13[476]},
      {stage1_13[246]}
   );
   gpc1_1 gpc825 (
      {stage0_13[477]},
      {stage1_13[247]}
   );
   gpc1_1 gpc826 (
      {stage0_13[478]},
      {stage1_13[248]}
   );
   gpc1_1 gpc827 (
      {stage0_13[479]},
      {stage1_13[249]}
   );
   gpc1_1 gpc828 (
      {stage0_13[480]},
      {stage1_13[250]}
   );
   gpc1_1 gpc829 (
      {stage0_13[481]},
      {stage1_13[251]}
   );
   gpc1_1 gpc830 (
      {stage0_13[482]},
      {stage1_13[252]}
   );
   gpc1_1 gpc831 (
      {stage0_13[483]},
      {stage1_13[253]}
   );
   gpc1_1 gpc832 (
      {stage0_13[484]},
      {stage1_13[254]}
   );
   gpc1_1 gpc833 (
      {stage0_13[485]},
      {stage1_13[255]}
   );
   gpc1_1 gpc834 (
      {stage0_13[486]},
      {stage1_13[256]}
   );
   gpc1_1 gpc835 (
      {stage0_13[487]},
      {stage1_13[257]}
   );
   gpc1_1 gpc836 (
      {stage0_13[488]},
      {stage1_13[258]}
   );
   gpc1_1 gpc837 (
      {stage0_13[489]},
      {stage1_13[259]}
   );
   gpc1_1 gpc838 (
      {stage0_13[490]},
      {stage1_13[260]}
   );
   gpc1_1 gpc839 (
      {stage0_13[491]},
      {stage1_13[261]}
   );
   gpc1_1 gpc840 (
      {stage0_13[492]},
      {stage1_13[262]}
   );
   gpc1_1 gpc841 (
      {stage0_13[493]},
      {stage1_13[263]}
   );
   gpc1_1 gpc842 (
      {stage0_13[494]},
      {stage1_13[264]}
   );
   gpc1_1 gpc843 (
      {stage0_13[495]},
      {stage1_13[265]}
   );
   gpc1_1 gpc844 (
      {stage0_13[496]},
      {stage1_13[266]}
   );
   gpc1_1 gpc845 (
      {stage0_13[497]},
      {stage1_13[267]}
   );
   gpc1_1 gpc846 (
      {stage0_13[498]},
      {stage1_13[268]}
   );
   gpc1_1 gpc847 (
      {stage0_13[499]},
      {stage1_13[269]}
   );
   gpc1_1 gpc848 (
      {stage0_13[500]},
      {stage1_13[270]}
   );
   gpc1_1 gpc849 (
      {stage0_13[501]},
      {stage1_13[271]}
   );
   gpc1_1 gpc850 (
      {stage0_13[502]},
      {stage1_13[272]}
   );
   gpc1_1 gpc851 (
      {stage0_13[503]},
      {stage1_13[273]}
   );
   gpc1_1 gpc852 (
      {stage0_13[504]},
      {stage1_13[274]}
   );
   gpc1_1 gpc853 (
      {stage0_13[505]},
      {stage1_13[275]}
   );
   gpc1_1 gpc854 (
      {stage0_13[506]},
      {stage1_13[276]}
   );
   gpc1_1 gpc855 (
      {stage0_13[507]},
      {stage1_13[277]}
   );
   gpc1_1 gpc856 (
      {stage0_13[508]},
      {stage1_13[278]}
   );
   gpc1_1 gpc857 (
      {stage0_13[509]},
      {stage1_13[279]}
   );
   gpc1_1 gpc858 (
      {stage0_13[510]},
      {stage1_13[280]}
   );
   gpc1_1 gpc859 (
      {stage0_13[511]},
      {stage1_13[281]}
   );
   gpc1_1 gpc860 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc861 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc862 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc863 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc864 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc865 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc866 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc867 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc868 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc869 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc870 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc871 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc872 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc873 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc874 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc875 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc876 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc877 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc878 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc879 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc880 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc881 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc882 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc883 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc884 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc885 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc886 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc887 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc888 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc889 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc890 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc891 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc892 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc893 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc894 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc895 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc896 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc897 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc898 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc899 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc900 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc901 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc902 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc903 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc904 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc905 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc906 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc907 (
      {stage0_14[486]},
      {stage1_14[219]}
   );
   gpc1_1 gpc908 (
      {stage0_14[487]},
      {stage1_14[220]}
   );
   gpc1_1 gpc909 (
      {stage0_14[488]},
      {stage1_14[221]}
   );
   gpc1_1 gpc910 (
      {stage0_14[489]},
      {stage1_14[222]}
   );
   gpc1_1 gpc911 (
      {stage0_14[490]},
      {stage1_14[223]}
   );
   gpc1_1 gpc912 (
      {stage0_14[491]},
      {stage1_14[224]}
   );
   gpc1_1 gpc913 (
      {stage0_14[492]},
      {stage1_14[225]}
   );
   gpc1_1 gpc914 (
      {stage0_14[493]},
      {stage1_14[226]}
   );
   gpc1_1 gpc915 (
      {stage0_14[494]},
      {stage1_14[227]}
   );
   gpc1_1 gpc916 (
      {stage0_14[495]},
      {stage1_14[228]}
   );
   gpc1_1 gpc917 (
      {stage0_14[496]},
      {stage1_14[229]}
   );
   gpc1_1 gpc918 (
      {stage0_14[497]},
      {stage1_14[230]}
   );
   gpc1_1 gpc919 (
      {stage0_14[498]},
      {stage1_14[231]}
   );
   gpc1_1 gpc920 (
      {stage0_14[499]},
      {stage1_14[232]}
   );
   gpc1_1 gpc921 (
      {stage0_14[500]},
      {stage1_14[233]}
   );
   gpc1_1 gpc922 (
      {stage0_14[501]},
      {stage1_14[234]}
   );
   gpc1_1 gpc923 (
      {stage0_14[502]},
      {stage1_14[235]}
   );
   gpc1_1 gpc924 (
      {stage0_14[503]},
      {stage1_14[236]}
   );
   gpc1_1 gpc925 (
      {stage0_14[504]},
      {stage1_14[237]}
   );
   gpc1_1 gpc926 (
      {stage0_14[505]},
      {stage1_14[238]}
   );
   gpc1_1 gpc927 (
      {stage0_14[506]},
      {stage1_14[239]}
   );
   gpc1_1 gpc928 (
      {stage0_14[507]},
      {stage1_14[240]}
   );
   gpc1_1 gpc929 (
      {stage0_14[508]},
      {stage1_14[241]}
   );
   gpc1_1 gpc930 (
      {stage0_14[509]},
      {stage1_14[242]}
   );
   gpc1_1 gpc931 (
      {stage0_14[510]},
      {stage1_14[243]}
   );
   gpc1_1 gpc932 (
      {stage0_14[511]},
      {stage1_14[244]}
   );
   gpc1_1 gpc933 (
      {stage0_15[384]},
      {stage1_15[144]}
   );
   gpc1_1 gpc934 (
      {stage0_15[385]},
      {stage1_15[145]}
   );
   gpc1_1 gpc935 (
      {stage0_15[386]},
      {stage1_15[146]}
   );
   gpc1_1 gpc936 (
      {stage0_15[387]},
      {stage1_15[147]}
   );
   gpc1_1 gpc937 (
      {stage0_15[388]},
      {stage1_15[148]}
   );
   gpc1_1 gpc938 (
      {stage0_15[389]},
      {stage1_15[149]}
   );
   gpc1_1 gpc939 (
      {stage0_15[390]},
      {stage1_15[150]}
   );
   gpc1_1 gpc940 (
      {stage0_15[391]},
      {stage1_15[151]}
   );
   gpc1_1 gpc941 (
      {stage0_15[392]},
      {stage1_15[152]}
   );
   gpc1_1 gpc942 (
      {stage0_15[393]},
      {stage1_15[153]}
   );
   gpc1_1 gpc943 (
      {stage0_15[394]},
      {stage1_15[154]}
   );
   gpc1_1 gpc944 (
      {stage0_15[395]},
      {stage1_15[155]}
   );
   gpc1_1 gpc945 (
      {stage0_15[396]},
      {stage1_15[156]}
   );
   gpc1_1 gpc946 (
      {stage0_15[397]},
      {stage1_15[157]}
   );
   gpc1_1 gpc947 (
      {stage0_15[398]},
      {stage1_15[158]}
   );
   gpc1_1 gpc948 (
      {stage0_15[399]},
      {stage1_15[159]}
   );
   gpc1_1 gpc949 (
      {stage0_15[400]},
      {stage1_15[160]}
   );
   gpc1_1 gpc950 (
      {stage0_15[401]},
      {stage1_15[161]}
   );
   gpc1_1 gpc951 (
      {stage0_15[402]},
      {stage1_15[162]}
   );
   gpc1_1 gpc952 (
      {stage0_15[403]},
      {stage1_15[163]}
   );
   gpc1_1 gpc953 (
      {stage0_15[404]},
      {stage1_15[164]}
   );
   gpc1_1 gpc954 (
      {stage0_15[405]},
      {stage1_15[165]}
   );
   gpc1_1 gpc955 (
      {stage0_15[406]},
      {stage1_15[166]}
   );
   gpc1_1 gpc956 (
      {stage0_15[407]},
      {stage1_15[167]}
   );
   gpc1_1 gpc957 (
      {stage0_15[408]},
      {stage1_15[168]}
   );
   gpc1_1 gpc958 (
      {stage0_15[409]},
      {stage1_15[169]}
   );
   gpc1_1 gpc959 (
      {stage0_15[410]},
      {stage1_15[170]}
   );
   gpc1_1 gpc960 (
      {stage0_15[411]},
      {stage1_15[171]}
   );
   gpc1_1 gpc961 (
      {stage0_15[412]},
      {stage1_15[172]}
   );
   gpc1_1 gpc962 (
      {stage0_15[413]},
      {stage1_15[173]}
   );
   gpc1_1 gpc963 (
      {stage0_15[414]},
      {stage1_15[174]}
   );
   gpc1_1 gpc964 (
      {stage0_15[415]},
      {stage1_15[175]}
   );
   gpc1_1 gpc965 (
      {stage0_15[416]},
      {stage1_15[176]}
   );
   gpc1_1 gpc966 (
      {stage0_15[417]},
      {stage1_15[177]}
   );
   gpc1_1 gpc967 (
      {stage0_15[418]},
      {stage1_15[178]}
   );
   gpc1_1 gpc968 (
      {stage0_15[419]},
      {stage1_15[179]}
   );
   gpc1_1 gpc969 (
      {stage0_15[420]},
      {stage1_15[180]}
   );
   gpc1_1 gpc970 (
      {stage0_15[421]},
      {stage1_15[181]}
   );
   gpc1_1 gpc971 (
      {stage0_15[422]},
      {stage1_15[182]}
   );
   gpc1_1 gpc972 (
      {stage0_15[423]},
      {stage1_15[183]}
   );
   gpc1_1 gpc973 (
      {stage0_15[424]},
      {stage1_15[184]}
   );
   gpc1_1 gpc974 (
      {stage0_15[425]},
      {stage1_15[185]}
   );
   gpc1_1 gpc975 (
      {stage0_15[426]},
      {stage1_15[186]}
   );
   gpc1_1 gpc976 (
      {stage0_15[427]},
      {stage1_15[187]}
   );
   gpc1_1 gpc977 (
      {stage0_15[428]},
      {stage1_15[188]}
   );
   gpc1_1 gpc978 (
      {stage0_15[429]},
      {stage1_15[189]}
   );
   gpc1_1 gpc979 (
      {stage0_15[430]},
      {stage1_15[190]}
   );
   gpc1_1 gpc980 (
      {stage0_15[431]},
      {stage1_15[191]}
   );
   gpc1_1 gpc981 (
      {stage0_15[432]},
      {stage1_15[192]}
   );
   gpc1_1 gpc982 (
      {stage0_15[433]},
      {stage1_15[193]}
   );
   gpc1_1 gpc983 (
      {stage0_15[434]},
      {stage1_15[194]}
   );
   gpc1_1 gpc984 (
      {stage0_15[435]},
      {stage1_15[195]}
   );
   gpc1_1 gpc985 (
      {stage0_15[436]},
      {stage1_15[196]}
   );
   gpc1_1 gpc986 (
      {stage0_15[437]},
      {stage1_15[197]}
   );
   gpc1_1 gpc987 (
      {stage0_15[438]},
      {stage1_15[198]}
   );
   gpc1_1 gpc988 (
      {stage0_15[439]},
      {stage1_15[199]}
   );
   gpc1_1 gpc989 (
      {stage0_15[440]},
      {stage1_15[200]}
   );
   gpc1_1 gpc990 (
      {stage0_15[441]},
      {stage1_15[201]}
   );
   gpc1_1 gpc991 (
      {stage0_15[442]},
      {stage1_15[202]}
   );
   gpc1_1 gpc992 (
      {stage0_15[443]},
      {stage1_15[203]}
   );
   gpc1_1 gpc993 (
      {stage0_15[444]},
      {stage1_15[204]}
   );
   gpc1_1 gpc994 (
      {stage0_15[445]},
      {stage1_15[205]}
   );
   gpc1_1 gpc995 (
      {stage0_15[446]},
      {stage1_15[206]}
   );
   gpc1_1 gpc996 (
      {stage0_15[447]},
      {stage1_15[207]}
   );
   gpc1_1 gpc997 (
      {stage0_15[448]},
      {stage1_15[208]}
   );
   gpc1_1 gpc998 (
      {stage0_15[449]},
      {stage1_15[209]}
   );
   gpc1_1 gpc999 (
      {stage0_15[450]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[451]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[452]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[453]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[454]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[455]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[456]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[457]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1007 (
      {stage0_15[458]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1008 (
      {stage0_15[459]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1009 (
      {stage0_15[460]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1010 (
      {stage0_15[461]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1011 (
      {stage0_15[462]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1012 (
      {stage0_15[463]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1013 (
      {stage0_15[464]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1014 (
      {stage0_15[465]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1015 (
      {stage0_15[466]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1016 (
      {stage0_15[467]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1017 (
      {stage0_15[468]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1018 (
      {stage0_15[469]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1019 (
      {stage0_15[470]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1020 (
      {stage0_15[471]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1021 (
      {stage0_15[472]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1022 (
      {stage0_15[473]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1023 (
      {stage0_15[474]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1024 (
      {stage0_15[475]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1025 (
      {stage0_15[476]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1026 (
      {stage0_15[477]},
      {stage1_15[237]}
   );
   gpc1_1 gpc1027 (
      {stage0_15[478]},
      {stage1_15[238]}
   );
   gpc1_1 gpc1028 (
      {stage0_15[479]},
      {stage1_15[239]}
   );
   gpc1_1 gpc1029 (
      {stage0_15[480]},
      {stage1_15[240]}
   );
   gpc1_1 gpc1030 (
      {stage0_15[481]},
      {stage1_15[241]}
   );
   gpc1_1 gpc1031 (
      {stage0_15[482]},
      {stage1_15[242]}
   );
   gpc1_1 gpc1032 (
      {stage0_15[483]},
      {stage1_15[243]}
   );
   gpc1_1 gpc1033 (
      {stage0_15[484]},
      {stage1_15[244]}
   );
   gpc1_1 gpc1034 (
      {stage0_15[485]},
      {stage1_15[245]}
   );
   gpc1_1 gpc1035 (
      {stage0_15[486]},
      {stage1_15[246]}
   );
   gpc1_1 gpc1036 (
      {stage0_15[487]},
      {stage1_15[247]}
   );
   gpc1_1 gpc1037 (
      {stage0_15[488]},
      {stage1_15[248]}
   );
   gpc1_1 gpc1038 (
      {stage0_15[489]},
      {stage1_15[249]}
   );
   gpc1_1 gpc1039 (
      {stage0_15[490]},
      {stage1_15[250]}
   );
   gpc1_1 gpc1040 (
      {stage0_15[491]},
      {stage1_15[251]}
   );
   gpc1_1 gpc1041 (
      {stage0_15[492]},
      {stage1_15[252]}
   );
   gpc1_1 gpc1042 (
      {stage0_15[493]},
      {stage1_15[253]}
   );
   gpc1_1 gpc1043 (
      {stage0_15[494]},
      {stage1_15[254]}
   );
   gpc1_1 gpc1044 (
      {stage0_15[495]},
      {stage1_15[255]}
   );
   gpc1_1 gpc1045 (
      {stage0_15[496]},
      {stage1_15[256]}
   );
   gpc1_1 gpc1046 (
      {stage0_15[497]},
      {stage1_15[257]}
   );
   gpc1_1 gpc1047 (
      {stage0_15[498]},
      {stage1_15[258]}
   );
   gpc1_1 gpc1048 (
      {stage0_15[499]},
      {stage1_15[259]}
   );
   gpc1_1 gpc1049 (
      {stage0_15[500]},
      {stage1_15[260]}
   );
   gpc1_1 gpc1050 (
      {stage0_15[501]},
      {stage1_15[261]}
   );
   gpc1_1 gpc1051 (
      {stage0_15[502]},
      {stage1_15[262]}
   );
   gpc1_1 gpc1052 (
      {stage0_15[503]},
      {stage1_15[263]}
   );
   gpc1_1 gpc1053 (
      {stage0_15[504]},
      {stage1_15[264]}
   );
   gpc1_1 gpc1054 (
      {stage0_15[505]},
      {stage1_15[265]}
   );
   gpc1_1 gpc1055 (
      {stage0_15[506]},
      {stage1_15[266]}
   );
   gpc1_1 gpc1056 (
      {stage0_15[507]},
      {stage1_15[267]}
   );
   gpc1_1 gpc1057 (
      {stage0_15[508]},
      {stage1_15[268]}
   );
   gpc1_1 gpc1058 (
      {stage0_15[509]},
      {stage1_15[269]}
   );
   gpc1_1 gpc1059 (
      {stage0_15[510]},
      {stage1_15[270]}
   );
   gpc1_1 gpc1060 (
      {stage0_15[511]},
      {stage1_15[271]}
   );
   gpc1163_5 gpc1061 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1062 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1063 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1064 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1065 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1066 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1067 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1068 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1069 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1070 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1071 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1072 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1073 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1074 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1075 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1076 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1077 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1078 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1079 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1080 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1081 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1082 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc615_5 gpc1083 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100]},
      {stage1_1[72]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1084 (
      {stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc1085 (
      {stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc1086 (
      {stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc1087 (
      {stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc1088 (
      {stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc1089 (
      {stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1090 (
      {stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1091 (
      {stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1092 (
      {stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1093 (
      {stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1094 (
      {stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1095 (
      {stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1096 (
      {stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc1097 (
      {stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc1098 (
      {stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc1099 (
      {stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc1100 (
      {stage1_1[169], stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc1101 (
      {stage1_1[175], stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], 1'b0},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc615_5 gpc1102 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[120]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1103 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[121]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1104 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[122]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1105 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[123]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc1106 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[124]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc1107 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[125]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc1108 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[126]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc1109 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[127]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc1110 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[128]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc1111 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[129]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc1112 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[130]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc1113 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[131]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc1114 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[132]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc1115 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[133]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[31],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc1116 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[134]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[32],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc1117 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[135]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[33],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc1118 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[136]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[34],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc1119 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[137]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[35],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc1120 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[138]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[36],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc615_5 gpc1121 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[114]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[19],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1122 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[115]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[20],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1123 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[116]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[21],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1124 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[117]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[22],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1125 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[118]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[23],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1126 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[119]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[24],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1127 (
      {stage1_3[169], stage1_3[170], stage1_3[171], stage1_3[172], stage1_3[173]},
      {stage1_4[120]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[25],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1128 (
      {stage1_3[174], stage1_3[175], stage1_3[176], stage1_3[177], stage1_3[178]},
      {stage1_4[121]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[26],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1129 (
      {stage1_3[179], stage1_3[180], stage1_3[181], stage1_3[182], stage1_3[183]},
      {stage1_4[122]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[27],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1130 (
      {stage1_3[184], stage1_3[185], stage1_3[186], stage1_3[187], stage1_3[188]},
      {stage1_4[123]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[28],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1131 (
      {stage1_3[189], stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193]},
      {stage1_4[124]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[29],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1132 (
      {stage1_3[194], stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198]},
      {stage1_4[125]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[30],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1133 (
      {stage1_3[199], stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203]},
      {stage1_4[126]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[31],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1134 (
      {stage1_3[204], stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208]},
      {stage1_4[127]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[32],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1135 (
      {stage1_3[209], stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213]},
      {stage1_4[128]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[33],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1136 (
      {stage1_3[214], stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218]},
      {stage1_4[129]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[34],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc606_5 gpc1137 (
      {stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[16],stage2_6[35],stage2_5[53],stage2_4[76]}
   );
   gpc606_5 gpc1138 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[17],stage2_6[36],stage2_5[54],stage2_4[77]}
   );
   gpc606_5 gpc1139 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[18],stage2_6[37],stage2_5[55],stage2_4[78]}
   );
   gpc606_5 gpc1140 (
      {stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[19],stage2_6[38],stage2_5[56],stage2_4[79]}
   );
   gpc606_5 gpc1141 (
      {stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[20],stage2_6[39],stage2_5[57],stage2_4[80]}
   );
   gpc606_5 gpc1142 (
      {stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[21],stage2_6[40],stage2_5[58],stage2_4[81]}
   );
   gpc606_5 gpc1143 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[22],stage2_6[41],stage2_5[59],stage2_4[82]}
   );
   gpc606_5 gpc1144 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[23],stage2_6[42],stage2_5[60],stage2_4[83]}
   );
   gpc606_5 gpc1145 (
      {stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[24],stage2_6[43],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc1146 (
      {stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[25],stage2_6[44],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc1147 (
      {stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[26],stage2_6[45],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc1148 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[27],stage2_6[46],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc1149 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206], stage1_4[207]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[28],stage2_6[47],stage2_5[65],stage2_4[88]}
   );
   gpc606_5 gpc1150 (
      {stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211], stage1_4[212], stage1_4[213]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[29],stage2_6[48],stage2_5[66],stage2_4[89]}
   );
   gpc606_5 gpc1151 (
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[14],stage2_7[30],stage2_6[49],stage2_5[67]}
   );
   gpc606_5 gpc1152 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[15],stage2_7[31],stage2_6[50],stage2_5[68]}
   );
   gpc606_5 gpc1153 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[16],stage2_7[32],stage2_6[51],stage2_5[69]}
   );
   gpc606_5 gpc1154 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[17],stage2_7[33],stage2_6[52],stage2_5[70]}
   );
   gpc606_5 gpc1155 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[18],stage2_7[34],stage2_6[53],stage2_5[71]}
   );
   gpc606_5 gpc1156 (
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[19],stage2_7[35],stage2_6[54],stage2_5[72]}
   );
   gpc606_5 gpc1157 (
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[20],stage2_7[36],stage2_6[55],stage2_5[73]}
   );
   gpc606_5 gpc1158 (
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[21],stage2_7[37],stage2_6[56],stage2_5[74]}
   );
   gpc606_5 gpc1159 (
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[22],stage2_7[38],stage2_6[57],stage2_5[75]}
   );
   gpc606_5 gpc1160 (
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[23],stage2_7[39],stage2_6[58],stage2_5[76]}
   );
   gpc606_5 gpc1161 (
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[24],stage2_7[40],stage2_6[59],stage2_5[77]}
   );
   gpc606_5 gpc1162 (
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[25],stage2_7[41],stage2_6[60],stage2_5[78]}
   );
   gpc606_5 gpc1163 (
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[26],stage2_7[42],stage2_6[61],stage2_5[79]}
   );
   gpc606_5 gpc1164 (
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[27],stage2_7[43],stage2_6[62],stage2_5[80]}
   );
   gpc606_5 gpc1165 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[28],stage2_7[44],stage2_6[63],stage2_5[81]}
   );
   gpc606_5 gpc1166 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[29],stage2_7[45],stage2_6[64],stage2_5[82]}
   );
   gpc606_5 gpc1167 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[30],stage2_7[46],stage2_6[65],stage2_5[83]}
   );
   gpc606_5 gpc1168 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[31],stage2_7[47],stage2_6[66],stage2_5[84]}
   );
   gpc606_5 gpc1169 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[32],stage2_7[48],stage2_6[67],stage2_5[85]}
   );
   gpc606_5 gpc1170 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[19],stage2_8[33],stage2_7[49],stage2_6[68]}
   );
   gpc606_5 gpc1171 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[20],stage2_8[34],stage2_7[50],stage2_6[69]}
   );
   gpc606_5 gpc1172 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[21],stage2_8[35],stage2_7[51],stage2_6[70]}
   );
   gpc606_5 gpc1173 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[22],stage2_8[36],stage2_7[52],stage2_6[71]}
   );
   gpc606_5 gpc1174 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[23],stage2_8[37],stage2_7[53],stage2_6[72]}
   );
   gpc606_5 gpc1175 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[24],stage2_8[38],stage2_7[54],stage2_6[73]}
   );
   gpc606_5 gpc1176 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[25],stage2_8[39],stage2_7[55],stage2_6[74]}
   );
   gpc606_5 gpc1177 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[26],stage2_8[40],stage2_7[56],stage2_6[75]}
   );
   gpc606_5 gpc1178 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[27],stage2_8[41],stage2_7[57],stage2_6[76]}
   );
   gpc606_5 gpc1179 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[28],stage2_8[42],stage2_7[58],stage2_6[77]}
   );
   gpc606_5 gpc1180 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[29],stage2_8[43],stage2_7[59],stage2_6[78]}
   );
   gpc606_5 gpc1181 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[30],stage2_8[44],stage2_7[60],stage2_6[79]}
   );
   gpc606_5 gpc1182 (
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[31],stage2_8[45],stage2_7[61],stage2_6[80]}
   );
   gpc606_5 gpc1183 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[32],stage2_8[46],stage2_7[62],stage2_6[81]}
   );
   gpc606_5 gpc1184 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[33],stage2_8[47],stage2_7[63],stage2_6[82]}
   );
   gpc615_5 gpc1185 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178]},
      {stage1_7[114]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[34],stage2_8[48],stage2_7[64],stage2_6[83]}
   );
   gpc615_5 gpc1186 (
      {stage1_6[179], stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183]},
      {stage1_7[115]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[35],stage2_8[49],stage2_7[65],stage2_6[84]}
   );
   gpc615_5 gpc1187 (
      {stage1_6[184], stage1_6[185], stage1_6[186], stage1_6[187], stage1_6[188]},
      {stage1_7[116]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[36],stage2_8[50],stage2_7[66],stage2_6[85]}
   );
   gpc615_5 gpc1188 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[108]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[18],stage2_9[37],stage2_8[51],stage2_7[67]}
   );
   gpc615_5 gpc1189 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[109]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[19],stage2_9[38],stage2_8[52],stage2_7[68]}
   );
   gpc615_5 gpc1190 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[110]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[20],stage2_9[39],stage2_8[53],stage2_7[69]}
   );
   gpc615_5 gpc1191 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[111]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[21],stage2_9[40],stage2_8[54],stage2_7[70]}
   );
   gpc615_5 gpc1192 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[112]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[22],stage2_9[41],stage2_8[55],stage2_7[71]}
   );
   gpc615_5 gpc1193 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[113]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[23],stage2_9[42],stage2_8[56],stage2_7[72]}
   );
   gpc615_5 gpc1194 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[114]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[24],stage2_9[43],stage2_8[57],stage2_7[73]}
   );
   gpc615_5 gpc1195 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[115]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[25],stage2_9[44],stage2_8[58],stage2_7[74]}
   );
   gpc615_5 gpc1196 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[116]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[26],stage2_9[45],stage2_8[59],stage2_7[75]}
   );
   gpc615_5 gpc1197 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[117]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[27],stage2_9[46],stage2_8[60],stage2_7[76]}
   );
   gpc615_5 gpc1198 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[118]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[28],stage2_9[47],stage2_8[61],stage2_7[77]}
   );
   gpc615_5 gpc1199 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[119]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[29],stage2_9[48],stage2_8[62],stage2_7[78]}
   );
   gpc615_5 gpc1200 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[120]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[30],stage2_9[49],stage2_8[63],stage2_7[79]}
   );
   gpc615_5 gpc1201 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[121]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[31],stage2_9[50],stage2_8[64],stage2_7[80]}
   );
   gpc615_5 gpc1202 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[122]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[32],stage2_9[51],stage2_8[65],stage2_7[81]}
   );
   gpc615_5 gpc1203 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[123]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[33],stage2_9[52],stage2_8[66],stage2_7[82]}
   );
   gpc615_5 gpc1204 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[124]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[34],stage2_9[53],stage2_8[67],stage2_7[83]}
   );
   gpc615_5 gpc1205 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[125]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[35],stage2_9[54],stage2_8[68],stage2_7[84]}
   );
   gpc606_5 gpc1206 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[18],stage2_10[36],stage2_9[55],stage2_8[69]}
   );
   gpc606_5 gpc1207 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[19],stage2_10[37],stage2_9[56],stage2_8[70]}
   );
   gpc615_5 gpc1208 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142]},
      {stage1_9[108]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[20],stage2_10[38],stage2_9[57],stage2_8[71]}
   );
   gpc615_5 gpc1209 (
      {stage1_8[143], stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147]},
      {stage1_9[109]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[21],stage2_10[39],stage2_9[58],stage2_8[72]}
   );
   gpc615_5 gpc1210 (
      {stage1_8[148], stage1_8[149], stage1_8[150], stage1_8[151], stage1_8[152]},
      {stage1_9[110]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[22],stage2_10[40],stage2_9[59],stage2_8[73]}
   );
   gpc615_5 gpc1211 (
      {stage1_8[153], stage1_8[154], stage1_8[155], stage1_8[156], stage1_8[157]},
      {stage1_9[111]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[23],stage2_10[41],stage2_9[60],stage2_8[74]}
   );
   gpc615_5 gpc1212 (
      {stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161], stage1_8[162]},
      {stage1_9[112]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[24],stage2_10[42],stage2_9[61],stage2_8[75]}
   );
   gpc615_5 gpc1213 (
      {stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_9[113]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[25],stage2_10[43],stage2_9[62],stage2_8[76]}
   );
   gpc615_5 gpc1214 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172]},
      {stage1_9[114]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[26],stage2_10[44],stage2_9[63],stage2_8[77]}
   );
   gpc615_5 gpc1215 (
      {stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_9[115]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[27],stage2_10[45],stage2_9[64],stage2_8[78]}
   );
   gpc615_5 gpc1216 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_9[116]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[28],stage2_10[46],stage2_9[65],stage2_8[79]}
   );
   gpc615_5 gpc1217 (
      {stage1_8[183], stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187]},
      {stage1_9[117]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[29],stage2_10[47],stage2_9[66],stage2_8[80]}
   );
   gpc615_5 gpc1218 (
      {stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_9[118]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[30],stage2_10[48],stage2_9[67],stage2_8[81]}
   );
   gpc615_5 gpc1219 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197]},
      {stage1_9[119]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[31],stage2_10[49],stage2_9[68],stage2_8[82]}
   );
   gpc615_5 gpc1220 (
      {stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202]},
      {stage1_9[120]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[32],stage2_10[50],stage2_9[69],stage2_8[83]}
   );
   gpc615_5 gpc1221 (
      {stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_9[121]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[33],stage2_10[51],stage2_9[70],stage2_8[84]}
   );
   gpc615_5 gpc1222 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212]},
      {stage1_9[122]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[34],stage2_10[52],stage2_9[71],stage2_8[85]}
   );
   gpc615_5 gpc1223 (
      {stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217]},
      {stage1_9[123]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[35],stage2_10[53],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc1224 (
      {stage1_9[124], stage1_9[125], stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[36],stage2_10[54],stage2_9[73]}
   );
   gpc606_5 gpc1225 (
      {stage1_9[130], stage1_9[131], stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[37],stage2_10[55],stage2_9[74]}
   );
   gpc606_5 gpc1226 (
      {stage1_9[136], stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[38],stage2_10[56],stage2_9[75]}
   );
   gpc606_5 gpc1227 (
      {stage1_9[142], stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[21],stage2_11[39],stage2_10[57],stage2_9[76]}
   );
   gpc606_5 gpc1228 (
      {stage1_9[148], stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[22],stage2_11[40],stage2_10[58],stage2_9[77]}
   );
   gpc606_5 gpc1229 (
      {stage1_9[154], stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[23],stage2_11[41],stage2_10[59],stage2_9[78]}
   );
   gpc606_5 gpc1230 (
      {stage1_9[160], stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[24],stage2_11[42],stage2_10[60],stage2_9[79]}
   );
   gpc606_5 gpc1231 (
      {stage1_9[166], stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[25],stage2_11[43],stage2_10[61],stage2_9[80]}
   );
   gpc606_5 gpc1232 (
      {stage1_9[172], stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[26],stage2_11[44],stage2_10[62],stage2_9[81]}
   );
   gpc606_5 gpc1233 (
      {stage1_9[178], stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[27],stage2_11[45],stage2_10[63],stage2_9[82]}
   );
   gpc606_5 gpc1234 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[28],stage2_11[46],stage2_10[64],stage2_9[83]}
   );
   gpc606_5 gpc1235 (
      {stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[29],stage2_11[47],stage2_10[65],stage2_9[84]}
   );
   gpc606_5 gpc1236 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[30],stage2_11[48],stage2_10[66],stage2_9[85]}
   );
   gpc606_5 gpc1237 (
      {stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[31],stage2_11[49],stage2_10[67],stage2_9[86]}
   );
   gpc606_5 gpc1238 (
      {stage1_9[208], stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[32],stage2_11[50],stage2_10[68],stage2_9[87]}
   );
   gpc606_5 gpc1239 (
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[15],stage2_12[33],stage2_11[51],stage2_10[69]}
   );
   gpc606_5 gpc1240 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[16],stage2_12[34],stage2_11[52],stage2_10[70]}
   );
   gpc606_5 gpc1241 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[17],stage2_12[35],stage2_11[53],stage2_10[71]}
   );
   gpc606_5 gpc1242 (
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[18],stage2_12[36],stage2_11[54],stage2_10[72]}
   );
   gpc606_5 gpc1243 (
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[19],stage2_12[37],stage2_11[55],stage2_10[73]}
   );
   gpc606_5 gpc1244 (
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[20],stage2_12[38],stage2_11[56],stage2_10[74]}
   );
   gpc606_5 gpc1245 (
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[21],stage2_12[39],stage2_11[57],stage2_10[75]}
   );
   gpc606_5 gpc1246 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[22],stage2_12[40],stage2_11[58],stage2_10[76]}
   );
   gpc606_5 gpc1247 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[23],stage2_12[41],stage2_11[59],stage2_10[77]}
   );
   gpc606_5 gpc1248 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[24],stage2_12[42],stage2_11[60],stage2_10[78]}
   );
   gpc606_5 gpc1249 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[25],stage2_12[43],stage2_11[61],stage2_10[79]}
   );
   gpc606_5 gpc1250 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[26],stage2_12[44],stage2_11[62],stage2_10[80]}
   );
   gpc606_5 gpc1251 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[27],stage2_12[45],stage2_11[63],stage2_10[81]}
   );
   gpc606_5 gpc1252 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[28],stage2_12[46],stage2_11[64],stage2_10[82]}
   );
   gpc606_5 gpc1253 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[29],stage2_12[47],stage2_11[65],stage2_10[83]}
   );
   gpc606_5 gpc1254 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[30],stage2_12[48],stage2_11[66],stage2_10[84]}
   );
   gpc606_5 gpc1255 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[31],stage2_12[49],stage2_11[67],stage2_10[85]}
   );
   gpc615_5 gpc1256 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[17],stage2_13[32],stage2_12[50],stage2_11[68]}
   );
   gpc615_5 gpc1257 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[103]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[18],stage2_13[33],stage2_12[51],stage2_11[69]}
   );
   gpc615_5 gpc1258 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[104]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[19],stage2_13[34],stage2_12[52],stage2_11[70]}
   );
   gpc615_5 gpc1259 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[105]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[20],stage2_13[35],stage2_12[53],stage2_11[71]}
   );
   gpc615_5 gpc1260 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[106]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[21],stage2_13[36],stage2_12[54],stage2_11[72]}
   );
   gpc615_5 gpc1261 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[107]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[22],stage2_13[37],stage2_12[55],stage2_11[73]}
   );
   gpc606_5 gpc1262 (
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[23],stage2_13[38],stage2_12[56]}
   );
   gpc606_5 gpc1263 (
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[24],stage2_13[39],stage2_12[57]}
   );
   gpc606_5 gpc1264 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[8],stage2_14[25],stage2_13[40],stage2_12[58]}
   );
   gpc606_5 gpc1265 (
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[9],stage2_14[26],stage2_13[41],stage2_12[59]}
   );
   gpc606_5 gpc1266 (
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[10],stage2_14[27],stage2_13[42],stage2_12[60]}
   );
   gpc606_5 gpc1267 (
      {stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[11],stage2_14[28],stage2_13[43],stage2_12[61]}
   );
   gpc606_5 gpc1268 (
      {stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[12],stage2_14[29],stage2_13[44],stage2_12[62]}
   );
   gpc606_5 gpc1269 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[13],stage2_14[30],stage2_13[45],stage2_12[63]}
   );
   gpc606_5 gpc1270 (
      {stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[14],stage2_14[31],stage2_13[46],stage2_12[64]}
   );
   gpc606_5 gpc1271 (
      {stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[15],stage2_14[32],stage2_13[47],stage2_12[65]}
   );
   gpc606_5 gpc1272 (
      {stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[16],stage2_14[33],stage2_13[48],stage2_12[66]}
   );
   gpc606_5 gpc1273 (
      {stage1_12[174], stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[17],stage2_14[34],stage2_13[49],stage2_12[67]}
   );
   gpc606_5 gpc1274 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[18],stage2_14[35],stage2_13[50],stage2_12[68]}
   );
   gpc606_5 gpc1275 (
      {stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[19],stage2_14[36],stage2_13[51],stage2_12[69]}
   );
   gpc606_5 gpc1276 (
      {stage1_12[192], stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[20],stage2_14[37],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc1277 (
      {stage1_12[198], stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[21],stage2_14[38],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc1278 (
      {stage1_12[204], stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[22],stage2_14[39],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc1279 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[17],stage2_15[23],stage2_14[40],stage2_13[55]}
   );
   gpc606_5 gpc1280 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[18],stage2_15[24],stage2_14[41],stage2_13[56]}
   );
   gpc606_5 gpc1281 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[19],stage2_15[25],stage2_14[42],stage2_13[57]}
   );
   gpc606_5 gpc1282 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[20],stage2_15[26],stage2_14[43],stage2_13[58]}
   );
   gpc606_5 gpc1283 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[21],stage2_15[27],stage2_14[44],stage2_13[59]}
   );
   gpc606_5 gpc1284 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[22],stage2_15[28],stage2_14[45],stage2_13[60]}
   );
   gpc606_5 gpc1285 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[23],stage2_15[29],stage2_14[46],stage2_13[61]}
   );
   gpc606_5 gpc1286 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[24],stage2_15[30],stage2_14[47],stage2_13[62]}
   );
   gpc606_5 gpc1287 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[25],stage2_15[31],stage2_14[48],stage2_13[63]}
   );
   gpc606_5 gpc1288 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[26],stage2_15[32],stage2_14[49],stage2_13[64]}
   );
   gpc606_5 gpc1289 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[27],stage2_15[33],stage2_14[50],stage2_13[65]}
   );
   gpc606_5 gpc1290 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[28],stage2_15[34],stage2_14[51],stage2_13[66]}
   );
   gpc606_5 gpc1291 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[29],stage2_15[35],stage2_14[52],stage2_13[67]}
   );
   gpc606_5 gpc1292 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[30],stage2_15[36],stage2_14[53],stage2_13[68]}
   );
   gpc606_5 gpc1293 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[31],stage2_15[37],stage2_14[54],stage2_13[69]}
   );
   gpc606_5 gpc1294 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[32],stage2_15[38],stage2_14[55],stage2_13[70]}
   );
   gpc615_5 gpc1295 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136]},
      {stage1_14[102]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[33],stage2_15[39],stage2_14[56],stage2_13[71]}
   );
   gpc615_5 gpc1296 (
      {stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141]},
      {stage1_14[103]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[34],stage2_15[40],stage2_14[57],stage2_13[72]}
   );
   gpc615_5 gpc1297 (
      {stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage1_14[104]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[35],stage2_15[41],stage2_14[58],stage2_13[73]}
   );
   gpc615_5 gpc1298 (
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151]},
      {stage1_14[105]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[36],stage2_15[42],stage2_14[59],stage2_13[74]}
   );
   gpc615_5 gpc1299 (
      {stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156]},
      {stage1_14[106]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[37],stage2_15[43],stage2_14[60],stage2_13[75]}
   );
   gpc615_5 gpc1300 (
      {stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_14[107]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[38],stage2_15[44],stage2_14[61],stage2_13[76]}
   );
   gpc615_5 gpc1301 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166]},
      {stage1_14[108]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage2_17[22],stage2_16[39],stage2_15[45],stage2_14[62],stage2_13[77]}
   );
   gpc615_5 gpc1302 (
      {stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171]},
      {stage1_14[109]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage2_17[23],stage2_16[40],stage2_15[46],stage2_14[63],stage2_13[78]}
   );
   gpc615_5 gpc1303 (
      {stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage1_14[110]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage2_17[24],stage2_16[41],stage2_15[47],stage2_14[64],stage2_13[79]}
   );
   gpc615_5 gpc1304 (
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181]},
      {stage1_14[111]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage2_17[25],stage2_16[42],stage2_15[48],stage2_14[65],stage2_13[80]}
   );
   gpc615_5 gpc1305 (
      {stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185], stage1_13[186]},
      {stage1_14[112]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage2_17[26],stage2_16[43],stage2_15[49],stage2_14[66],stage2_13[81]}
   );
   gpc615_5 gpc1306 (
      {stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_14[113]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage2_17[27],stage2_16[44],stage2_15[50],stage2_14[67],stage2_13[82]}
   );
   gpc615_5 gpc1307 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196]},
      {stage1_14[114]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage2_17[28],stage2_16[45],stage2_15[51],stage2_14[68],stage2_13[83]}
   );
   gpc615_5 gpc1308 (
      {stage1_13[197], stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201]},
      {stage1_14[115]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage2_17[29],stage2_16[46],stage2_15[52],stage2_14[69],stage2_13[84]}
   );
   gpc615_5 gpc1309 (
      {stage1_13[202], stage1_13[203], stage1_13[204], stage1_13[205], stage1_13[206]},
      {stage1_14[116]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage2_17[30],stage2_16[47],stage2_15[53],stage2_14[70],stage2_13[85]}
   );
   gpc615_5 gpc1310 (
      {stage1_13[207], stage1_13[208], stage1_13[209], stage1_13[210], stage1_13[211]},
      {stage1_14[117]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage2_17[31],stage2_16[48],stage2_15[54],stage2_14[71],stage2_13[86]}
   );
   gpc615_5 gpc1311 (
      {stage1_13[212], stage1_13[213], stage1_13[214], stage1_13[215], stage1_13[216]},
      {stage1_14[118]},
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196], stage1_15[197]},
      {stage2_17[32],stage2_16[49],stage2_15[55],stage2_14[72],stage2_13[87]}
   );
   gpc615_5 gpc1312 (
      {stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_14[119]},
      {stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201], stage1_15[202], stage1_15[203]},
      {stage2_17[33],stage2_16[50],stage2_15[56],stage2_14[73],stage2_13[88]}
   );
   gpc615_5 gpc1313 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226]},
      {stage1_14[120]},
      {stage1_15[204], stage1_15[205], stage1_15[206], stage1_15[207], stage1_15[208], stage1_15[209]},
      {stage2_17[34],stage2_16[51],stage2_15[57],stage2_14[74],stage2_13[89]}
   );
   gpc615_5 gpc1314 (
      {stage1_13[227], stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231]},
      {stage1_14[121]},
      {stage1_15[210], stage1_15[211], stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215]},
      {stage2_17[35],stage2_16[52],stage2_15[58],stage2_14[75],stage2_13[90]}
   );
   gpc606_5 gpc1315 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[36],stage2_16[53],stage2_15[59],stage2_14[76]}
   );
   gpc606_5 gpc1316 (
      {stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[37],stage2_16[54],stage2_15[60],stage2_14[77]}
   );
   gpc606_5 gpc1317 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[38],stage2_16[55],stage2_15[61],stage2_14[78]}
   );
   gpc606_5 gpc1318 (
      {stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[39],stage2_16[56],stage2_15[62],stage2_14[79]}
   );
   gpc606_5 gpc1319 (
      {stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[40],stage2_16[57],stage2_15[63],stage2_14[80]}
   );
   gpc606_5 gpc1320 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[41],stage2_16[58],stage2_15[64],stage2_14[81]}
   );
   gpc606_5 gpc1321 (
      {stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[42],stage2_16[59],stage2_15[65],stage2_14[82]}
   );
   gpc606_5 gpc1322 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[43],stage2_16[60],stage2_15[66],stage2_14[83]}
   );
   gpc606_5 gpc1323 (
      {stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[44],stage2_16[61],stage2_15[67],stage2_14[84]}
   );
   gpc606_5 gpc1324 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[45],stage2_16[62],stage2_15[68],stage2_14[85]}
   );
   gpc606_5 gpc1325 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186], stage1_14[187]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[46],stage2_16[63],stage2_15[69],stage2_14[86]}
   );
   gpc606_5 gpc1326 (
      {stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191], stage1_14[192], stage1_14[193]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[47],stage2_16[64],stage2_15[70],stage2_14[87]}
   );
   gpc606_5 gpc1327 (
      {stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[48],stage2_16[65],stage2_15[71],stage2_14[88]}
   );
   gpc606_5 gpc1328 (
      {stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[49],stage2_16[66],stage2_15[72],stage2_14[89]}
   );
   gpc615_5 gpc1329 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[216]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[50],stage2_16[67],stage2_15[73],stage2_14[90]}
   );
   gpc615_5 gpc1330 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[90]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[15],stage2_17[51],stage2_16[68],stage2_15[74]}
   );
   gpc615_5 gpc1331 (
      {stage1_15[222], stage1_15[223], stage1_15[224], stage1_15[225], stage1_15[226]},
      {stage1_16[91]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[16],stage2_17[52],stage2_16[69],stage2_15[75]}
   );
   gpc615_5 gpc1332 (
      {stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230], stage1_15[231]},
      {stage1_16[92]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[17],stage2_17[53],stage2_16[70],stage2_15[76]}
   );
   gpc615_5 gpc1333 (
      {stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_16[93]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[18],stage2_17[54],stage2_16[71],stage2_15[77]}
   );
   gpc615_5 gpc1334 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241]},
      {stage1_16[94]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[19],stage2_17[55],stage2_16[72],stage2_15[78]}
   );
   gpc615_5 gpc1335 (
      {stage1_15[242], stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246]},
      {stage1_16[95]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[20],stage2_17[56],stage2_16[73],stage2_15[79]}
   );
   gpc615_5 gpc1336 (
      {stage1_15[247], stage1_15[248], stage1_15[249], stage1_15[250], stage1_15[251]},
      {stage1_16[96]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[21],stage2_17[57],stage2_16[74],stage2_15[80]}
   );
   gpc615_5 gpc1337 (
      {stage1_15[252], stage1_15[253], stage1_15[254], stage1_15[255], stage1_15[256]},
      {stage1_16[97]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[22],stage2_17[58],stage2_16[75],stage2_15[81]}
   );
   gpc615_5 gpc1338 (
      {stage1_15[257], stage1_15[258], stage1_15[259], stage1_15[260], stage1_15[261]},
      {stage1_16[98]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[23],stage2_17[59],stage2_16[76],stage2_15[82]}
   );
   gpc615_5 gpc1339 (
      {stage1_15[262], stage1_15[263], stage1_15[264], stage1_15[265], stage1_15[266]},
      {stage1_16[99]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[24],stage2_17[60],stage2_16[77],stage2_15[83]}
   );
   gpc615_5 gpc1340 (
      {stage1_15[267], stage1_15[268], stage1_15[269], stage1_15[270], stage1_15[271]},
      {stage1_16[100]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], 1'b0, 1'b0},
      {stage2_19[10],stage2_18[25],stage2_17[61],stage2_16[78],stage2_15[84]}
   );
   gpc1_1 gpc1341 (
      {stage1_3[219]},
      {stage2_3[76]}
   );
   gpc1_1 gpc1342 (
      {stage1_3[220]},
      {stage2_3[77]}
   );
   gpc1_1 gpc1343 (
      {stage1_3[221]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1344 (
      {stage1_3[222]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1345 (
      {stage1_3[223]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1346 (
      {stage1_3[224]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1347 (
      {stage1_3[225]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1348 (
      {stage1_3[226]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1349 (
      {stage1_3[227]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1350 (
      {stage1_3[228]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1351 (
      {stage1_3[229]},
      {stage2_3[86]}
   );
   gpc1_1 gpc1352 (
      {stage1_3[230]},
      {stage2_3[87]}
   );
   gpc1_1 gpc1353 (
      {stage1_3[231]},
      {stage2_3[88]}
   );
   gpc1_1 gpc1354 (
      {stage1_3[232]},
      {stage2_3[89]}
   );
   gpc1_1 gpc1355 (
      {stage1_3[233]},
      {stage2_3[90]}
   );
   gpc1_1 gpc1356 (
      {stage1_3[234]},
      {stage2_3[91]}
   );
   gpc1_1 gpc1357 (
      {stage1_3[235]},
      {stage2_3[92]}
   );
   gpc1_1 gpc1358 (
      {stage1_3[236]},
      {stage2_3[93]}
   );
   gpc1_1 gpc1359 (
      {stage1_3[237]},
      {stage2_3[94]}
   );
   gpc1_1 gpc1360 (
      {stage1_3[238]},
      {stage2_3[95]}
   );
   gpc1_1 gpc1361 (
      {stage1_3[239]},
      {stage2_3[96]}
   );
   gpc1_1 gpc1362 (
      {stage1_3[240]},
      {stage2_3[97]}
   );
   gpc1_1 gpc1363 (
      {stage1_3[241]},
      {stage2_3[98]}
   );
   gpc1_1 gpc1364 (
      {stage1_3[242]},
      {stage2_3[99]}
   );
   gpc1_1 gpc1365 (
      {stage1_3[243]},
      {stage2_3[100]}
   );
   gpc1_1 gpc1366 (
      {stage1_3[244]},
      {stage2_3[101]}
   );
   gpc1_1 gpc1367 (
      {stage1_3[245]},
      {stage2_3[102]}
   );
   gpc1_1 gpc1368 (
      {stage1_4[214]},
      {stage2_4[90]}
   );
   gpc1_1 gpc1369 (
      {stage1_4[215]},
      {stage2_4[91]}
   );
   gpc1_1 gpc1370 (
      {stage1_4[216]},
      {stage2_4[92]}
   );
   gpc1_1 gpc1371 (
      {stage1_4[217]},
      {stage2_4[93]}
   );
   gpc1_1 gpc1372 (
      {stage1_4[218]},
      {stage2_4[94]}
   );
   gpc1_1 gpc1373 (
      {stage1_4[219]},
      {stage2_4[95]}
   );
   gpc1_1 gpc1374 (
      {stage1_4[220]},
      {stage2_4[96]}
   );
   gpc1_1 gpc1375 (
      {stage1_4[221]},
      {stage2_4[97]}
   );
   gpc1_1 gpc1376 (
      {stage1_4[222]},
      {stage2_4[98]}
   );
   gpc1_1 gpc1377 (
      {stage1_4[223]},
      {stage2_4[99]}
   );
   gpc1_1 gpc1378 (
      {stage1_4[224]},
      {stage2_4[100]}
   );
   gpc1_1 gpc1379 (
      {stage1_4[225]},
      {stage2_4[101]}
   );
   gpc1_1 gpc1380 (
      {stage1_4[226]},
      {stage2_4[102]}
   );
   gpc1_1 gpc1381 (
      {stage1_4[227]},
      {stage2_4[103]}
   );
   gpc1_1 gpc1382 (
      {stage1_4[228]},
      {stage2_4[104]}
   );
   gpc1_1 gpc1383 (
      {stage1_4[229]},
      {stage2_4[105]}
   );
   gpc1_1 gpc1384 (
      {stage1_4[230]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1385 (
      {stage1_4[231]},
      {stage2_4[107]}
   );
   gpc1_1 gpc1386 (
      {stage1_4[232]},
      {stage2_4[108]}
   );
   gpc1_1 gpc1387 (
      {stage1_4[233]},
      {stage2_4[109]}
   );
   gpc1_1 gpc1388 (
      {stage1_4[234]},
      {stage2_4[110]}
   );
   gpc1_1 gpc1389 (
      {stage1_4[235]},
      {stage2_4[111]}
   );
   gpc1_1 gpc1390 (
      {stage1_4[236]},
      {stage2_4[112]}
   );
   gpc1_1 gpc1391 (
      {stage1_4[237]},
      {stage2_4[113]}
   );
   gpc1_1 gpc1392 (
      {stage1_4[238]},
      {stage2_4[114]}
   );
   gpc1_1 gpc1393 (
      {stage1_4[239]},
      {stage2_4[115]}
   );
   gpc1_1 gpc1394 (
      {stage1_4[240]},
      {stage2_4[116]}
   );
   gpc1_1 gpc1395 (
      {stage1_5[210]},
      {stage2_5[86]}
   );
   gpc1_1 gpc1396 (
      {stage1_5[211]},
      {stage2_5[87]}
   );
   gpc1_1 gpc1397 (
      {stage1_5[212]},
      {stage2_5[88]}
   );
   gpc1_1 gpc1398 (
      {stage1_5[213]},
      {stage2_5[89]}
   );
   gpc1_1 gpc1399 (
      {stage1_5[214]},
      {stage2_5[90]}
   );
   gpc1_1 gpc1400 (
      {stage1_5[215]},
      {stage2_5[91]}
   );
   gpc1_1 gpc1401 (
      {stage1_5[216]},
      {stage2_5[92]}
   );
   gpc1_1 gpc1402 (
      {stage1_5[217]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1403 (
      {stage1_6[189]},
      {stage2_6[86]}
   );
   gpc1_1 gpc1404 (
      {stage1_6[190]},
      {stage2_6[87]}
   );
   gpc1_1 gpc1405 (
      {stage1_6[191]},
      {stage2_6[88]}
   );
   gpc1_1 gpc1406 (
      {stage1_6[192]},
      {stage2_6[89]}
   );
   gpc1_1 gpc1407 (
      {stage1_6[193]},
      {stage2_6[90]}
   );
   gpc1_1 gpc1408 (
      {stage1_6[194]},
      {stage2_6[91]}
   );
   gpc1_1 gpc1409 (
      {stage1_6[195]},
      {stage2_6[92]}
   );
   gpc1_1 gpc1410 (
      {stage1_6[196]},
      {stage2_6[93]}
   );
   gpc1_1 gpc1411 (
      {stage1_6[197]},
      {stage2_6[94]}
   );
   gpc1_1 gpc1412 (
      {stage1_6[198]},
      {stage2_6[95]}
   );
   gpc1_1 gpc1413 (
      {stage1_6[199]},
      {stage2_6[96]}
   );
   gpc1_1 gpc1414 (
      {stage1_6[200]},
      {stage2_6[97]}
   );
   gpc1_1 gpc1415 (
      {stage1_6[201]},
      {stage2_6[98]}
   );
   gpc1_1 gpc1416 (
      {stage1_6[202]},
      {stage2_6[99]}
   );
   gpc1_1 gpc1417 (
      {stage1_6[203]},
      {stage2_6[100]}
   );
   gpc1_1 gpc1418 (
      {stage1_6[204]},
      {stage2_6[101]}
   );
   gpc1_1 gpc1419 (
      {stage1_6[205]},
      {stage2_6[102]}
   );
   gpc1_1 gpc1420 (
      {stage1_6[206]},
      {stage2_6[103]}
   );
   gpc1_1 gpc1421 (
      {stage1_9[214]},
      {stage2_9[88]}
   );
   gpc1_1 gpc1422 (
      {stage1_9[215]},
      {stage2_9[89]}
   );
   gpc1_1 gpc1423 (
      {stage1_9[216]},
      {stage2_9[90]}
   );
   gpc1_1 gpc1424 (
      {stage1_9[217]},
      {stage2_9[91]}
   );
   gpc1_1 gpc1425 (
      {stage1_9[218]},
      {stage2_9[92]}
   );
   gpc1_1 gpc1426 (
      {stage1_9[219]},
      {stage2_9[93]}
   );
   gpc1_1 gpc1427 (
      {stage1_9[220]},
      {stage2_9[94]}
   );
   gpc1_1 gpc1428 (
      {stage1_9[221]},
      {stage2_9[95]}
   );
   gpc1_1 gpc1429 (
      {stage1_9[222]},
      {stage2_9[96]}
   );
   gpc1_1 gpc1430 (
      {stage1_9[223]},
      {stage2_9[97]}
   );
   gpc1_1 gpc1431 (
      {stage1_9[224]},
      {stage2_9[98]}
   );
   gpc1_1 gpc1432 (
      {stage1_9[225]},
      {stage2_9[99]}
   );
   gpc1_1 gpc1433 (
      {stage1_9[226]},
      {stage2_9[100]}
   );
   gpc1_1 gpc1434 (
      {stage1_9[227]},
      {stage2_9[101]}
   );
   gpc1_1 gpc1435 (
      {stage1_9[228]},
      {stage2_9[102]}
   );
   gpc1_1 gpc1436 (
      {stage1_9[229]},
      {stage2_9[103]}
   );
   gpc1_1 gpc1437 (
      {stage1_9[230]},
      {stage2_9[104]}
   );
   gpc1_1 gpc1438 (
      {stage1_9[231]},
      {stage2_9[105]}
   );
   gpc1_1 gpc1439 (
      {stage1_9[232]},
      {stage2_9[106]}
   );
   gpc1_1 gpc1440 (
      {stage1_9[233]},
      {stage2_9[107]}
   );
   gpc1_1 gpc1441 (
      {stage1_9[234]},
      {stage2_9[108]}
   );
   gpc1_1 gpc1442 (
      {stage1_9[235]},
      {stage2_9[109]}
   );
   gpc1_1 gpc1443 (
      {stage1_9[236]},
      {stage2_9[110]}
   );
   gpc1_1 gpc1444 (
      {stage1_9[237]},
      {stage2_9[111]}
   );
   gpc1_1 gpc1445 (
      {stage1_9[238]},
      {stage2_9[112]}
   );
   gpc1_1 gpc1446 (
      {stage1_9[239]},
      {stage2_9[113]}
   );
   gpc1_1 gpc1447 (
      {stage1_9[240]},
      {stage2_9[114]}
   );
   gpc1_1 gpc1448 (
      {stage1_9[241]},
      {stage2_9[115]}
   );
   gpc1_1 gpc1449 (
      {stage1_9[242]},
      {stage2_9[116]}
   );
   gpc1_1 gpc1450 (
      {stage1_9[243]},
      {stage2_9[117]}
   );
   gpc1_1 gpc1451 (
      {stage1_9[244]},
      {stage2_9[118]}
   );
   gpc1_1 gpc1452 (
      {stage1_9[245]},
      {stage2_9[119]}
   );
   gpc1_1 gpc1453 (
      {stage1_9[246]},
      {stage2_9[120]}
   );
   gpc1_1 gpc1454 (
      {stage1_9[247]},
      {stage2_9[121]}
   );
   gpc1_1 gpc1455 (
      {stage1_9[248]},
      {stage2_9[122]}
   );
   gpc1_1 gpc1456 (
      {stage1_9[249]},
      {stage2_9[123]}
   );
   gpc1_1 gpc1457 (
      {stage1_9[250]},
      {stage2_9[124]}
   );
   gpc1_1 gpc1458 (
      {stage1_9[251]},
      {stage2_9[125]}
   );
   gpc1_1 gpc1459 (
      {stage1_9[252]},
      {stage2_9[126]}
   );
   gpc1_1 gpc1460 (
      {stage1_9[253]},
      {stage2_9[127]}
   );
   gpc1_1 gpc1461 (
      {stage1_9[254]},
      {stage2_9[128]}
   );
   gpc1_1 gpc1462 (
      {stage1_9[255]},
      {stage2_9[129]}
   );
   gpc1_1 gpc1463 (
      {stage1_9[256]},
      {stage2_9[130]}
   );
   gpc1_1 gpc1464 (
      {stage1_9[257]},
      {stage2_9[131]}
   );
   gpc1_1 gpc1465 (
      {stage1_9[258]},
      {stage2_9[132]}
   );
   gpc1_1 gpc1466 (
      {stage1_9[259]},
      {stage2_9[133]}
   );
   gpc1_1 gpc1467 (
      {stage1_9[260]},
      {stage2_9[134]}
   );
   gpc1_1 gpc1468 (
      {stage1_9[261]},
      {stage2_9[135]}
   );
   gpc1_1 gpc1469 (
      {stage1_9[262]},
      {stage2_9[136]}
   );
   gpc1_1 gpc1470 (
      {stage1_9[263]},
      {stage2_9[137]}
   );
   gpc1_1 gpc1471 (
      {stage1_11[120]},
      {stage2_11[74]}
   );
   gpc1_1 gpc1472 (
      {stage1_11[121]},
      {stage2_11[75]}
   );
   gpc1_1 gpc1473 (
      {stage1_11[122]},
      {stage2_11[76]}
   );
   gpc1_1 gpc1474 (
      {stage1_11[123]},
      {stage2_11[77]}
   );
   gpc1_1 gpc1475 (
      {stage1_11[124]},
      {stage2_11[78]}
   );
   gpc1_1 gpc1476 (
      {stage1_11[125]},
      {stage2_11[79]}
   );
   gpc1_1 gpc1477 (
      {stage1_11[126]},
      {stage2_11[80]}
   );
   gpc1_1 gpc1478 (
      {stage1_11[127]},
      {stage2_11[81]}
   );
   gpc1_1 gpc1479 (
      {stage1_11[128]},
      {stage2_11[82]}
   );
   gpc1_1 gpc1480 (
      {stage1_11[129]},
      {stage2_11[83]}
   );
   gpc1_1 gpc1481 (
      {stage1_11[130]},
      {stage2_11[84]}
   );
   gpc1_1 gpc1482 (
      {stage1_11[131]},
      {stage2_11[85]}
   );
   gpc1_1 gpc1483 (
      {stage1_11[132]},
      {stage2_11[86]}
   );
   gpc1_1 gpc1484 (
      {stage1_11[133]},
      {stage2_11[87]}
   );
   gpc1_1 gpc1485 (
      {stage1_11[134]},
      {stage2_11[88]}
   );
   gpc1_1 gpc1486 (
      {stage1_11[135]},
      {stage2_11[89]}
   );
   gpc1_1 gpc1487 (
      {stage1_11[136]},
      {stage2_11[90]}
   );
   gpc1_1 gpc1488 (
      {stage1_11[137]},
      {stage2_11[91]}
   );
   gpc1_1 gpc1489 (
      {stage1_11[138]},
      {stage2_11[92]}
   );
   gpc1_1 gpc1490 (
      {stage1_11[139]},
      {stage2_11[93]}
   );
   gpc1_1 gpc1491 (
      {stage1_11[140]},
      {stage2_11[94]}
   );
   gpc1_1 gpc1492 (
      {stage1_11[141]},
      {stage2_11[95]}
   );
   gpc1_1 gpc1493 (
      {stage1_11[142]},
      {stage2_11[96]}
   );
   gpc1_1 gpc1494 (
      {stage1_11[143]},
      {stage2_11[97]}
   );
   gpc1_1 gpc1495 (
      {stage1_11[144]},
      {stage2_11[98]}
   );
   gpc1_1 gpc1496 (
      {stage1_11[145]},
      {stage2_11[99]}
   );
   gpc1_1 gpc1497 (
      {stage1_11[146]},
      {stage2_11[100]}
   );
   gpc1_1 gpc1498 (
      {stage1_11[147]},
      {stage2_11[101]}
   );
   gpc1_1 gpc1499 (
      {stage1_11[148]},
      {stage2_11[102]}
   );
   gpc1_1 gpc1500 (
      {stage1_11[149]},
      {stage2_11[103]}
   );
   gpc1_1 gpc1501 (
      {stage1_11[150]},
      {stage2_11[104]}
   );
   gpc1_1 gpc1502 (
      {stage1_11[151]},
      {stage2_11[105]}
   );
   gpc1_1 gpc1503 (
      {stage1_11[152]},
      {stage2_11[106]}
   );
   gpc1_1 gpc1504 (
      {stage1_11[153]},
      {stage2_11[107]}
   );
   gpc1_1 gpc1505 (
      {stage1_11[154]},
      {stage2_11[108]}
   );
   gpc1_1 gpc1506 (
      {stage1_11[155]},
      {stage2_11[109]}
   );
   gpc1_1 gpc1507 (
      {stage1_11[156]},
      {stage2_11[110]}
   );
   gpc1_1 gpc1508 (
      {stage1_11[157]},
      {stage2_11[111]}
   );
   gpc1_1 gpc1509 (
      {stage1_11[158]},
      {stage2_11[112]}
   );
   gpc1_1 gpc1510 (
      {stage1_11[159]},
      {stage2_11[113]}
   );
   gpc1_1 gpc1511 (
      {stage1_11[160]},
      {stage2_11[114]}
   );
   gpc1_1 gpc1512 (
      {stage1_11[161]},
      {stage2_11[115]}
   );
   gpc1_1 gpc1513 (
      {stage1_11[162]},
      {stage2_11[116]}
   );
   gpc1_1 gpc1514 (
      {stage1_11[163]},
      {stage2_11[117]}
   );
   gpc1_1 gpc1515 (
      {stage1_11[164]},
      {stage2_11[118]}
   );
   gpc1_1 gpc1516 (
      {stage1_11[165]},
      {stage2_11[119]}
   );
   gpc1_1 gpc1517 (
      {stage1_11[166]},
      {stage2_11[120]}
   );
   gpc1_1 gpc1518 (
      {stage1_11[167]},
      {stage2_11[121]}
   );
   gpc1_1 gpc1519 (
      {stage1_11[168]},
      {stage2_11[122]}
   );
   gpc1_1 gpc1520 (
      {stage1_11[169]},
      {stage2_11[123]}
   );
   gpc1_1 gpc1521 (
      {stage1_11[170]},
      {stage2_11[124]}
   );
   gpc1_1 gpc1522 (
      {stage1_11[171]},
      {stage2_11[125]}
   );
   gpc1_1 gpc1523 (
      {stage1_11[172]},
      {stage2_11[126]}
   );
   gpc1_1 gpc1524 (
      {stage1_11[173]},
      {stage2_11[127]}
   );
   gpc1_1 gpc1525 (
      {stage1_11[174]},
      {stage2_11[128]}
   );
   gpc1_1 gpc1526 (
      {stage1_11[175]},
      {stage2_11[129]}
   );
   gpc1_1 gpc1527 (
      {stage1_11[176]},
      {stage2_11[130]}
   );
   gpc1_1 gpc1528 (
      {stage1_11[177]},
      {stage2_11[131]}
   );
   gpc1_1 gpc1529 (
      {stage1_11[178]},
      {stage2_11[132]}
   );
   gpc1_1 gpc1530 (
      {stage1_11[179]},
      {stage2_11[133]}
   );
   gpc1_1 gpc1531 (
      {stage1_11[180]},
      {stage2_11[134]}
   );
   gpc1_1 gpc1532 (
      {stage1_11[181]},
      {stage2_11[135]}
   );
   gpc1_1 gpc1533 (
      {stage1_11[182]},
      {stage2_11[136]}
   );
   gpc1_1 gpc1534 (
      {stage1_11[183]},
      {stage2_11[137]}
   );
   gpc1_1 gpc1535 (
      {stage1_11[184]},
      {stage2_11[138]}
   );
   gpc1_1 gpc1536 (
      {stage1_11[185]},
      {stage2_11[139]}
   );
   gpc1_1 gpc1537 (
      {stage1_11[186]},
      {stage2_11[140]}
   );
   gpc1_1 gpc1538 (
      {stage1_11[187]},
      {stage2_11[141]}
   );
   gpc1_1 gpc1539 (
      {stage1_11[188]},
      {stage2_11[142]}
   );
   gpc1_1 gpc1540 (
      {stage1_11[189]},
      {stage2_11[143]}
   );
   gpc1_1 gpc1541 (
      {stage1_12[210]},
      {stage2_12[73]}
   );
   gpc1_1 gpc1542 (
      {stage1_12[211]},
      {stage2_12[74]}
   );
   gpc1_1 gpc1543 (
      {stage1_12[212]},
      {stage2_12[75]}
   );
   gpc1_1 gpc1544 (
      {stage1_12[213]},
      {stage2_12[76]}
   );
   gpc1_1 gpc1545 (
      {stage1_12[214]},
      {stage2_12[77]}
   );
   gpc1_1 gpc1546 (
      {stage1_12[215]},
      {stage2_12[78]}
   );
   gpc1_1 gpc1547 (
      {stage1_12[216]},
      {stage2_12[79]}
   );
   gpc1_1 gpc1548 (
      {stage1_12[217]},
      {stage2_12[80]}
   );
   gpc1_1 gpc1549 (
      {stage1_12[218]},
      {stage2_12[81]}
   );
   gpc1_1 gpc1550 (
      {stage1_12[219]},
      {stage2_12[82]}
   );
   gpc1_1 gpc1551 (
      {stage1_12[220]},
      {stage2_12[83]}
   );
   gpc1_1 gpc1552 (
      {stage1_12[221]},
      {stage2_12[84]}
   );
   gpc1_1 gpc1553 (
      {stage1_13[232]},
      {stage2_13[91]}
   );
   gpc1_1 gpc1554 (
      {stage1_13[233]},
      {stage2_13[92]}
   );
   gpc1_1 gpc1555 (
      {stage1_13[234]},
      {stage2_13[93]}
   );
   gpc1_1 gpc1556 (
      {stage1_13[235]},
      {stage2_13[94]}
   );
   gpc1_1 gpc1557 (
      {stage1_13[236]},
      {stage2_13[95]}
   );
   gpc1_1 gpc1558 (
      {stage1_13[237]},
      {stage2_13[96]}
   );
   gpc1_1 gpc1559 (
      {stage1_13[238]},
      {stage2_13[97]}
   );
   gpc1_1 gpc1560 (
      {stage1_13[239]},
      {stage2_13[98]}
   );
   gpc1_1 gpc1561 (
      {stage1_13[240]},
      {stage2_13[99]}
   );
   gpc1_1 gpc1562 (
      {stage1_13[241]},
      {stage2_13[100]}
   );
   gpc1_1 gpc1563 (
      {stage1_13[242]},
      {stage2_13[101]}
   );
   gpc1_1 gpc1564 (
      {stage1_13[243]},
      {stage2_13[102]}
   );
   gpc1_1 gpc1565 (
      {stage1_13[244]},
      {stage2_13[103]}
   );
   gpc1_1 gpc1566 (
      {stage1_13[245]},
      {stage2_13[104]}
   );
   gpc1_1 gpc1567 (
      {stage1_13[246]},
      {stage2_13[105]}
   );
   gpc1_1 gpc1568 (
      {stage1_13[247]},
      {stage2_13[106]}
   );
   gpc1_1 gpc1569 (
      {stage1_13[248]},
      {stage2_13[107]}
   );
   gpc1_1 gpc1570 (
      {stage1_13[249]},
      {stage2_13[108]}
   );
   gpc1_1 gpc1571 (
      {stage1_13[250]},
      {stage2_13[109]}
   );
   gpc1_1 gpc1572 (
      {stage1_13[251]},
      {stage2_13[110]}
   );
   gpc1_1 gpc1573 (
      {stage1_13[252]},
      {stage2_13[111]}
   );
   gpc1_1 gpc1574 (
      {stage1_13[253]},
      {stage2_13[112]}
   );
   gpc1_1 gpc1575 (
      {stage1_13[254]},
      {stage2_13[113]}
   );
   gpc1_1 gpc1576 (
      {stage1_13[255]},
      {stage2_13[114]}
   );
   gpc1_1 gpc1577 (
      {stage1_13[256]},
      {stage2_13[115]}
   );
   gpc1_1 gpc1578 (
      {stage1_13[257]},
      {stage2_13[116]}
   );
   gpc1_1 gpc1579 (
      {stage1_13[258]},
      {stage2_13[117]}
   );
   gpc1_1 gpc1580 (
      {stage1_13[259]},
      {stage2_13[118]}
   );
   gpc1_1 gpc1581 (
      {stage1_13[260]},
      {stage2_13[119]}
   );
   gpc1_1 gpc1582 (
      {stage1_13[261]},
      {stage2_13[120]}
   );
   gpc1_1 gpc1583 (
      {stage1_13[262]},
      {stage2_13[121]}
   );
   gpc1_1 gpc1584 (
      {stage1_13[263]},
      {stage2_13[122]}
   );
   gpc1_1 gpc1585 (
      {stage1_13[264]},
      {stage2_13[123]}
   );
   gpc1_1 gpc1586 (
      {stage1_13[265]},
      {stage2_13[124]}
   );
   gpc1_1 gpc1587 (
      {stage1_13[266]},
      {stage2_13[125]}
   );
   gpc1_1 gpc1588 (
      {stage1_13[267]},
      {stage2_13[126]}
   );
   gpc1_1 gpc1589 (
      {stage1_13[268]},
      {stage2_13[127]}
   );
   gpc1_1 gpc1590 (
      {stage1_13[269]},
      {stage2_13[128]}
   );
   gpc1_1 gpc1591 (
      {stage1_13[270]},
      {stage2_13[129]}
   );
   gpc1_1 gpc1592 (
      {stage1_13[271]},
      {stage2_13[130]}
   );
   gpc1_1 gpc1593 (
      {stage1_13[272]},
      {stage2_13[131]}
   );
   gpc1_1 gpc1594 (
      {stage1_13[273]},
      {stage2_13[132]}
   );
   gpc1_1 gpc1595 (
      {stage1_13[274]},
      {stage2_13[133]}
   );
   gpc1_1 gpc1596 (
      {stage1_13[275]},
      {stage2_13[134]}
   );
   gpc1_1 gpc1597 (
      {stage1_13[276]},
      {stage2_13[135]}
   );
   gpc1_1 gpc1598 (
      {stage1_13[277]},
      {stage2_13[136]}
   );
   gpc1_1 gpc1599 (
      {stage1_13[278]},
      {stage2_13[137]}
   );
   gpc1_1 gpc1600 (
      {stage1_13[279]},
      {stage2_13[138]}
   );
   gpc1_1 gpc1601 (
      {stage1_13[280]},
      {stage2_13[139]}
   );
   gpc1_1 gpc1602 (
      {stage1_13[281]},
      {stage2_13[140]}
   );
   gpc1_1 gpc1603 (
      {stage1_14[211]},
      {stage2_14[91]}
   );
   gpc1_1 gpc1604 (
      {stage1_14[212]},
      {stage2_14[92]}
   );
   gpc1_1 gpc1605 (
      {stage1_14[213]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1606 (
      {stage1_14[214]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1607 (
      {stage1_14[215]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1608 (
      {stage1_14[216]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1609 (
      {stage1_14[217]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1610 (
      {stage1_14[218]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1611 (
      {stage1_14[219]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1612 (
      {stage1_14[220]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1613 (
      {stage1_14[221]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1614 (
      {stage1_14[222]},
      {stage2_14[102]}
   );
   gpc1_1 gpc1615 (
      {stage1_14[223]},
      {stage2_14[103]}
   );
   gpc1_1 gpc1616 (
      {stage1_14[224]},
      {stage2_14[104]}
   );
   gpc1_1 gpc1617 (
      {stage1_14[225]},
      {stage2_14[105]}
   );
   gpc1_1 gpc1618 (
      {stage1_14[226]},
      {stage2_14[106]}
   );
   gpc1_1 gpc1619 (
      {stage1_14[227]},
      {stage2_14[107]}
   );
   gpc1_1 gpc1620 (
      {stage1_14[228]},
      {stage2_14[108]}
   );
   gpc1_1 gpc1621 (
      {stage1_14[229]},
      {stage2_14[109]}
   );
   gpc1_1 gpc1622 (
      {stage1_14[230]},
      {stage2_14[110]}
   );
   gpc1_1 gpc1623 (
      {stage1_14[231]},
      {stage2_14[111]}
   );
   gpc1_1 gpc1624 (
      {stage1_14[232]},
      {stage2_14[112]}
   );
   gpc1_1 gpc1625 (
      {stage1_14[233]},
      {stage2_14[113]}
   );
   gpc1_1 gpc1626 (
      {stage1_14[234]},
      {stage2_14[114]}
   );
   gpc1_1 gpc1627 (
      {stage1_14[235]},
      {stage2_14[115]}
   );
   gpc1_1 gpc1628 (
      {stage1_14[236]},
      {stage2_14[116]}
   );
   gpc1_1 gpc1629 (
      {stage1_14[237]},
      {stage2_14[117]}
   );
   gpc1_1 gpc1630 (
      {stage1_14[238]},
      {stage2_14[118]}
   );
   gpc1_1 gpc1631 (
      {stage1_14[239]},
      {stage2_14[119]}
   );
   gpc1_1 gpc1632 (
      {stage1_14[240]},
      {stage2_14[120]}
   );
   gpc1_1 gpc1633 (
      {stage1_14[241]},
      {stage2_14[121]}
   );
   gpc1_1 gpc1634 (
      {stage1_14[242]},
      {stage2_14[122]}
   );
   gpc1_1 gpc1635 (
      {stage1_14[243]},
      {stage2_14[123]}
   );
   gpc1_1 gpc1636 (
      {stage1_14[244]},
      {stage2_14[124]}
   );
   gpc1_1 gpc1637 (
      {stage1_16[101]},
      {stage2_16[79]}
   );
   gpc1_1 gpc1638 (
      {stage1_16[102]},
      {stage2_16[80]}
   );
   gpc1_1 gpc1639 (
      {stage1_16[103]},
      {stage2_16[81]}
   );
   gpc1_1 gpc1640 (
      {stage1_16[104]},
      {stage2_16[82]}
   );
   gpc1_1 gpc1641 (
      {stage1_16[105]},
      {stage2_16[83]}
   );
   gpc1_1 gpc1642 (
      {stage1_16[106]},
      {stage2_16[84]}
   );
   gpc1_1 gpc1643 (
      {stage1_16[107]},
      {stage2_16[85]}
   );
   gpc1_1 gpc1644 (
      {stage1_16[108]},
      {stage2_16[86]}
   );
   gpc1_1 gpc1645 (
      {stage1_16[109]},
      {stage2_16[87]}
   );
   gpc1_1 gpc1646 (
      {stage1_16[110]},
      {stage2_16[88]}
   );
   gpc1_1 gpc1647 (
      {stage1_16[111]},
      {stage2_16[89]}
   );
   gpc1_1 gpc1648 (
      {stage1_16[112]},
      {stage2_16[90]}
   );
   gpc1_1 gpc1649 (
      {stage1_16[113]},
      {stage2_16[91]}
   );
   gpc1_1 gpc1650 (
      {stage1_16[114]},
      {stage2_16[92]}
   );
   gpc1_1 gpc1651 (
      {stage1_16[115]},
      {stage2_16[93]}
   );
   gpc1_1 gpc1652 (
      {stage1_16[116]},
      {stage2_16[94]}
   );
   gpc1_1 gpc1653 (
      {stage1_16[117]},
      {stage2_16[95]}
   );
   gpc1_1 gpc1654 (
      {stage1_16[118]},
      {stage2_16[96]}
   );
   gpc1_1 gpc1655 (
      {stage1_16[119]},
      {stage2_16[97]}
   );
   gpc1_1 gpc1656 (
      {stage1_16[120]},
      {stage2_16[98]}
   );
   gpc1_1 gpc1657 (
      {stage1_16[121]},
      {stage2_16[99]}
   );
   gpc1_1 gpc1658 (
      {stage1_16[122]},
      {stage2_16[100]}
   );
   gpc1_1 gpc1659 (
      {stage1_16[123]},
      {stage2_16[101]}
   );
   gpc1_1 gpc1660 (
      {stage1_16[124]},
      {stage2_16[102]}
   );
   gpc1_1 gpc1661 (
      {stage1_16[125]},
      {stage2_16[103]}
   );
   gpc1_1 gpc1662 (
      {stage1_16[126]},
      {stage2_16[104]}
   );
   gpc606_5 gpc1663 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc1664 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_1[0]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc1665 (
      {stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15]},
      {stage2_1[1]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc1666 (
      {stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[2]},
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1667 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc1668 (
      {stage2_1[9], stage2_1[10], stage2_1[11], stage2_1[12], stage2_1[13], stage2_1[14]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc1669 (
      {stage2_1[15], stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1670 (
      {stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24], stage2_1[25], stage2_1[26]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1671 (
      {stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30], stage2_1[31], stage2_1[32]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1672 (
      {stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36], stage2_1[37], stage2_1[38]},
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1673 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc1674 (
      {stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[36]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc1675 (
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38], stage2_2[39]},
      {stage2_3[37]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc1676 (
      {stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_3[38]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc1677 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49]},
      {stage2_3[39]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1678 (
      {stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage2_3[40]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1679 (
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59]},
      {stage2_3[41]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc606_5 gpc1680 (
      {stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc1681 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52]},
      {stage2_4[42]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc1682 (
      {stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57]},
      {stage2_4[43]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1683 (
      {stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62]},
      {stage2_4[44]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1684 (
      {stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67]},
      {stage2_4[45]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1685 (
      {stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage2_4[46]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1686 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[47]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc1687 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[48]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc1688 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[49]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc1689 (
      {stage2_3[88], stage2_3[89], stage2_3[90], stage2_3[91], stage2_3[92]},
      {stage2_4[50]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc1690 (
      {stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96], stage2_3[97]},
      {stage2_4[51]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc1691 (
      {stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102]},
      {stage2_4[52]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc1692 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc1693 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc1694 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[14],stage3_6[21],stage3_5[27],stage3_4[31]}
   );
   gpc606_5 gpc1695 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[15],stage3_6[22],stage3_5[28],stage3_4[32]}
   );
   gpc606_5 gpc1696 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[16],stage3_6[23],stage3_5[29],stage3_4[33]}
   );
   gpc606_5 gpc1697 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[17],stage3_6[24],stage3_5[30],stage3_4[34]}
   );
   gpc606_5 gpc1698 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[18],stage3_6[25],stage3_5[31],stage3_4[35]}
   );
   gpc606_5 gpc1699 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[19],stage3_6[26],stage3_5[32],stage3_4[36]}
   );
   gpc606_5 gpc1700 (
      {stage2_4[101], stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[20],stage3_6[27],stage3_5[33],stage3_4[37]}
   );
   gpc615_5 gpc1701 (
      {stage2_4[107], stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111]},
      {stage2_5[72]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[21],stage3_6[28],stage3_5[34],stage3_4[38]}
   );
   gpc615_5 gpc1702 (
      {stage2_4[112], stage2_4[113], stage2_4[114], stage2_4[115], stage2_4[116]},
      {stage2_5[73]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[22],stage3_6[29],stage3_5[35],stage3_4[39]}
   );
   gpc615_5 gpc1703 (
      {stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77], stage2_5[78]},
      {stage2_6[66]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[11],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc615_5 gpc1704 (
      {stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_6[67]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[12],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1705 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[13],stage3_7[25],stage3_6[32]}
   );
   gpc606_5 gpc1706 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78], stage2_6[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[14],stage3_7[26],stage3_6[33]}
   );
   gpc606_5 gpc1707 (
      {stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83], stage2_6[84], stage2_6[85]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[15],stage3_7[27],stage3_6[34]}
   );
   gpc606_5 gpc1708 (
      {stage2_6[86], stage2_6[87], stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[5],stage3_8[16],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc1709 (
      {stage2_6[92], stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[6],stage3_8[17],stage3_7[29],stage3_6[36]}
   );
   gpc606_5 gpc1710 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102], stage2_6[103]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[7],stage3_8[18],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1711 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[8],stage3_8[19],stage3_7[31]}
   );
   gpc615_5 gpc1712 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[9],stage3_8[20],stage3_7[32]}
   );
   gpc615_5 gpc1713 (
      {stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[10],stage3_8[21],stage3_7[33]}
   );
   gpc615_5 gpc1714 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[11],stage3_8[22],stage3_7[34]}
   );
   gpc615_5 gpc1715 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[40]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[10],stage3_9[12],stage3_8[23],stage3_7[35]}
   );
   gpc615_5 gpc1716 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[41]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[11],stage3_9[13],stage3_8[24],stage3_7[36]}
   );
   gpc615_5 gpc1717 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[42]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[12],stage3_9[14],stage3_8[25],stage3_7[37]}
   );
   gpc615_5 gpc1718 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[43]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[13],stage3_9[15],stage3_8[26],stage3_7[38]}
   );
   gpc615_5 gpc1719 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[44]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[14],stage3_9[16],stage3_8[27],stage3_7[39]}
   );
   gpc615_5 gpc1720 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[45]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[15],stage3_9[17],stage3_8[28],stage3_7[40]}
   );
   gpc615_5 gpc1721 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[46]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[16],stage3_9[18],stage3_8[29],stage3_7[41]}
   );
   gpc615_5 gpc1722 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[47]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[17],stage3_9[19],stage3_8[30],stage3_7[42]}
   );
   gpc615_5 gpc1723 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[48]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[18],stage3_9[20],stage3_8[31],stage3_7[43]}
   );
   gpc615_5 gpc1724 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[49]},
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage3_11[13],stage3_10[19],stage3_9[21],stage3_8[32],stage3_7[44]}
   );
   gpc615_5 gpc1725 (
      {stage2_7[82], stage2_7[83], stage2_7[84], 1'b0, 1'b0},
      {stage2_8[50]},
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage3_11[14],stage3_10[20],stage3_9[22],stage3_8[33],stage3_7[45]}
   );
   gpc606_5 gpc1726 (
      {stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[15],stage3_10[21],stage3_9[23],stage3_8[34]}
   );
   gpc615_5 gpc1727 (
      {stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61]},
      {stage2_9[90]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[16],stage3_10[22],stage3_9[24],stage3_8[35]}
   );
   gpc615_5 gpc1728 (
      {stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65], stage2_8[66]},
      {stage2_9[91]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[17],stage3_10[23],stage3_9[25],stage3_8[36]}
   );
   gpc615_5 gpc1729 (
      {stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_9[92]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[18],stage3_10[24],stage3_9[26],stage3_8[37]}
   );
   gpc615_5 gpc1730 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_9[93]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[19],stage3_10[25],stage3_9[27],stage3_8[38]}
   );
   gpc615_5 gpc1731 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_9[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[20],stage3_10[26],stage3_9[28],stage3_8[39]}
   );
   gpc615_5 gpc1732 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86]},
      {stage2_9[95]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[21],stage3_10[27],stage3_9[29],stage3_8[40]}
   );
   gpc606_5 gpc1733 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[22],stage3_10[28],stage3_9[30]}
   );
   gpc606_5 gpc1734 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[8],stage3_11[23],stage3_10[29],stage3_9[31]}
   );
   gpc606_5 gpc1735 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[9],stage3_11[24],stage3_10[30],stage3_9[32]}
   );
   gpc606_5 gpc1736 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[10],stage3_11[25],stage3_10[31],stage3_9[33]}
   );
   gpc615_5 gpc1737 (
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[11],stage3_11[26],stage3_10[32]}
   );
   gpc615_5 gpc1738 (
      {stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51]},
      {stage2_11[25]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[5],stage3_12[12],stage3_11[27],stage3_10[33]}
   );
   gpc615_5 gpc1739 (
      {stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_11[26]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[6],stage3_12[13],stage3_11[28],stage3_10[34]}
   );
   gpc606_5 gpc1740 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[7],stage3_12[14],stage3_11[29]}
   );
   gpc606_5 gpc1741 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[8],stage3_12[15],stage3_11[30]}
   );
   gpc606_5 gpc1742 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[9],stage3_12[16],stage3_11[31]}
   );
   gpc606_5 gpc1743 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[10],stage3_12[17],stage3_11[32]}
   );
   gpc606_5 gpc1744 (
      {stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[11],stage3_12[18],stage3_11[33]}
   );
   gpc606_5 gpc1745 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[12],stage3_12[19],stage3_11[34]}
   );
   gpc606_5 gpc1746 (
      {stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[9],stage3_13[13],stage3_12[20],stage3_11[35]}
   );
   gpc606_5 gpc1747 (
      {stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[10],stage3_13[14],stage3_12[21],stage3_11[36]}
   );
   gpc606_5 gpc1748 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[11],stage3_13[15],stage3_12[22],stage3_11[37]}
   );
   gpc606_5 gpc1749 (
      {stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[12],stage3_13[16],stage3_12[23],stage3_11[38]}
   );
   gpc606_5 gpc1750 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91], stage2_11[92]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[13],stage3_13[17],stage3_12[24],stage3_11[39]}
   );
   gpc606_5 gpc1751 (
      {stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[14],stage3_13[18],stage3_12[25],stage3_11[40]}
   );
   gpc606_5 gpc1752 (
      {stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[15],stage3_13[19],stage3_12[26],stage3_11[41]}
   );
   gpc606_5 gpc1753 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109], stage2_11[110]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[16],stage3_13[20],stage3_12[27],stage3_11[42]}
   );
   gpc606_5 gpc1754 (
      {stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114], stage2_11[115], stage2_11[116]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[17],stage3_13[21],stage3_12[28],stage3_11[43]}
   );
   gpc606_5 gpc1755 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121], stage2_11[122]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[18],stage3_13[22],stage3_12[29],stage3_11[44]}
   );
   gpc606_5 gpc1756 (
      {stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126], stage2_11[127], stage2_11[128]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[19],stage3_13[23],stage3_12[30],stage3_11[45]}
   );
   gpc606_5 gpc1757 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[17],stage3_14[20],stage3_13[24],stage3_12[31]}
   );
   gpc606_5 gpc1758 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[18],stage3_14[21],stage3_13[25],stage3_12[32]}
   );
   gpc606_5 gpc1759 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[19],stage3_14[22],stage3_13[26],stage3_12[33]}
   );
   gpc606_5 gpc1760 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[20],stage3_14[23],stage3_13[27],stage3_12[34]}
   );
   gpc606_5 gpc1761 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[21],stage3_14[24],stage3_13[28],stage3_12[35]}
   );
   gpc606_5 gpc1762 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[22],stage3_14[25],stage3_13[29],stage3_12[36]}
   );
   gpc606_5 gpc1763 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[23],stage3_14[26],stage3_13[30],stage3_12[37]}
   );
   gpc606_5 gpc1764 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[24],stage3_14[27],stage3_13[31],stage3_12[38]}
   );
   gpc606_5 gpc1765 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[25],stage3_14[28],stage3_13[32],stage3_12[39]}
   );
   gpc606_5 gpc1766 (
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[9],stage3_15[26],stage3_14[29],stage3_13[33]}
   );
   gpc606_5 gpc1767 (
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[10],stage3_15[27],stage3_14[30],stage3_13[34]}
   );
   gpc606_5 gpc1768 (
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[11],stage3_15[28],stage3_14[31],stage3_13[35]}
   );
   gpc606_5 gpc1769 (
      {stage2_13[120], stage2_13[121], stage2_13[122], stage2_13[123], stage2_13[124], stage2_13[125]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[12],stage3_15[29],stage3_14[32],stage3_13[36]}
   );
   gpc606_5 gpc1770 (
      {stage2_13[126], stage2_13[127], stage2_13[128], stage2_13[129], stage2_13[130], stage2_13[131]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[13],stage3_15[30],stage3_14[33],stage3_13[37]}
   );
   gpc606_5 gpc1771 (
      {stage2_13[132], stage2_13[133], stage2_13[134], stage2_13[135], stage2_13[136], stage2_13[137]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[14],stage3_15[31],stage3_14[34],stage3_13[38]}
   );
   gpc606_5 gpc1772 (
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[15],stage3_15[32],stage3_14[35]}
   );
   gpc606_5 gpc1773 (
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[16],stage3_15[33],stage3_14[36]}
   );
   gpc606_5 gpc1774 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[17],stage3_15[34],stage3_14[37]}
   );
   gpc606_5 gpc1775 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[18],stage3_15[35],stage3_14[38]}
   );
   gpc606_5 gpc1776 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[19],stage3_15[36],stage3_14[39]}
   );
   gpc606_5 gpc1777 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[20],stage3_15[37],stage3_14[40]}
   );
   gpc606_5 gpc1778 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[21],stage3_15[38],stage3_14[41]}
   );
   gpc606_5 gpc1779 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[13],stage3_16[22],stage3_15[39],stage3_14[42]}
   );
   gpc615_5 gpc1780 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106]},
      {stage2_15[36]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[14],stage3_16[23],stage3_15[40],stage3_14[43]}
   );
   gpc615_5 gpc1781 (
      {stage2_14[107], stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111]},
      {stage2_15[37]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[15],stage3_16[24],stage3_15[41],stage3_14[44]}
   );
   gpc615_5 gpc1782 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[16],stage3_16[25],stage3_15[42]}
   );
   gpc615_5 gpc1783 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[17],stage3_16[26],stage3_15[43]}
   );
   gpc615_5 gpc1784 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[18],stage3_16[27],stage3_15[44]}
   );
   gpc615_5 gpc1785 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[19],stage3_16[28],stage3_15[45]}
   );
   gpc615_5 gpc1786 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[20],stage3_16[29],stage3_15[46]}
   );
   gpc615_5 gpc1787 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[21],stage3_16[30],stage3_15[47]}
   );
   gpc615_5 gpc1788 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[22],stage3_16[31],stage3_15[48]}
   );
   gpc615_5 gpc1789 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[23],stage3_16[32],stage3_15[49]}
   );
   gpc606_5 gpc1790 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[18],stage3_17[24],stage3_16[33]}
   );
   gpc606_5 gpc1791 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[9],stage3_18[19],stage3_17[25],stage3_16[34]}
   );
   gpc606_5 gpc1792 (
      {stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83], stage2_16[84], stage2_16[85]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[10],stage3_18[20],stage3_17[26],stage3_16[35]}
   );
   gpc606_5 gpc1793 (
      {stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89], stage2_16[90], stage2_16[91]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[11],stage3_18[21],stage3_17[27],stage3_16[36]}
   );
   gpc606_5 gpc1794 (
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[4],stage3_19[12],stage3_18[22],stage3_17[28]}
   );
   gpc606_5 gpc1795 (
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], 1'b0},
      {stage3_21[1],stage3_20[5],stage3_19[13],stage3_18[23],stage3_17[29]}
   );
   gpc1_1 gpc1796 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1797 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1798 (
      {stage2_1[39]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1799 (
      {stage2_1[40]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1800 (
      {stage2_5[84]},
      {stage3_5[38]}
   );
   gpc1_1 gpc1801 (
      {stage2_5[85]},
      {stage3_5[39]}
   );
   gpc1_1 gpc1802 (
      {stage2_5[86]},
      {stage3_5[40]}
   );
   gpc1_1 gpc1803 (
      {stage2_5[87]},
      {stage3_5[41]}
   );
   gpc1_1 gpc1804 (
      {stage2_5[88]},
      {stage3_5[42]}
   );
   gpc1_1 gpc1805 (
      {stage2_5[89]},
      {stage3_5[43]}
   );
   gpc1_1 gpc1806 (
      {stage2_5[90]},
      {stage3_5[44]}
   );
   gpc1_1 gpc1807 (
      {stage2_5[91]},
      {stage3_5[45]}
   );
   gpc1_1 gpc1808 (
      {stage2_5[92]},
      {stage3_5[46]}
   );
   gpc1_1 gpc1809 (
      {stage2_5[93]},
      {stage3_5[47]}
   );
   gpc1_1 gpc1810 (
      {stage2_9[120]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_9[121]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_9[122]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_9[123]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_9[124]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_9[125]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_9[126]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1817 (
      {stage2_9[127]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1818 (
      {stage2_9[128]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1819 (
      {stage2_9[129]},
      {stage3_9[43]}
   );
   gpc1_1 gpc1820 (
      {stage2_9[130]},
      {stage3_9[44]}
   );
   gpc1_1 gpc1821 (
      {stage2_9[131]},
      {stage3_9[45]}
   );
   gpc1_1 gpc1822 (
      {stage2_9[132]},
      {stage3_9[46]}
   );
   gpc1_1 gpc1823 (
      {stage2_9[133]},
      {stage3_9[47]}
   );
   gpc1_1 gpc1824 (
      {stage2_9[134]},
      {stage3_9[48]}
   );
   gpc1_1 gpc1825 (
      {stage2_9[135]},
      {stage3_9[49]}
   );
   gpc1_1 gpc1826 (
      {stage2_9[136]},
      {stage3_9[50]}
   );
   gpc1_1 gpc1827 (
      {stage2_9[137]},
      {stage3_9[51]}
   );
   gpc1_1 gpc1828 (
      {stage2_10[57]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1829 (
      {stage2_10[58]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1830 (
      {stage2_10[59]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1831 (
      {stage2_10[60]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1832 (
      {stage2_10[61]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1833 (
      {stage2_10[62]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1834 (
      {stage2_10[63]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1835 (
      {stage2_10[64]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1836 (
      {stage2_10[65]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1837 (
      {stage2_10[66]},
      {stage3_10[44]}
   );
   gpc1_1 gpc1838 (
      {stage2_10[67]},
      {stage3_10[45]}
   );
   gpc1_1 gpc1839 (
      {stage2_10[68]},
      {stage3_10[46]}
   );
   gpc1_1 gpc1840 (
      {stage2_10[69]},
      {stage3_10[47]}
   );
   gpc1_1 gpc1841 (
      {stage2_10[70]},
      {stage3_10[48]}
   );
   gpc1_1 gpc1842 (
      {stage2_10[71]},
      {stage3_10[49]}
   );
   gpc1_1 gpc1843 (
      {stage2_10[72]},
      {stage3_10[50]}
   );
   gpc1_1 gpc1844 (
      {stage2_10[73]},
      {stage3_10[51]}
   );
   gpc1_1 gpc1845 (
      {stage2_10[74]},
      {stage3_10[52]}
   );
   gpc1_1 gpc1846 (
      {stage2_10[75]},
      {stage3_10[53]}
   );
   gpc1_1 gpc1847 (
      {stage2_10[76]},
      {stage3_10[54]}
   );
   gpc1_1 gpc1848 (
      {stage2_10[77]},
      {stage3_10[55]}
   );
   gpc1_1 gpc1849 (
      {stage2_10[78]},
      {stage3_10[56]}
   );
   gpc1_1 gpc1850 (
      {stage2_10[79]},
      {stage3_10[57]}
   );
   gpc1_1 gpc1851 (
      {stage2_10[80]},
      {stage3_10[58]}
   );
   gpc1_1 gpc1852 (
      {stage2_10[81]},
      {stage3_10[59]}
   );
   gpc1_1 gpc1853 (
      {stage2_10[82]},
      {stage3_10[60]}
   );
   gpc1_1 gpc1854 (
      {stage2_10[83]},
      {stage3_10[61]}
   );
   gpc1_1 gpc1855 (
      {stage2_10[84]},
      {stage3_10[62]}
   );
   gpc1_1 gpc1856 (
      {stage2_10[85]},
      {stage3_10[63]}
   );
   gpc1_1 gpc1857 (
      {stage2_11[129]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1858 (
      {stage2_11[130]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1859 (
      {stage2_11[131]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1860 (
      {stage2_11[132]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1861 (
      {stage2_11[133]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1862 (
      {stage2_11[134]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1863 (
      {stage2_11[135]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1864 (
      {stage2_11[136]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1865 (
      {stage2_11[137]},
      {stage3_11[54]}
   );
   gpc1_1 gpc1866 (
      {stage2_11[138]},
      {stage3_11[55]}
   );
   gpc1_1 gpc1867 (
      {stage2_11[139]},
      {stage3_11[56]}
   );
   gpc1_1 gpc1868 (
      {stage2_11[140]},
      {stage3_11[57]}
   );
   gpc1_1 gpc1869 (
      {stage2_11[141]},
      {stage3_11[58]}
   );
   gpc1_1 gpc1870 (
      {stage2_11[142]},
      {stage3_11[59]}
   );
   gpc1_1 gpc1871 (
      {stage2_11[143]},
      {stage3_11[60]}
   );
   gpc1_1 gpc1872 (
      {stage2_12[72]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1873 (
      {stage2_12[73]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1874 (
      {stage2_12[74]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1875 (
      {stage2_12[75]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1876 (
      {stage2_12[76]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1877 (
      {stage2_12[77]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1878 (
      {stage2_12[78]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1879 (
      {stage2_12[79]},
      {stage3_12[47]}
   );
   gpc1_1 gpc1880 (
      {stage2_12[80]},
      {stage3_12[48]}
   );
   gpc1_1 gpc1881 (
      {stage2_12[81]},
      {stage3_12[49]}
   );
   gpc1_1 gpc1882 (
      {stage2_12[82]},
      {stage3_12[50]}
   );
   gpc1_1 gpc1883 (
      {stage2_12[83]},
      {stage3_12[51]}
   );
   gpc1_1 gpc1884 (
      {stage2_12[84]},
      {stage3_12[52]}
   );
   gpc1_1 gpc1885 (
      {stage2_13[138]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1886 (
      {stage2_13[139]},
      {stage3_13[40]}
   );
   gpc1_1 gpc1887 (
      {stage2_13[140]},
      {stage3_13[41]}
   );
   gpc1_1 gpc1888 (
      {stage2_14[112]},
      {stage3_14[45]}
   );
   gpc1_1 gpc1889 (
      {stage2_14[113]},
      {stage3_14[46]}
   );
   gpc1_1 gpc1890 (
      {stage2_14[114]},
      {stage3_14[47]}
   );
   gpc1_1 gpc1891 (
      {stage2_14[115]},
      {stage3_14[48]}
   );
   gpc1_1 gpc1892 (
      {stage2_14[116]},
      {stage3_14[49]}
   );
   gpc1_1 gpc1893 (
      {stage2_14[117]},
      {stage3_14[50]}
   );
   gpc1_1 gpc1894 (
      {stage2_14[118]},
      {stage3_14[51]}
   );
   gpc1_1 gpc1895 (
      {stage2_14[119]},
      {stage3_14[52]}
   );
   gpc1_1 gpc1896 (
      {stage2_14[120]},
      {stage3_14[53]}
   );
   gpc1_1 gpc1897 (
      {stage2_14[121]},
      {stage3_14[54]}
   );
   gpc1_1 gpc1898 (
      {stage2_14[122]},
      {stage3_14[55]}
   );
   gpc1_1 gpc1899 (
      {stage2_14[123]},
      {stage3_14[56]}
   );
   gpc1_1 gpc1900 (
      {stage2_14[124]},
      {stage3_14[57]}
   );
   gpc1_1 gpc1901 (
      {stage2_15[78]},
      {stage3_15[50]}
   );
   gpc1_1 gpc1902 (
      {stage2_15[79]},
      {stage3_15[51]}
   );
   gpc1_1 gpc1903 (
      {stage2_15[80]},
      {stage3_15[52]}
   );
   gpc1_1 gpc1904 (
      {stage2_15[81]},
      {stage3_15[53]}
   );
   gpc1_1 gpc1905 (
      {stage2_15[82]},
      {stage3_15[54]}
   );
   gpc1_1 gpc1906 (
      {stage2_15[83]},
      {stage3_15[55]}
   );
   gpc1_1 gpc1907 (
      {stage2_15[84]},
      {stage3_15[56]}
   );
   gpc1_1 gpc1908 (
      {stage2_16[92]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1909 (
      {stage2_16[93]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1910 (
      {stage2_16[94]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1911 (
      {stage2_16[95]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1912 (
      {stage2_16[96]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1913 (
      {stage2_16[97]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1914 (
      {stage2_16[98]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1915 (
      {stage2_16[99]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1916 (
      {stage2_16[100]},
      {stage3_16[45]}
   );
   gpc1_1 gpc1917 (
      {stage2_16[101]},
      {stage3_16[46]}
   );
   gpc1_1 gpc1918 (
      {stage2_16[102]},
      {stage3_16[47]}
   );
   gpc1_1 gpc1919 (
      {stage2_16[103]},
      {stage3_16[48]}
   );
   gpc1_1 gpc1920 (
      {stage2_16[104]},
      {stage3_16[49]}
   );
   gpc1_1 gpc1921 (
      {stage2_17[60]},
      {stage3_17[30]}
   );
   gpc1_1 gpc1922 (
      {stage2_17[61]},
      {stage3_17[31]}
   );
   gpc1_1 gpc1923 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1924 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc606_5 gpc1925 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc1926 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1927 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[12]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc615_5 gpc1928 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[13]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc615_5 gpc1929 (
      {stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17], stage3_3[18]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc1930 (
      {stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5]}
   );
   gpc606_5 gpc1931 (
      {stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[4],stage4_5[6],stage4_4[6]}
   );
   gpc615_5 gpc1932 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16]},
      {stage3_6[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[5],stage4_5[7]}
   );
   gpc615_5 gpc1933 (
      {stage3_5[17], stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21]},
      {stage3_6[7]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[6],stage4_5[8]}
   );
   gpc615_5 gpc1934 (
      {stage3_5[22], stage3_5[23], stage3_5[24], stage3_5[25], stage3_5[26]},
      {stage3_6[8]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[7],stage4_5[9]}
   );
   gpc615_5 gpc1935 (
      {stage3_5[27], stage3_5[28], stage3_5[29], stage3_5[30], stage3_5[31]},
      {stage3_6[9]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc1936 (
      {stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35], stage3_5[36]},
      {stage3_6[10]},
      {stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage4_9[4],stage4_8[5],stage4_7[7],stage4_6[9],stage4_5[11]}
   );
   gpc615_5 gpc1937 (
      {stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[11]},
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35]},
      {stage4_9[5],stage4_8[6],stage4_7[8],stage4_6[10],stage4_5[12]}
   );
   gpc615_5 gpc1938 (
      {stage3_5[42], stage3_5[43], stage3_5[44], stage3_5[45], stage3_5[46]},
      {stage3_6[12]},
      {stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41]},
      {stage4_9[6],stage4_8[7],stage4_7[9],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc1939 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[7],stage4_8[8],stage4_7[10],stage4_6[12]}
   );
   gpc606_5 gpc1940 (
      {stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[8],stage4_8[9],stage4_7[11],stage4_6[13]}
   );
   gpc606_5 gpc1941 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29], stage3_6[30]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[9],stage4_8[10],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1942 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[10],stage4_8[11]}
   );
   gpc615_5 gpc1943 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[11],stage4_8[12]}
   );
   gpc606_5 gpc1944 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[12]}
   );
   gpc615_5 gpc1945 (
      {stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12]},
      {stage3_10[12]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[13]}
   );
   gpc615_5 gpc1946 (
      {stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_10[13]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[4],stage4_10[7],stage4_9[14]}
   );
   gpc615_5 gpc1947 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22]},
      {stage3_10[14]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[5],stage4_11[5],stage4_10[8],stage4_9[15]}
   );
   gpc615_5 gpc1948 (
      {stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[6],stage4_11[6],stage4_10[9],stage4_9[16]}
   );
   gpc615_5 gpc1949 (
      {stage3_9[28], stage3_9[29], stage3_9[30], stage3_9[31], stage3_9[32]},
      {stage3_10[16]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[7],stage4_11[7],stage4_10[10],stage4_9[17]}
   );
   gpc615_5 gpc1950 (
      {stage3_9[33], stage3_9[34], stage3_9[35], stage3_9[36], stage3_9[37]},
      {stage3_10[17]},
      {stage3_11[36], stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage4_13[6],stage4_12[8],stage4_11[8],stage4_10[11],stage4_9[18]}
   );
   gpc615_5 gpc1951 (
      {stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41], stage3_9[42]},
      {stage3_10[18]},
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage4_13[7],stage4_12[9],stage4_11[9],stage4_10[12],stage4_9[19]}
   );
   gpc615_5 gpc1952 (
      {stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_10[19]},
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52], stage3_11[53]},
      {stage4_13[8],stage4_12[10],stage4_11[10],stage4_10[13],stage4_9[20]}
   );
   gpc606_5 gpc1953 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[9],stage4_12[11],stage4_11[11],stage4_10[14]}
   );
   gpc606_5 gpc1954 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[10],stage4_12[12],stage4_11[12],stage4_10[15]}
   );
   gpc606_5 gpc1955 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[11],stage4_12[13],stage4_11[13],stage4_10[16]}
   );
   gpc606_5 gpc1956 (
      {stage3_10[38], stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[12],stage4_12[14],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1957 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[4],stage4_13[13],stage4_12[15]}
   );
   gpc606_5 gpc1958 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[5],stage4_13[14],stage4_12[16]}
   );
   gpc606_5 gpc1959 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[2],stage4_14[6],stage4_13[15],stage4_12[17]}
   );
   gpc606_5 gpc1960 (
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[3],stage4_14[7],stage4_13[16],stage4_12[18]}
   );
   gpc1163_5 gpc1961 (
      {stage3_13[0], stage3_13[1], stage3_13[2]},
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[0]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[4],stage4_15[4],stage4_14[8],stage4_13[17]}
   );
   gpc1163_5 gpc1962 (
      {stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[30], stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[1]},
      {stage3_16[1]},
      {stage4_17[1],stage4_16[5],stage4_15[5],stage4_14[9],stage4_13[18]}
   );
   gpc1163_5 gpc1963 (
      {stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[36], stage3_14[37], stage3_14[38], stage3_14[39], stage3_14[40], stage3_14[41]},
      {stage3_15[2]},
      {stage3_16[2]},
      {stage4_17[2],stage4_16[6],stage4_15[6],stage4_14[10],stage4_13[19]}
   );
   gpc1163_5 gpc1964 (
      {stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_14[42], stage3_14[43], stage3_14[44], stage3_14[45], stage3_14[46], stage3_14[47]},
      {stage3_15[3]},
      {stage3_16[3]},
      {stage4_17[3],stage4_16[7],stage4_15[7],stage4_14[11],stage4_13[20]}
   );
   gpc606_5 gpc1965 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[4],stage4_16[8],stage4_15[8],stage4_14[12],stage4_13[21]}
   );
   gpc606_5 gpc1966 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[5],stage4_16[9],stage4_15[9],stage4_14[13],stage4_13[22]}
   );
   gpc606_5 gpc1967 (
      {stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29]},
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage4_17[6],stage4_16[10],stage4_15[10],stage4_14[14],stage4_13[23]}
   );
   gpc606_5 gpc1968 (
      {stage3_13[30], stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35]},
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27]},
      {stage4_17[7],stage4_16[11],stage4_15[11],stage4_14[15],stage4_13[24]}
   );
   gpc606_5 gpc1969 (
      {stage3_13[36], stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41]},
      {stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33]},
      {stage4_17[8],stage4_16[12],stage4_15[12],stage4_14[16],stage4_13[25]}
   );
   gpc615_5 gpc1970 (
      {stage3_14[48], stage3_14[49], stage3_14[50], stage3_14[51], stage3_14[52]},
      {stage3_15[34]},
      {stage3_16[4], stage3_16[5], stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9]},
      {stage4_18[0],stage4_17[9],stage4_16[13],stage4_15[13],stage4_14[17]}
   );
   gpc615_5 gpc1971 (
      {stage3_14[53], stage3_14[54], stage3_14[55], stage3_14[56], stage3_14[57]},
      {stage3_15[35]},
      {stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage4_18[1],stage4_17[10],stage4_16[14],stage4_15[14],stage4_14[18]}
   );
   gpc606_5 gpc1972 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40], stage3_15[41]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[2],stage4_17[11],stage4_16[15],stage4_15[15]}
   );
   gpc606_5 gpc1973 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46], stage3_15[47]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[3],stage4_17[12],stage4_16[16],stage4_15[16]}
   );
   gpc615_5 gpc1974 (
      {stage3_15[48], stage3_15[49], stage3_15[50], stage3_15[51], stage3_15[52]},
      {stage3_16[16]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[4],stage4_17[13],stage4_16[17],stage4_15[17]}
   );
   gpc606_5 gpc1975 (
      {stage3_16[17], stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[5],stage4_17[14],stage4_16[18]}
   );
   gpc606_5 gpc1976 (
      {stage3_16[23], stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[6],stage4_17[15],stage4_16[19]}
   );
   gpc606_5 gpc1977 (
      {stage3_16[29], stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34]},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[5],stage4_18[7],stage4_17[16],stage4_16[20]}
   );
   gpc606_5 gpc1978 (
      {stage3_16[35], stage3_16[36], stage3_16[37], stage3_16[38], stage3_16[39], stage3_16[40]},
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23]},
      {stage4_20[3],stage4_19[6],stage4_18[8],stage4_17[17],stage4_16[21]}
   );
   gpc606_5 gpc1979 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[7],stage4_18[9],stage4_17[18]}
   );
   gpc606_5 gpc1980 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[8],stage4_18[10],stage4_17[19]}
   );
   gpc1_1 gpc1981 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1982 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1983 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1984 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1985 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1986 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1987 (
      {stage3_2[10]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1988 (
      {stage3_2[11]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1989 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1990 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1991 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1992 (
      {stage3_2[15]},
      {stage4_2[9]}
   );
   gpc1_1 gpc1993 (
      {stage3_2[16]},
      {stage4_2[10]}
   );
   gpc1_1 gpc1994 (
      {stage3_3[24]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1995 (
      {stage3_3[25]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1996 (
      {stage3_3[26]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1997 (
      {stage3_3[27]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1998 (
      {stage3_3[28]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1999 (
      {stage3_4[20]},
      {stage4_4[7]}
   );
   gpc1_1 gpc2000 (
      {stage3_4[21]},
      {stage4_4[8]}
   );
   gpc1_1 gpc2001 (
      {stage3_4[22]},
      {stage4_4[9]}
   );
   gpc1_1 gpc2002 (
      {stage3_4[23]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2003 (
      {stage3_4[24]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2004 (
      {stage3_4[25]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2005 (
      {stage3_4[26]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2006 (
      {stage3_4[27]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2007 (
      {stage3_4[28]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2008 (
      {stage3_4[29]},
      {stage4_4[16]}
   );
   gpc1_1 gpc2009 (
      {stage3_4[30]},
      {stage4_4[17]}
   );
   gpc1_1 gpc2010 (
      {stage3_4[31]},
      {stage4_4[18]}
   );
   gpc1_1 gpc2011 (
      {stage3_4[32]},
      {stage4_4[19]}
   );
   gpc1_1 gpc2012 (
      {stage3_4[33]},
      {stage4_4[20]}
   );
   gpc1_1 gpc2013 (
      {stage3_4[34]},
      {stage4_4[21]}
   );
   gpc1_1 gpc2014 (
      {stage3_4[35]},
      {stage4_4[22]}
   );
   gpc1_1 gpc2015 (
      {stage3_4[36]},
      {stage4_4[23]}
   );
   gpc1_1 gpc2016 (
      {stage3_4[37]},
      {stage4_4[24]}
   );
   gpc1_1 gpc2017 (
      {stage3_4[38]},
      {stage4_4[25]}
   );
   gpc1_1 gpc2018 (
      {stage3_4[39]},
      {stage4_4[26]}
   );
   gpc1_1 gpc2019 (
      {stage3_5[47]},
      {stage4_5[14]}
   );
   gpc1_1 gpc2020 (
      {stage3_6[31]},
      {stage4_6[15]}
   );
   gpc1_1 gpc2021 (
      {stage3_6[32]},
      {stage4_6[16]}
   );
   gpc1_1 gpc2022 (
      {stage3_6[33]},
      {stage4_6[17]}
   );
   gpc1_1 gpc2023 (
      {stage3_6[34]},
      {stage4_6[18]}
   );
   gpc1_1 gpc2024 (
      {stage3_6[35]},
      {stage4_6[19]}
   );
   gpc1_1 gpc2025 (
      {stage3_6[36]},
      {stage4_6[20]}
   );
   gpc1_1 gpc2026 (
      {stage3_6[37]},
      {stage4_6[21]}
   );
   gpc1_1 gpc2027 (
      {stage3_7[42]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2028 (
      {stage3_7[43]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2029 (
      {stage3_7[44]},
      {stage4_7[15]}
   );
   gpc1_1 gpc2030 (
      {stage3_7[45]},
      {stage4_7[16]}
   );
   gpc1_1 gpc2031 (
      {stage3_8[28]},
      {stage4_8[13]}
   );
   gpc1_1 gpc2032 (
      {stage3_8[29]},
      {stage4_8[14]}
   );
   gpc1_1 gpc2033 (
      {stage3_8[30]},
      {stage4_8[15]}
   );
   gpc1_1 gpc2034 (
      {stage3_8[31]},
      {stage4_8[16]}
   );
   gpc1_1 gpc2035 (
      {stage3_8[32]},
      {stage4_8[17]}
   );
   gpc1_1 gpc2036 (
      {stage3_8[33]},
      {stage4_8[18]}
   );
   gpc1_1 gpc2037 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc2038 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc2039 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc2040 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc2041 (
      {stage3_8[38]},
      {stage4_8[23]}
   );
   gpc1_1 gpc2042 (
      {stage3_8[39]},
      {stage4_8[24]}
   );
   gpc1_1 gpc2043 (
      {stage3_8[40]},
      {stage4_8[25]}
   );
   gpc1_1 gpc2044 (
      {stage3_9[48]},
      {stage4_9[21]}
   );
   gpc1_1 gpc2045 (
      {stage3_9[49]},
      {stage4_9[22]}
   );
   gpc1_1 gpc2046 (
      {stage3_9[50]},
      {stage4_9[23]}
   );
   gpc1_1 gpc2047 (
      {stage3_9[51]},
      {stage4_9[24]}
   );
   gpc1_1 gpc2048 (
      {stage3_10[44]},
      {stage4_10[18]}
   );
   gpc1_1 gpc2049 (
      {stage3_10[45]},
      {stage4_10[19]}
   );
   gpc1_1 gpc2050 (
      {stage3_10[46]},
      {stage4_10[20]}
   );
   gpc1_1 gpc2051 (
      {stage3_10[47]},
      {stage4_10[21]}
   );
   gpc1_1 gpc2052 (
      {stage3_10[48]},
      {stage4_10[22]}
   );
   gpc1_1 gpc2053 (
      {stage3_10[49]},
      {stage4_10[23]}
   );
   gpc1_1 gpc2054 (
      {stage3_10[50]},
      {stage4_10[24]}
   );
   gpc1_1 gpc2055 (
      {stage3_10[51]},
      {stage4_10[25]}
   );
   gpc1_1 gpc2056 (
      {stage3_10[52]},
      {stage4_10[26]}
   );
   gpc1_1 gpc2057 (
      {stage3_10[53]},
      {stage4_10[27]}
   );
   gpc1_1 gpc2058 (
      {stage3_10[54]},
      {stage4_10[28]}
   );
   gpc1_1 gpc2059 (
      {stage3_10[55]},
      {stage4_10[29]}
   );
   gpc1_1 gpc2060 (
      {stage3_10[56]},
      {stage4_10[30]}
   );
   gpc1_1 gpc2061 (
      {stage3_10[57]},
      {stage4_10[31]}
   );
   gpc1_1 gpc2062 (
      {stage3_10[58]},
      {stage4_10[32]}
   );
   gpc1_1 gpc2063 (
      {stage3_10[59]},
      {stage4_10[33]}
   );
   gpc1_1 gpc2064 (
      {stage3_10[60]},
      {stage4_10[34]}
   );
   gpc1_1 gpc2065 (
      {stage3_10[61]},
      {stage4_10[35]}
   );
   gpc1_1 gpc2066 (
      {stage3_10[62]},
      {stage4_10[36]}
   );
   gpc1_1 gpc2067 (
      {stage3_10[63]},
      {stage4_10[37]}
   );
   gpc1_1 gpc2068 (
      {stage3_11[54]},
      {stage4_11[15]}
   );
   gpc1_1 gpc2069 (
      {stage3_11[55]},
      {stage4_11[16]}
   );
   gpc1_1 gpc2070 (
      {stage3_11[56]},
      {stage4_11[17]}
   );
   gpc1_1 gpc2071 (
      {stage3_11[57]},
      {stage4_11[18]}
   );
   gpc1_1 gpc2072 (
      {stage3_11[58]},
      {stage4_11[19]}
   );
   gpc1_1 gpc2073 (
      {stage3_11[59]},
      {stage4_11[20]}
   );
   gpc1_1 gpc2074 (
      {stage3_11[60]},
      {stage4_11[21]}
   );
   gpc1_1 gpc2075 (
      {stage3_12[48]},
      {stage4_12[19]}
   );
   gpc1_1 gpc2076 (
      {stage3_12[49]},
      {stage4_12[20]}
   );
   gpc1_1 gpc2077 (
      {stage3_12[50]},
      {stage4_12[21]}
   );
   gpc1_1 gpc2078 (
      {stage3_12[51]},
      {stage4_12[22]}
   );
   gpc1_1 gpc2079 (
      {stage3_12[52]},
      {stage4_12[23]}
   );
   gpc1_1 gpc2080 (
      {stage3_15[53]},
      {stage4_15[18]}
   );
   gpc1_1 gpc2081 (
      {stage3_15[54]},
      {stage4_15[19]}
   );
   gpc1_1 gpc2082 (
      {stage3_15[55]},
      {stage4_15[20]}
   );
   gpc1_1 gpc2083 (
      {stage3_15[56]},
      {stage4_15[21]}
   );
   gpc1_1 gpc2084 (
      {stage3_16[41]},
      {stage4_16[22]}
   );
   gpc1_1 gpc2085 (
      {stage3_16[42]},
      {stage4_16[23]}
   );
   gpc1_1 gpc2086 (
      {stage3_16[43]},
      {stage4_16[24]}
   );
   gpc1_1 gpc2087 (
      {stage3_16[44]},
      {stage4_16[25]}
   );
   gpc1_1 gpc2088 (
      {stage3_16[45]},
      {stage4_16[26]}
   );
   gpc1_1 gpc2089 (
      {stage3_16[46]},
      {stage4_16[27]}
   );
   gpc1_1 gpc2090 (
      {stage3_16[47]},
      {stage4_16[28]}
   );
   gpc1_1 gpc2091 (
      {stage3_16[48]},
      {stage4_16[29]}
   );
   gpc1_1 gpc2092 (
      {stage3_16[49]},
      {stage4_16[30]}
   );
   gpc1_1 gpc2093 (
      {stage3_17[30]},
      {stage4_17[20]}
   );
   gpc1_1 gpc2094 (
      {stage3_17[31]},
      {stage4_17[21]}
   );
   gpc1_1 gpc2095 (
      {stage3_18[24]},
      {stage4_18[11]}
   );
   gpc1_1 gpc2096 (
      {stage3_18[25]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2097 (
      {stage3_19[12]},
      {stage4_19[9]}
   );
   gpc1_1 gpc2098 (
      {stage3_19[13]},
      {stage4_19[10]}
   );
   gpc1_1 gpc2099 (
      {stage3_20[0]},
      {stage4_20[6]}
   );
   gpc1_1 gpc2100 (
      {stage3_20[1]},
      {stage4_20[7]}
   );
   gpc1_1 gpc2101 (
      {stage3_20[2]},
      {stage4_20[8]}
   );
   gpc1_1 gpc2102 (
      {stage3_20[3]},
      {stage4_20[9]}
   );
   gpc1_1 gpc2103 (
      {stage3_20[4]},
      {stage4_20[10]}
   );
   gpc1_1 gpc2104 (
      {stage3_20[5]},
      {stage4_20[11]}
   );
   gpc1_1 gpc2105 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc1_1 gpc2106 (
      {stage3_21[1]},
      {stage4_21[3]}
   );
   gpc615_5 gpc2107 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc606_5 gpc2108 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1406_5 gpc2109 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc606_5 gpc2110 (
      {stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16], stage4_4[17]},
      {stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9]},
      {stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc606_5 gpc2111 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc615_5 gpc2112 (
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[3],stage5_7[4]}
   );
   gpc615_5 gpc2113 (
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[2],stage5_8[4],stage5_7[5]}
   );
   gpc1163_5 gpc2114 (
      {stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17]},
      {stage4_10[0]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[3],stage5_8[5]}
   );
   gpc1163_5 gpc2115 (
      {stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_9[18], stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23]},
      {stage4_10[1]},
      {stage4_11[1]},
      {stage5_12[1],stage5_11[3],stage5_10[3],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc2116 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12], stage4_8[13]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[2],stage5_11[4],stage5_10[4],stage5_9[5],stage5_8[7]}
   );
   gpc606_5 gpc2117 (
      {stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17], stage4_8[18], stage4_8[19]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[3],stage5_11[5],stage5_10[5],stage5_9[6],stage5_8[8]}
   );
   gpc606_5 gpc2118 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19]},
      {stage5_12[4],stage5_11[6],stage5_10[6],stage5_9[7],stage5_8[9]}
   );
   gpc606_5 gpc2119 (
      {stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24], stage4_10[25]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[5],stage5_11[7],stage5_10[7]}
   );
   gpc606_5 gpc2120 (
      {stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30], stage4_10[31]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[1],stage5_12[6],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc2121 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[12]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc2122 (
      {stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage4_12[13]},
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[8],stage5_11[10]}
   );
   gpc615_5 gpc2123 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16]},
      {stage4_12[14]},
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[9],stage5_11[11]}
   );
   gpc615_5 gpc2124 (
      {stage4_11[17], stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21]},
      {stage4_12[15]},
      {stage4_13[18], stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[10],stage5_11[12]}
   );
   gpc606_5 gpc2125 (
      {stage4_12[16], stage4_12[17], stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[11]}
   );
   gpc615_5 gpc2126 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc2127 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc2128 (
      {stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage4_16[12]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7]}
   );
   gpc615_5 gpc2129 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[13]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8]}
   );
   gpc615_5 gpc2130 (
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16]},
      {stage4_16[14]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc606_5 gpc2131 (
      {stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18], stage4_16[19], stage4_16[20]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[3],stage5_18[5],stage5_17[5],stage5_16[6]}
   );
   gpc606_5 gpc2132 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], 1'b0, 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[4],stage5_18[6],stage5_17[6]}
   );
   gpc606_5 gpc2133 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[5],stage5_18[7]}
   );
   gpc1343_5 gpc2134 (
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {1'b0},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[6]}
   );
   gpc1_1 gpc2135 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc2136 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc2137 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc2138 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc2139 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc2140 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc2141 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2142 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2143 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2144 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2145 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2146 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2147 (
      {stage4_2[9]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2148 (
      {stage4_2[10]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2149 (
      {stage4_3[7]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2150 (
      {stage4_3[8]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2151 (
      {stage4_3[9]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2152 (
      {stage4_3[10]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2153 (
      {stage4_4[18]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2154 (
      {stage4_4[19]},
      {stage5_4[5]}
   );
   gpc1_1 gpc2155 (
      {stage4_4[20]},
      {stage5_4[6]}
   );
   gpc1_1 gpc2156 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc2157 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc2158 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc2159 (
      {stage4_4[24]},
      {stage5_4[10]}
   );
   gpc1_1 gpc2160 (
      {stage4_4[25]},
      {stage5_4[11]}
   );
   gpc1_1 gpc2161 (
      {stage4_4[26]},
      {stage5_4[12]}
   );
   gpc1_1 gpc2162 (
      {stage4_5[12]},
      {stage5_5[5]}
   );
   gpc1_1 gpc2163 (
      {stage4_5[13]},
      {stage5_5[6]}
   );
   gpc1_1 gpc2164 (
      {stage4_5[14]},
      {stage5_5[7]}
   );
   gpc1_1 gpc2165 (
      {stage4_6[10]},
      {stage5_6[5]}
   );
   gpc1_1 gpc2166 (
      {stage4_6[11]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2167 (
      {stage4_6[12]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2168 (
      {stage4_6[13]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2169 (
      {stage4_6[14]},
      {stage5_6[9]}
   );
   gpc1_1 gpc2170 (
      {stage4_6[15]},
      {stage5_6[10]}
   );
   gpc1_1 gpc2171 (
      {stage4_6[16]},
      {stage5_6[11]}
   );
   gpc1_1 gpc2172 (
      {stage4_6[17]},
      {stage5_6[12]}
   );
   gpc1_1 gpc2173 (
      {stage4_6[18]},
      {stage5_6[13]}
   );
   gpc1_1 gpc2174 (
      {stage4_6[19]},
      {stage5_6[14]}
   );
   gpc1_1 gpc2175 (
      {stage4_6[20]},
      {stage5_6[15]}
   );
   gpc1_1 gpc2176 (
      {stage4_6[21]},
      {stage5_6[16]}
   );
   gpc1_1 gpc2177 (
      {stage4_9[24]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2178 (
      {stage4_10[32]},
      {stage5_10[9]}
   );
   gpc1_1 gpc2179 (
      {stage4_10[33]},
      {stage5_10[10]}
   );
   gpc1_1 gpc2180 (
      {stage4_10[34]},
      {stage5_10[11]}
   );
   gpc1_1 gpc2181 (
      {stage4_10[35]},
      {stage5_10[12]}
   );
   gpc1_1 gpc2182 (
      {stage4_10[36]},
      {stage5_10[13]}
   );
   gpc1_1 gpc2183 (
      {stage4_10[37]},
      {stage5_10[14]}
   );
   gpc1_1 gpc2184 (
      {stage4_12[22]},
      {stage5_12[12]}
   );
   gpc1_1 gpc2185 (
      {stage4_12[23]},
      {stage5_12[13]}
   );
   gpc1_1 gpc2186 (
      {stage4_13[24]},
      {stage5_13[7]}
   );
   gpc1_1 gpc2187 (
      {stage4_13[25]},
      {stage5_13[8]}
   );
   gpc1_1 gpc2188 (
      {stage4_14[16]},
      {stage5_14[9]}
   );
   gpc1_1 gpc2189 (
      {stage4_14[17]},
      {stage5_14[10]}
   );
   gpc1_1 gpc2190 (
      {stage4_14[18]},
      {stage5_14[11]}
   );
   gpc1_1 gpc2191 (
      {stage4_15[17]},
      {stage5_15[10]}
   );
   gpc1_1 gpc2192 (
      {stage4_15[18]},
      {stage5_15[11]}
   );
   gpc1_1 gpc2193 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc2194 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc2195 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc2196 (
      {stage4_16[21]},
      {stage5_16[7]}
   );
   gpc1_1 gpc2197 (
      {stage4_16[22]},
      {stage5_16[8]}
   );
   gpc1_1 gpc2198 (
      {stage4_16[23]},
      {stage5_16[9]}
   );
   gpc1_1 gpc2199 (
      {stage4_16[24]},
      {stage5_16[10]}
   );
   gpc1_1 gpc2200 (
      {stage4_16[25]},
      {stage5_16[11]}
   );
   gpc1_1 gpc2201 (
      {stage4_16[26]},
      {stage5_16[12]}
   );
   gpc1_1 gpc2202 (
      {stage4_16[27]},
      {stage5_16[13]}
   );
   gpc1_1 gpc2203 (
      {stage4_16[28]},
      {stage5_16[14]}
   );
   gpc1_1 gpc2204 (
      {stage4_16[29]},
      {stage5_16[15]}
   );
   gpc1_1 gpc2205 (
      {stage4_16[30]},
      {stage5_16[16]}
   );
   gpc1_1 gpc2206 (
      {stage4_18[12]},
      {stage5_18[8]}
   );
   gpc1_1 gpc2207 (
      {stage4_19[9]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2208 (
      {stage4_19[10]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2209 (
      {stage4_20[10]},
      {stage5_20[4]}
   );
   gpc1_1 gpc2210 (
      {stage4_20[11]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2211 (
      {stage4_21[3]},
      {stage5_21[3]}
   );
   gpc1163_5 gpc2212 (
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[0]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc207_4 gpc2213 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[0],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc7_3 gpc2214 (
      {stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5], stage5_5[6], stage5_5[7]},
      {stage6_7[1],stage6_6[2],stage6_5[2]}
   );
   gpc1325_5 gpc2215 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[3]}
   );
   gpc1325_5 gpc2216 (
      {stage5_6[7], stage5_6[8], stage5_6[9], stage5_6[10], stage5_6[11]},
      {stage5_7[2], stage5_7[3]},
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[4]}
   );
   gpc1325_5 gpc2217 (
      {stage5_6[12], stage5_6[13], stage5_6[14], stage5_6[15], stage5_6[16]},
      {stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7], stage5_8[8]},
      {stage5_9[2]},
      {stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[5]}
   );
   gpc1163_5 gpc2218 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[3]}
   );
   gpc1163_5 gpc2219 (
      {stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage5_11[6], stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11]},
      {stage5_12[1]},
      {stage5_13[1]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[1],stage6_10[4]}
   );
   gpc615_5 gpc2220 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10]},
      {stage5_11[12]},
      {stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7]},
      {stage6_14[2],stage6_13[2],stage6_12[2],stage6_11[2],stage6_10[5]}
   );
   gpc2116_5 gpc2221 (
      {stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {stage5_13[2]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[3]}
   );
   gpc623_5 gpc2222 (
      {stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[1], stage5_14[2]},
      {stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc1423_5 gpc2223 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5]}
   );
   gpc615_5 gpc2224 (
      {stage5_14[6], stage5_14[7], stage5_14[8], stage5_14[9], stage5_14[10]},
      {stage5_15[10]},
      {stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], stage5_16[8], stage5_16[9]},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[3],stage6_14[6]}
   );
   gpc606_5 gpc2225 (
      {stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14], stage5_16[15]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[3],stage6_16[4]}
   );
   gpc606_5 gpc2226 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[1],stage6_19[1],stage6_18[3],stage6_17[4]}
   );
   gpc1_1 gpc2227 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc2228 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2229 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2230 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2231 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2232 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2233 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc2234 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2235 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc2236 (
      {stage5_2[4]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2237 (
      {stage5_2[5]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2238 (
      {stage5_2[6]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2239 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2240 (
      {stage5_4[9]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2241 (
      {stage5_4[10]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2242 (
      {stage5_4[11]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2243 (
      {stage5_4[12]},
      {stage6_4[6]}
   );
   gpc1_1 gpc2244 (
      {stage5_8[9]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2245 (
      {stage5_9[3]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2246 (
      {stage5_9[4]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2247 (
      {stage5_9[5]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2248 (
      {stage5_9[6]},
      {stage6_9[6]}
   );
   gpc1_1 gpc2249 (
      {stage5_9[7]},
      {stage6_9[7]}
   );
   gpc1_1 gpc2250 (
      {stage5_9[8]},
      {stage6_9[8]}
   );
   gpc1_1 gpc2251 (
      {stage5_10[11]},
      {stage6_10[6]}
   );
   gpc1_1 gpc2252 (
      {stage5_10[12]},
      {stage6_10[7]}
   );
   gpc1_1 gpc2253 (
      {stage5_10[13]},
      {stage6_10[8]}
   );
   gpc1_1 gpc2254 (
      {stage5_10[14]},
      {stage6_10[9]}
   );
   gpc1_1 gpc2255 (
      {stage5_13[6]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2256 (
      {stage5_13[7]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2257 (
      {stage5_13[8]},
      {stage6_13[7]}
   );
   gpc1_1 gpc2258 (
      {stage5_14[11]},
      {stage6_14[7]}
   );
   gpc1_1 gpc2259 (
      {stage5_15[11]},
      {stage6_15[4]}
   );
   gpc1_1 gpc2260 (
      {stage5_15[12]},
      {stage6_15[5]}
   );
   gpc1_1 gpc2261 (
      {stage5_15[13]},
      {stage6_15[6]}
   );
   gpc1_1 gpc2262 (
      {stage5_15[14]},
      {stage6_15[7]}
   );
   gpc1_1 gpc2263 (
      {stage5_16[16]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2264 (
      {stage5_18[6]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2265 (
      {stage5_18[7]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2266 (
      {stage5_18[8]},
      {stage6_18[6]}
   );
   gpc1_1 gpc2267 (
      {stage5_19[6]},
      {stage6_19[2]}
   );
   gpc1_1 gpc2268 (
      {stage5_19[7]},
      {stage6_19[3]}
   );
   gpc1_1 gpc2269 (
      {stage5_19[8]},
      {stage6_19[4]}
   );
   gpc1_1 gpc2270 (
      {stage5_20[0]},
      {stage6_20[2]}
   );
   gpc1_1 gpc2271 (
      {stage5_20[1]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2272 (
      {stage5_20[2]},
      {stage6_20[4]}
   );
   gpc1_1 gpc2273 (
      {stage5_20[3]},
      {stage6_20[5]}
   );
   gpc1_1 gpc2274 (
      {stage5_20[4]},
      {stage6_20[6]}
   );
   gpc1_1 gpc2275 (
      {stage5_20[5]},
      {stage6_20[7]}
   );
   gpc1_1 gpc2276 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc2277 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc2278 (
      {stage5_21[2]},
      {stage6_21[3]}
   );
   gpc1_1 gpc2279 (
      {stage5_21[3]},
      {stage6_21[4]}
   );
   gpc1_1 gpc2280 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
   gpc1_1 gpc2281 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc2282 (
      {stage5_23[0]},
      {stage6_23[0]}
   );
   gpc1406_5 gpc2283 (
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[0]}
   );
   gpc117_4 gpc2284 (
      {stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5], stage6_9[6], stage6_9[7]},
      {stage6_10[0]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc1415_5 gpc2285 (
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[2]}
   );
   gpc606_5 gpc2286 (
      {stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc606_5 gpc2287 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[1],stage7_16[1],stage7_15[1],stage7_14[2]}
   );
   gpc606_5 gpc2288 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc1406_5 gpc2289 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc1_1 gpc2290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc2291 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2292 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc2293 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc2294 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc2295 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc2296 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc2297 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2298 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc2299 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc2300 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc2301 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc2302 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc2303 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc2304 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc2305 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc2306 (
      {stage6_4[2]},
      {stage7_4[2]}
   );
   gpc1_1 gpc2307 (
      {stage6_4[3]},
      {stage7_4[3]}
   );
   gpc1_1 gpc2308 (
      {stage6_4[4]},
      {stage7_4[4]}
   );
   gpc1_1 gpc2309 (
      {stage6_4[5]},
      {stage7_4[5]}
   );
   gpc1_1 gpc2310 (
      {stage6_4[6]},
      {stage7_4[6]}
   );
   gpc1_1 gpc2311 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc2312 (
      {stage6_5[1]},
      {stage7_5[1]}
   );
   gpc1_1 gpc2313 (
      {stage6_5[2]},
      {stage7_5[2]}
   );
   gpc1_1 gpc2314 (
      {stage6_7[0]},
      {stage7_7[1]}
   );
   gpc1_1 gpc2315 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc2316 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc2317 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc2318 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc2319 (
      {stage6_9[8]},
      {stage7_9[2]}
   );
   gpc1_1 gpc2320 (
      {stage6_10[6]},
      {stage7_10[3]}
   );
   gpc1_1 gpc2321 (
      {stage6_10[7]},
      {stage7_10[4]}
   );
   gpc1_1 gpc2322 (
      {stage6_10[8]},
      {stage7_10[5]}
   );
   gpc1_1 gpc2323 (
      {stage6_10[9]},
      {stage7_10[6]}
   );
   gpc1_1 gpc2324 (
      {stage6_11[2]},
      {stage7_11[2]}
   );
   gpc1_1 gpc2325 (
      {stage6_13[7]},
      {stage7_13[2]}
   );
   gpc1_1 gpc2326 (
      {stage6_14[6]},
      {stage7_14[3]}
   );
   gpc1_1 gpc2327 (
      {stage6_14[7]},
      {stage7_14[4]}
   );
   gpc1_1 gpc2328 (
      {stage6_15[6]},
      {stage7_15[2]}
   );
   gpc1_1 gpc2329 (
      {stage6_15[7]},
      {stage7_15[3]}
   );
   gpc1_1 gpc2330 (
      {stage6_17[0]},
      {stage7_17[2]}
   );
   gpc1_1 gpc2331 (
      {stage6_17[1]},
      {stage7_17[3]}
   );
   gpc1_1 gpc2332 (
      {stage6_17[2]},
      {stage7_17[4]}
   );
   gpc1_1 gpc2333 (
      {stage6_17[3]},
      {stage7_17[5]}
   );
   gpc1_1 gpc2334 (
      {stage6_17[4]},
      {stage7_17[6]}
   );
   gpc1_1 gpc2335 (
      {stage6_18[6]},
      {stage7_18[2]}
   );
   gpc1_1 gpc2336 (
      {stage6_20[6]},
      {stage7_20[2]}
   );
   gpc1_1 gpc2337 (
      {stage6_20[7]},
      {stage7_20[3]}
   );
   gpc1_1 gpc2338 (
      {stage6_21[4]},
      {stage7_21[2]}
   );
   gpc1_1 gpc2339 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc2340 (
      {stage6_23[0]},
      {stage7_23[1]}
   );
   gpc615_5 gpc2341 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc7_3 gpc2342 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc615_5 gpc2343 (
      {stage7_5[0], stage7_5[1], stage7_5[2], 1'b0, 1'b0},
      {stage7_6[0]},
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5]},
      {stage8_9[0],stage8_8[0],stage8_7[0],stage8_6[1],stage8_5[1]}
   );
   gpc23_3 gpc2344 (
      {stage7_9[0], stage7_9[1], stage7_9[2]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc135_4 gpc2345 (
      {stage7_10[2], stage7_10[3], stage7_10[4], stage7_10[5], stage7_10[6]},
      {stage7_11[0], stage7_11[1], stage7_11[2]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1]}
   );
   gpc1343_5 gpc2346 (
      {stage7_13[0], stage7_13[1], stage7_13[2]},
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3]},
      {stage7_15[0], stage7_15[1], stage7_15[2]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc7_3 gpc2347 (
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3], stage7_17[4], stage7_17[5], stage7_17[6]},
      {stage8_19[0],stage8_18[0],stage8_17[1]}
   );
   gpc1325_5 gpc2348 (
      {stage7_18[0], stage7_18[1], stage7_18[2], 1'b0, 1'b0},
      {stage7_19[0], stage7_19[1]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1],stage8_18[1]}
   );
   gpc1163_5 gpc2349 (
      {stage7_21[1], stage7_21[2], 1'b0},
      {stage7_22[0], stage7_22[1], stage7_22[2], 1'b0, 1'b0, 1'b0},
      {stage7_23[0]},
      {1'b0},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1]}
   );
   gpc1_1 gpc2350 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc2351 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc2352 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc2353 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc2354 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc2355 (
      {stage7_14[4]},
      {stage8_14[1]}
   );
   gpc1_1 gpc2356 (
      {stage7_15[3]},
      {stage8_15[1]}
   );
   gpc1_1 gpc2357 (
      {stage7_16[1]},
      {stage8_16[1]}
   );
   gpc1_1 gpc2358 (
      {stage7_20[3]},
      {stage8_20[1]}
   );
   gpc1_1 gpc2359 (
      {stage7_23[1]},
      {stage8_23[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor_CLA512_16 compressor_CLA512_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h24afeee679ed09d4e220026a03c1f8ef93d4ff8f88147a9ddded753d80bb95c7435d5babacd5c3fefda90c81e1622afd9786c7770f555ed98e616058c403ac66703e8a619be8e4e2a0b61e263d2a115f293b1ae1bed4de523a7124bc8a0aa7207b1ef3da41c0c81fcb3f3cd4dab67ccc4038ab81845e2748517a4760e7cbbc84ed2e38bca2a8cf1670a81a572a7bb38e7b9548deb6c3d1e4c309c3b2910a885b1c665c68a50a49be1fa140867a875cf99d248ef0692c8464ff4f948f283ce45eb7d897cf3eb067175cd190f71dcc536314202f052da35831cff6b88364518d7feda3c2ef383b936cc5656981e8055d9128cf849ec429b96d10039c1f09c6a9d52d362c792f5a5a6bae8c83883099cf9da80d43fc4e1c3e96a6b3e5d0b33cc632fdcffb9b61b9d5ceefcbd2e60034e1a176e9f04cca7e7feea4e2ec5682378df0a69e728a5f6bb6a3fc156b5505546e616c3303210784596dbaea2290b181090701612192f97cae764a3d38b4f32864511e6b1f3a6567aa65897b048afec7791667a419f3f00d694e57a0e9aaf5c280e903629cffbe749fd68ae4a3605eff813db219d0d55277c3f16ab875802708ea10e656cbb94e527d11774566114d9c884b3188d058e55202722a25140bd40572daba165cb2cda8bc933d3210e3d3962dfe893a62e2c16fb43adcd4333611f5716f29281a9812f76d80aeb35e608abb7c79651f46d3696d523ec8a0230a9d229ace80b1d0fe1442831a918248f6740cf472c8188e138e94e2f736a3f3efa7d2154b5f542f185656a3cddae9a0a5e452b6fcb0ae9f2f1d0fa3f8b6f845f8033fd01690adbbc37387f08dbc52bdb9061b16d123ad686d8a42969484df0a8067c7bf1496b5810793fcba43b3f50de4534bf0dbc120fb78daa615db1f25f96f7e8aaf5912fe51363c1b581d28c9954d2980a7affb3dbcb185c516a7fab09e8a993389ab03217d736f5169394b6fe602baf0c9dc4756756f0fcca6707bd9a6a976b02777c1482245703828004968f8d99f0f4be4285c1841be0d8a372f57818a08e3e6ca367e9b6920d071c3a33909ed7ee0c452acf7b4d1ff83366d30f600d05f190e00a4dd95566f15ca4df7836d19aa043d80cd1b10c5d59b8a06bc5e84fa10499c9e2fb5fb8ef46db76e092d868c4a31a3b1378507f858d0a8f94c0d6d1a317f3ec5a6f3a427863d5f5ef7f3899018aca30e9e447eccbcacbf5ce4e7b3de12841e5af7d9813a022868f7eb0883a9df1bb80ae1a3b5c4e6d723a5f9d184cf11349211abcd53c2ea16fa6ea67989553c4ea3cca4476f2c89f0bacaa3476817379e2894316e9711321a31289f2a620688350a75e0e6c76882be1e9a5cbf75258f957c877b2add0b28e4bb9827b9ed0c6294a584d929f1b3c254e9b808a9d95a9d43e92c288871e3c9b0b9bb204473c0dc93f3d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc0aa69acaebddd8136d22300325b29a56cad52ee627cf574026e552a290f55584a3372d93e7f413ac11b3324f830b4179a77f3a9b1f950e335a403f1f9ea4178bc81e91456ff279222986f44f08c548d72815ae67bbae6280616133a0d1cd6c439dc6435d9ec5e915142d2d7225654105a4bbf387033a1a7624c8474d9e0a93d8b533bec42dfa48db7487348a2390f0473b149b753b95c89b78d326247e8e929e83b810ff1e1d7cfb3a361d95d23be32a1e76716b8d9046a778554765ca00bad861d72f87e1020cf5061810eb1c047b27d4801165bb167b832ba00d49f73ac1e03aacd3915705e9396a0d2e62aad4d60f45473053df2da83804a4353bf685075631abae25be8feb21300723fdff4d8500191df21fbc6ccadb2d82cdc159d7a9133c0d32a99c304c3ff241c992055431a2a2edbc7eb2e1573f6131e1ddf8d1351a391f80ea3061a3d78aff21199bf0f54784359a648a17dfe1f2aed5221515f2e249ee45bf72f4d0f94021ad00022c7eb70b959c03f8b39cb0451ab9c2137cdf819c22047768c6eae33ac90797b0da6090feaea4afc7c81777ff80cb2acfd7f2329ab2a8d06558b5ef09693f01480aeddc1de02ecdc3e15ad27f6174322f9bfbe5af7138bc9e5d811808fa76b4d071b96e598f3d0dec4193c9bcbfcb289d86ac39ffa09353abf074638e0ffe4ce3b0b3079aaf2247560468bdc95b8565b47b1b1f5af0447d4b52ae33c08f7d9c0d7c320696cf93950bfc73b8c89db983f0eb265d4116974cebf176e9bde13dffccd8dfbadfbe3c60b76d43c85bda722783c9dc7196631c24dd2b02b61c9591f35bf100ed98ec74f88c9c42b22f6761c45074c3cb250a7d2d7f64fb7c9f7e9f124aae8842613748670bf3426d3faea14dfdf6c815756d4c127f4d944eb31b25625153e477932619281932164234ec81cea4fe86e842fcced3881ddd500eceea31e30acb47e70a160487fe861da03814cc96db0bfb65f833101d828eed3a70ea5c83334a3f865db25dc680fb038a68e93830f1b88b85d0f586d2298178283523a447ce66cb61b44c73ec6017f1e04d19b8348761a2a25f7fc44b5763a26c6889c1a938f474dfe1cd0b4b9443b8ca1f08d6e306f09f5973537b1d02ed78dbd9e963fb10a89668b4afa8a3a5e5e0686f786af2b5cf10782a93ce2943f1eb45a73bb907728b7898db0a8b226fb5ae8a0810598813a5e873401fff08fdb6fa88e22f343a5a3f2eee47c3db16f7507d2112f3f912085d7f8962d54b8dce4d8bd26a2f9110ebd1c4ce8d15f6831b890527e8e630d5bd68e2531f4d6f2071f2e468cf9dc042131def9e6f7e8993b4410e434201face99105c2e76086c3812047970c6a96e0ad4bb627b01b4371e134d4795594ccacd95e1451c93cc9147a49acab0ec42340410a95644cd5a1c9a4612216af830daea55ab9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he329f45b9b6c35bf706d53ab282a13de9f2d48913c976e935423e98f5c8ebb0c0dd96248bc2a4643488311f57b63297c3b4b89402d4703f6ae2f89253d1c00d49270556bfbf0de93ed1692bb19e841b47785c01a403c6a391b385d259af383783853c1598f768905d757d36e1ee19269ab69bbc3b1130da6ed5e0cf6b00ae8810cfc305d18362506172bccbe30b88c2990c0f21839ba004443bdb7411de3b3177eebac0c0e192d50055026e7740fead3027da6765e3d774b4157cee0ab137e70f16ea6fab8a2c2cd4d2fceab9e450c78dc67524780155fa849630987ae60f77079405ad62802de7acdce3b37917609f6788c2118949d0cc89dc1324831a184758b69d3896dc6a37522888fab361467b9fa3889256afe0c785e99783460d045bbcac3c78f4362a1573473efc0cbd814f7bc14d4241dacded33710c2000b19247097b1a271bc910739f3cf68931895b5450dc01ad0352ad93e0842bd2305cdaabc4f9c39a750f812a1434fd49ddc2423efa01d3c2d6a868f440e66ec70de3e61e9c482cc8ec6bbb61bf17da2de4d69890209561b6da04de6836402e43ca5428be7f865bcddc96be665843a5b57ca942d9bb822a15a8f646320c29d86ca4e44886981a2980d394c4742a73c93732ce4762b912837489b9f42de11addb5a01aa504a8e4b86fc5f4440737e7ee513a6c451351a29738d370bb2c9e456893e6b39bc11854bdb3daae1d14a5cfe4dfe290afc3146fd3b4e58a77f2fb140c46dcc377b043d9205f61b228c84a408739406b3d8d3d683c878af7875d9d3f1a82fe6146d8ac3b09965ef91815440a2cfe9b9350b11d517c3b8259528fc8efdf40912b2b8ecf7c876d51d3536c4cccf8b6d0d5f42abb6f3f1b17c04256aa0a531dd123777883944d390b54592190ff9005bf4db20b32779aab2268105fc28ea6a9e52deeaaff20106c630a1ff8bb6168913080a51d2e6c546e1f0928f6998ad991ff6d70d0e0b8c2f4809dc8602a5adbf244244427e344957ab5f7f2dd8fc72639788a5e31f831c2687269f8865793cb36383f4a1671690493eb248597a2b612f12cf3417543619190112919f7d4a32cc0291fb6b16f2df5e8ccdc55cd697e1e8f252d4991cde3635e9ae5dd79633c425a29b9bab88e04a038bbbc9f3b676ba2c747895e0db3daf31b2cab8e9f70f428c4c83216e56940d3c73353713f5b88a169216a27e28143fcba904461ecbb0252591a6c9f461ad9b26715f2868baacddb884bf3ad1f4609d8339f003c6531a95e81faa510a9d71f7f88fa3a629908a0b2104fce5bd575670e78ed6d08dd1ad0dcfb7eb904ddcb87dba76df501d1bf6740d9ce129b6258432244511c5170069ada716d5be3db13dc454678d82d467b62b6a9b26ac2a37e6f9fe6c56f6d29c75aa44d663b97b2981745a58f203ed685160e6f81f9e14de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h826fe49b8ad322fbdc75c577a06287fb85a9d573427e4b7c8e5179a018473897e020d5f868d9a584c98af58be71e288ac582ebebf26fd1b486fbc4817bdb86ed299383005ae5f7de7970114cfdad827b8ffe85a2b18f0f07d5f795c1f8cc51d49b990e1341ea4bdb2e5604c9b06a0fb4523901bc12a774b238b1965c0cc51506077653b209f03c041e227d5576bae0f970daa87ef76bdc0280add7ba26c044e87520b3e02ad99b0a12b28f1032625e0b4c6846448fb452fea617e409f4ded2417a31dcd7bd24e8ef68ea6884404c4bfcacff0ea24e7a6e15094919f288374471cbe15c495506ed3abcbe483d97d65bee6f4b22de08ddbfd8923ec222811b5f0fbb3ec585ee3728df759b3c4288fdc07e5d8cf653fe319039ad45922e53d885e22f5ccc8d691e2503a45ebc697fd5b0a395d926f3136c0dff5104887741351debfd90caecf5c068d4711127c03d0811a7ad39fada1901ee546cbc98f5d06358d806d660c12793e2c165b1920a2242f41a599c7901be60b12d4471f67d009b7f62b2f820074f98815cd3b72af4a4f09999bbe6f956b41bee3f6de23395dcb70caecf858944bac024c72d0bb769c1ca6e2f8c1a63cc85bfdc0e088a3266a61f4af281b169e86cec8f9fbd48ea7fc5c46227f81ee8e1a81f652e41d8f7011e6e5a301f26468a247396329cf3308d5f993e3e7eaacd89ae18fc65c415cd2d24f7cd53ee1e4931098fd33d510c726b32ea770266fef2bc751d00f4e537076d6a3f2adeef88a5cb60104e2ddf34883ebb600b15689cdadca98c1b68e9bb90179b781d4bd5cc9d9e4b006b3a91ab29398ba96d232e99b88940736696948fafbfcad9e68aa23029929aab64e032bcba385e2e3e877e91aaf002cf07ad62013a709f0a73aa9a0ee8e5e384d4629f555c8c49dedf59490344efab170671016f4829d62cfb2b3655ba88e0296ad664f02c1300b081270df03fa357facc716d3098c8b39200a2e313428224c92ed3d675226fcd716bd7fe2540425568befdcc72cdc4af83030de46c3cb08c189e133d0e6f9c1d83c0791397b4791a380654f00216833d31b7b548378565e2aa949efc8a408faabbd76fda97cb116a35e9bd3d912cc13cfa5c6a555f0a92749580a7e78c700928be448483987540bc693c44eef4c56c4b8f53ec34fa82d6344bae23301543d63aed816e5c7db6955ff870572f06e79172c53c201a41de1762d92f267d3fb92902a1cb3c7ea163e1b515b670041bdb627720e857f87e6bef7b3e558288f4fd1ce77e14aad73b02beaede3d68e100f2d14396717d4cff388274753d20349b7aa189fc849a902118625fcff00a6b4555e29b48bf08ae444fb17125317d70118a15daec009af436acbf9da1eed7037cac71975fd7ba434a0e962f0139cc5994f0ba718614de6bf2cd4a99cfad6b395d0c306d948f38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h387deeeba6e77d00bed764f1d18ff412cad02c485c45958bf2c0cc68cc9c0fd4cbed85e71f4a2194a20a7f036b8a67d74d295cf36b670db89e6f5c5b15b40301741f493191c48999c0200470f4c11020968ef439bd1dae29ae215ec353f1afdc827bf8564b7200ed7b4e1562f69c25961848f20f373822d2ff6441c6b404ac8b587da16a119a7142b20a34f54f7b8433eed27e8d3da4349c45c639eecdd130b900fba93f3891540d6fc18596d9393cf3c25374a7ec76dcdbc5b4128039e76d8430fa152273014b9d47b6768de951f5d448da2f9b126ce89ff98cec5b9259d1feeb5cce8c2b0052685a2c122697bdbb55aa634c1b7ea7e469ebca6f407bcf4d8a933af5567bc93159f8117a1539c2b737e0fca49dac72b66e6247af66ac6f184495febe93ca6a15638a6eb8c38cd227d172cf50f7c49ed0a2ed6826a0902ef533aeb98c88544666340682bade1b43e654c7fe68d32fd78c1126126197637d9f3719d029d32bed7b28e11e33d3158b95dd10e0c3958798c3d26dcec422896e23be13f3cac252f0052b3a078b5794fb56b5f2afc6429784046173833f3ce5025987b9ea4a32e5832f662ade1cf4adffaea1744dec2890727613eb9d3dd5b898c128caa54bf0ef926799ab01dd33e0f75fe77e2eeb176e25b06bb269158ca0a4f5c131f88f91321bf57238c7aaa4e53e6fca068b4744fe1bbab448d2af25a948ac601d162661a768e655aec476affd8aed8a578f2b2bd721e3c8e3fedd91358b0bd2a8595f6fe680727df7a435de63e3924f9fbe002189a7c85ca9ffcb4901210ce852049432950c4e30ab88344530537ea7b02387e0b6e4d5ea44641c02e3580de5a8a3e1c0274acb67c732f6e727853f57a2d3224a7146d9475edc7996316ca81576283f3bdf8cf90f3ad155fc4cf5381e27b3b7e11e2ab0f448ae6e90724127143f4e899c68c0667260b1d0ce5a77adbc36b1c9e2c57920b24c6127d1d3514468503ab3b59177aa738e48c7a30617af230a2dbe1651f1f5c1073e6761e467679ac689907a7fdb33454ff61826d88f872d7a1fc3d25179fa9f6bb838e7f5f3c6be7097aa83ca247ac104a3e0252eca9a60d177e3f63f5ef4ecbcd8f10f4d32d8f32e049dc2bca8fbb953731abb64f4846d1c9a22a88c220cddb868ecbfb0ce651bd6b9be2104c64b66697b5a04288faa99a389a3095cb217c1d20b5c4cf986bdfe841facbe10c2a7b93d8dce29f9c22a65e9a676875b5976042711e9150c302ede700855cb2969c873392a98964c087506e6236413a0ca7ac5747c18acbbb7534363c891be87e0784281c59b38ee68435259cb3e4f1ec73625a34ed0ceabf3e352fd2d3afb419d8b4bc296a2514d437457d46bbbafe635230bb0b4c0afe8bc569a0983b81a756dec85b4f35614f60cf21bcffc6397b7525f44876a5ebf03d722f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3fcf01d8658aa7326635f32d4c30ca34476b4ac63a8eb5189525159a97e79a1329f845cb7b49ca132b4ba93385e4797c4d3950750e9fce475d7f1a6ec4c1293ad619edfed3baee41d8d6dda5104e233f06892fa3fbd71c4160ca2c4fb6adab453695a008d517b9dc153d72c3a15f5d3d2ccc7bc5d54806850788c28d16a3beaa26073848a36fee05b8a85504692a9ac113430d7575763ab46d03a917834a3646c5931ecd1134a211dcc0baebb4187fcd9ad4e859f4d9df6e6479c17ba7ac73bcc34c646eab8284b73ce7fb2cc603281e9a07d55678b343023904cfb0a362e94039fe509d6d0cd810ffc7584bb1e73baf6bc5f4688d10c6048adc11bfc68e45ec7fe2f91eb9ce018bbe7fd76bbbf08006e742613e27b7381275e34bf50bb16eb77e9335da34d33d7601c05a6a673f4eecc6f8caf2b7ca66e3b4160b64d899a2ee05c148d895b9903ca4fa4702d59077bbfe1b1535f4431f62dcea20bbe96b3cc38c7f5c56552b170fbcc20b4e846cfc76ab47ce408007e8496c689e12a74cf79b3bd0fb5850e643cca017f55d8922d1e4c604ee057f131f14411ce3d6b3033e2126eda59da3609c2e905250f18adf8a5727d0d9fe79cd2be1fa8cae621a9a5e6d010359ec09570ad251fa5fe8f201b31a169723315d9765efa1303673d13b7fc88938dc5732f30d5d28d94f02850dd6c7bebc7d3f845b14a8c72dc809559dbfac2f07573315123685ac8033cc8b52b4776467cd36c2071ad91ea10ded2926000c7626fc0fa373b2489f7cd9f3e82cf2b0ab92d3150c8f84e21120b8eb82d6bd02eca610b31d393e930c9abd7724f9de3c8a712cc33814620ae52d8e5845e0e7bd1ba0a978faf31d0846b4f751825cce2fd9c481988eedc39914431f80c2e15398f040d9c257c18d067f17be5242a5fb2d6603b4157f90902763ef2e0a8cef2727e4ee57625aa554acb9d8f4e685b2a56a4983af25d6665ca97aa0ccb5e4c82a16e2d8e008db530de35dcab9ebe3db667ecb1e2f2b35a63b66dd9201eb6bf0d32214685d5c29b4b8374d91a6124830a5b6fa562fe0051d00d7cfee39946cd62d19cd2fc2650cf4a11e553b2c8582babdeb5045680ef10dd8dd12de9627f795359024fcc31a85b0e448ebb0ce3b11f7bbaf34af82fa2a343acc73b1cc5eedc57bdb416629ee653230dd4ba3d46325fe2726d7cca331bab8ad04d4c54d7b788df3f05a0421c2e40fc7de6555b036b4271b0baaf5ead0db6856f324c27de043a9da8916f1f17a137fd89f450d503a6dbf0f079387355547fb9993a9bf40ee4790060c1d7551b90ddcba64ac07eeab0f267f35a401535658a4c3d3b19dee9231bacdb5cf79c8feb4b0cf8c679919fd17fb3ef8c9595084f1810f6b685a3ce3342c2ad9ee300d98aef4673dddf476a5357765c7e24fd919b290ecc46877a5017994136b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hef51a10ba85a85bd503fef82f27401680bad72fdacd525d251d28f6f61dfccdd77ca7f37970f34272f88e916a28d51476dd10fd4a4ca696d71eb76846a69bc7aaf555ad9208c81371607daa3c37d9cd76a369c89f47bb3f1b68de49262dc30dac1423b7b3bc28992150a65ba511639647ae008ff55f9c5da75b72dbec7e5a67d415cd5b0db284e93ee4bc49928b7a4b9a425c80907ac23e8e5cb4f3e2fcfba37149b08de1fdac832f56f9488590337c8ba0a608722675b0af93f6e3119e14efb2d5f1fa248c9794a13cb5dfe8db433f50877934118cb95b49cf66e9606f7ab4f96b3c466b9fd762a366b261bf315d622493d81f4574680aef8794f670ad71c3d9764a80d542a7b2fd31fd8b67463e5be7d5b1521b7a107d15118700af02ba4fd6a5cc07b45645bca93f854ba2940f1e5f087ca66b0161c27d8c4cdf74f038b0f7fec96955e54c187d67a98ca59b9dc338d28df2ea895419653235a99a99bf65e0a14597edae51ac18367746d057bffb6f9f044bed0cb6ee0e397cc1deee3a2bf0d53628627a4208dd6d1c1a1841e38d0efe36f43d5bb7ef04e4c00ba6347fe65ac8eb652b12e1313b6f518211f74b28fc8edc0e6166d491ed69abd129d0b03a74d1fa0ec65736d80c32dcda6fb347039814abcf969eda6c10f46324bd1d3852496c51e410b0f2962b6b3d6905de89afd77b90ca03cb9d9c4b56a4133f4825363623eefc117e4997272d9bbb4c4c1891fa058a7e56fc5124bc606aeaebc19782b61f9cb3134cbc285fe956f29433a2a295472a0f77e5fe1de26f8a6ef0feb3548c80d02e9917e3d4e2e604703e15f35187b519ee507034f94bd351e63ee5574998ebff75ea3be10cccf056fb162bc69ba431577833ff0e3f4b37467cfe1ff140ea194912a840de9b2bd6495bef39995024357c92b5fbd92be1627db93dfa91b433432ea51f39284b5e8b838ac78ab26e5fc2b6c472d03c3e24df60c3bd3f80887f76a00493e155f7e9afa6a367a16b354988c9af5ef7993815976dfac54ac09b431ca439cdbed1778962f81364919cf8259ecd62ba31cafe83436390a703d49eb322c4936bb637e4cfc6de4f9db59468f5afd2f1ad7243f051c776d2b05d4b5fa441a9c5a0baed77119f1c894e6b425d837c5fa0ff403d4c1ff95275502a5394c9a6d6597f5524879b64321056fdbf46d58e4ceeaae2032390729e38a47c3ee74b5030995a866cdc7c1a57dfb201def11bbf6b4af16e2fb1cb339c9ef0aee7391a2646869e7df386a4e30d8367cc37ba64c1ce48caf1f39a69656ddb64fe5e66c0f5098311e8c3ff5cfbe84466d7e351681c0134b20fe2e8838372ca5e49f207e6c2c6187e0fb1d4b08847cc0048d8770a3502da1d114fb8b5a182877d61ffa237e08a41b8d7b7cb79006cfbb1950591a79892d62090a56d83d5be67d54593e52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hff2281160e8fb634a432c92900ac62e172d2891163e390fcd26f908df153c3f3d933d6c6c378c3437d94f835b02eff191d5388419b501d98274daa9b3760ed131357cc71aab22d4e2fcd07fc2983c2f90f30e9aae339e1ce53cafab1696544adf33e3848996704a8ea5cb3e6b8bd9b24e3484d7312b8c76b1ab879830a61f8f719ae2fbbd3b0c06c765505c20923b068435738975eed262b93d8534a614b753bc59b21428ae6e99288af2828c266011614c43d281a4236b867f43dd9091187f184a3ee2a32d99246e4204624350a1171c7bde769b8d058b32061e7171c96ffd3ac278d4615ecbdeeec824ac0c711bf79984ec8def6b254913ecadaf7e1fb685d5237a2376373d6f701e54a070097ffe1280d7ae59e6ae574b54ca16805474201ef97720c93d0f5df0147949020a3e9eff23b8ef2e063f80b1cda566a02720959082146ef63e2718eaad4b8ef9928dd0bdc6b05c0fec7e4417f05be024c17ae2a08918d3918edda0eac11b2d3d367ed1619823886de57ed0b05bf18da0de193da0671f7b687631699af9a790480c4929109f2643d3acd835246572fb88948fb1164665dd644395e14101475a73cbb2f28a92c9be2ea3a71863fcacc40c103488ef0682835f90f9d1ab2a06bb7dcf25b967dac86e00c65109f0d104ac22efd0891da936cbf82a302ecea9d73ff11884da1f0100560447e3257e957f6def0684f75cdc428ff4a46ed0499c565326507ab99c8f6525ca2990d253ee570099c8779525c3768a24cfd4fc5e05111bd1ab3bb1d2d41c5f3d053e65cf9b51e61cae1fa135afd7a1386f35af695589c39990f8515048b4f7a270a26761a4272034cc165e72f05f075d71950c806e2baff8d1e5e83445a8f75a8ec5a53a244eafe45e3e6d9f6e98035bf5fd5a8e78aea033b342324cad399c0d9943ebd9ad73f08ae17d69e01c7406f303494cfe0cedfd9541ebf50f26a6ff838534d3e284f3b7f543ad0cdce6c714a5bd6bf2b2c148f5b196e251cd581763da1007601e05b554b7079b395fd40a3abb57633933feb67fbd054f1ac676d4845a02bfb4af52d95252ca0d5b4bd7508c7190565f5e9ed255422f284ca8ff6cc5a6607c233efec19800d33a66e8b472581c0f60cefa4b6c33980a178392e2c15be05fbcbccf9d7f3a2089afa9323f542952f87e2c4a40e2c21a118d759d7afb128d5f6dba81c22c45767d45767ddea32b75ff1159148ca32891b6f1c4967d68111342592be2006256640dc9d087547d8ea512185863487fe78622f0157f255e0587a167592d8ebc5e591c63ebab55e22a527dab79af33c85fdde0cf09dec27b4d91f4eb962a7edce58dee1b07484297f916ef2bff761f5219178d4d02d0a1ade5944461aff6865f8a70388a4011aa299e0574edb0ed60f704edf3d0e5c9f9723437dc6819f612035244af2cd06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcbf2fcfea5f4d8fe8270bfdcde5aba3a42ee33c2e5d905a072951a433ed850a3435bdeb55b95e7a8177ff48fc7ccddca51a2f4f7968a15b3a8da17924f8d6d19bd206b06d18a4265ca84082b4018a275ee0c32ad1524d87c1806abe6cba36a87ce4284d007e3e2d155dff06f19c32d9b4207792f333fa09bd79f477403fda2b259a0a16306713e43d639e81f9473dc1eb3e4bca5aa9b80204f045c117f32336c726007eab27f5f6a06a6a96bb02ce0a23880ee445f1cf0781a533b40a1fe9f13f81e641e7802c6c47bc5d5a94afd3138da15c0cf67ec25b5bca03bb104d762a273b7b0afe1ae5126da2485e94657a9e42f74dfa0c5ab0701aa9fb1192e7684f5ae365c581cd7cd14e5f04afe37de3ff428a1792838f3b66bf5ae45c925808b7a7c766958b52db9194a92558bbc531c3558ea8194219b7cd75f69ad27f403e0458b80d0b6c2625da77353cb04dab558ff66d0fdadfeaa1c6386b8bb2afb768d40b855349f95c082d719e551b5ffcac59178a5efccb9be8dedef9f56c76ded635333881920a6b7e2da52cf35b62705b991606b62ed21ca8a07a497c84c6d366b8013de1976d4bd6ea264dc47fc72898be97705f0754b16cf1da118abd02cb9e57a1ef46a9ce0a9609a198cc43f9b2fff8b681ea58ee22053f1d934c62ffd4d9d2b8c75ff4ee0033279d61c58dbf186be5b12d353f05085d14726686144a38dffb04cef1a860345689b855b466b20e71b03f9c57b5a317daa1deb062b8e9d84a805ab87518c9202dd2bf7e588a2e6134ff02b3b24ea8f037728edd12bd5237a62801d1767b190953a5f9f75167fd7549a1cebe2baf1cc9831348751ab0f869dba44f1d6f60f151101a65fc34f4012047fdfa3348b5c66537c98bec9d8ac2124b7347a416c3697ffe800ab98a776fda1bf58f2625f925d950ed2abdcb429c9e90932b240cb7368c91a9cd0ab3763b0e4cc2bf0d4f0e330493ee9b9a405b3175a0177726fdfb05fc4f69ec6e9352312994a718cd17f2fb80d0ffd1c31fed546e4d1e553b430da6674952bfe0b38b4d35dc5f4d5f16641ffa6e5364d004dc2f0daa421b85b91a1e2a239550b29348e8f19a846e775b4cfb3d460e6dcaea1736ffbca2d60a20ae0bafe0acce49f55bbd158dc043f18fb28668980efdfed1e8566e30c96ad521649e954296342f7b69e694361f0c32d3630d0dfe4963c035cba3061b588e43d82b84b484dc0728fadae68ca18292aced8730f83148b35676e6d040992a70ac1836bd4d840c0214cb2d5ecff19315b20476c38326f86239541035bc7eec9c02e6b7713057b476ea3244ed00cbfd0ab682ae5c9c608f84df5a76bd4ae4aeef9485d70c8e131949a2087447b64a22b7d7e742c654e117afe351f75612b8ae70bddb34603b935e15a2f46a21d4a39fdde587c9d948208196a95e16b0464a655;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf1d8618f407c4d4ef1f011723b8cb64b1c47bd52d430f652083782f5c668fae3df8e8bbcfef613b476136bf040f835c6758b3e2e0ccbb7cad6821518fec4c298d44386506a67fbe4bca8e20752b1429769d5330271ea4d847f0446f11bbf7c1d4e5ac42bba4be869e6679186ea8522651b3088959727631e5b5648ed5f6176ebafbb8f7eaea4b4ef43fb730b24b73b4704d3fb442a065b6d940e52c6a71815251244f77cb46916d3e4c89316af9bad8a0d2e320071b2975d78e67fc8ef431d23b7a612e55438b2e367b80161c28860f6accaedf0398c869cf79715bc3ab1e1036855f980089582e3c95a3320dbc3c1a7b6b7663b88fd031aae8ab535263d1050b3d1edf18c6abef1ccb5f2923a02beecd8fc15da9d109ff00f8f05e501f32860b72c51b84547760f04a629131f64f4a4154fffbe16a8f149e9e13ad3bcc8f4fa038ce646f6ca0eeb8e5113c13f95658cc20e49901b414bbcf25ff0c32ab007d8803741bb1f03ba33d5c73c5dbad138deeea32efadb8693c83c4d5dd44dac5769faaaa72384ddde0c29534b991c4d8b37af050a92b19e0d9ce06a9c8386b70ab028ad9e9c2067016618dae5753ee4992846c7d2bb04d191599da54d20832b19ee7c8772f2952f11e2fdf7fed329e6f612173240a6c66326da59dff857c0b97b0bcbe583c2045daa7f74e3d3e7219dabca266ca1c21b057f9a9a6d10db09dbc05a176caae61f38d293bb5bb9ca13539c135536227e7e70e1e2406041afeada9ff77adbd676fec31e586683e38dd8c71ed3faec479a3ce1aeef779a49bafb5417d07e26e1c9a408f0d6acc32088064c8f5bdf01a5516667a3c6cda97de4ca6dca51ce658f5ca814c44bee6dfd6347aa79313dfe7691254c9a4cb6e5d5c8b7bf78b65af97757b78f73f3ab0f178074b77c7bd8ed32acefe8c6991e3b8c414cc392221909a1d572da50b70946fbde487ff187329591116c50110c0ef77342249856c3f6e04254ea7a6ec183168be67c87503f43321195cb990161b50b41cd06cc304768c6312cee22b7290f1193448b68e99904ff5865b208875ed3439e8c9a473bc0f89aa246f2da2e337001d6c0aba64bb32e99b6bc0d47ea3cebeb6f2788c6393e4db2dd53576d514fe4d2d40ee12e65b374cc758dfc665fea5869ac5f81a289568d5f4973f82347e435b69d271d8c9e5ab574a89fd50c3ebf6332b2e11021a62e119dbe0980cd97635757857daa71973d806772afec8933305fcf14c5c6f35ec9c7f5b3184e9d9ae0e209f8e51b3f68f7cac1046431d55a0a3c48f3b82808d42918bd8ffde16372e91e52e0ba8190ea107ce37fc22aa4561157fb0366b5de585ca822cda912a3bce0b44234c928cc7bdceda3ac5bf4d826be147043b5698c32673d133568331a611adbd0ddf8e80c8250a738e3b47ff32de482c45a5d09b72a72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h18a320ac67d8b707089354defda25e9f1f35430952a49ee4d32f31190871a0e0b975f2c78c3dbc1eba9bde4d74add5a931c4eb95a6230db28c485f1a49b34dc4e740d6f4393b16efab82e9a3fb74708af8866afc35ef09e886c9a34ccd353cbf9ce923cf748544a19fdb4dbed5b521f53d9bd0cd5b6fba6a277313eecda510c1654a9a4badec2822a272e2bb1378930f31a0129f7fd47623d521e1f1c4dfeb49e9676012690cabbcfe91c8938fed11f5700561ed5d6d4a3142af1b8d1e1f4d60256f079ed4ca0842da3e7b367b7f41e133baec2557c206e8158a8fa6c6e79c3eaf0e4ea7b1b281b9b2f018de552d6184d0341cc79d8d0c6e59f5e982188e4808e90ba1a20e90e83ff64c58645566bdceafde8fe3f1ce4d6f63185c7d7d8c4a936fbda0d8d73f9a44debe1d55897f2fe00885975eeff6f20148ce39f9b196e935336b27bdefa53aea000ecdadb615f6c633f5ca13213fbf98a35af0b60d16fb6394593e54f217aecd63645638d00d3b42b8b1ac36288129d9f91d5fba50858bb02011d4dd7449fc804f2ca12f35e3decc705a4def1ceb3bd29fdc9539cce0fad04b47fb03948038d5b36d2b2b83b9d9f87cbdea93b2f6afda1719263f70bcc761f45a1296eedb3800870a4b96694872a4d1f6c74bdabb38db44ffa99c5a6d108a57aea1e2e77a774ae64fce28e9d5008d3f0407753077e816f4aaec00cd2ec6e576a72a4e61f0a10342d8d5b7c5f9d92335dc68f0883282435946bf4cf2acadd23e3f206e41f95f92af49803b7b3ce8d79b17a643bbf67042a8a754a98159cf18aae19b7ce12ce57ce7520334b6a6be13b2156f7c7b18dae6a0b3bbac74592c909f1daf75f39d429bc300d3fe4dfa2e8c06a556f86340969b508e310b0f120a37b872c12be0bb5c8c266ae74e228954edea172a25081a58c3bb480949b1b27378c909a9006a19c8e08fe8bdc7bf39d60093df815ace870ed027ecd14cd5ec884255565a8704b85cd355e3fb5d1881b30d3820a8fbf6d11c9af45f822150d903b634dee8be3fdeebf333f45b7fdfa510af4ab1ecf6eec7fafdbdf5acb3e0041fd26752193b436b0ab56fc66be57a4ab5abcbaaf8964df0111bf6715c418f783ef55f354aac8673585789a5dd4d167e2e2c086c46136a969765ffdd9a5d03ac15e9622c1d7679bcf923e7f16a86fe8576262c23aebdf8e1719df135ad9a827c7cee4b61e95341bbf1ed0c251788ce51cefadf4a1ffc2910ee73b6dd6fc1b52b1b8459da7a1f0b4146f0b7651174c7fae60c7c0834971c1251255f8841750f02d5101e9604bf3ca19946bc38f7c79e13f576ec685b1b2bcc36caab2b561546c07be04685c734608ffcbd352ce7c65f8430a8db92702c5449eb0eb5628c98b2a8b2d0a570760800ab5f7732eda15961a67e23185fefc5180e4eab09c517c0614a2f0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h843394ec9580871b2191e1ffb9ff6d00295e66fc7a6cd03f64bacb2fe0b37610edee57b7a13f8bcbc8ff69b0ada1f85a1b0e73f6267972a3becbe90eaa228595f5c7e864d3758a7361678707c9ca067b184dd271b0d6bd812dc63433173a394266828e0098fcd39150fa60e80da476ceda9aa35cd3966dc3a967dc4ac159d80dd508f9e466d594e09d40edcf00c55e0c9cde4eaa9023cef62d11179127f8d63935f8a7f0814e842787a1d3ccc504bd89f1d880b72d9f1bb8ad1e088983ccf7aeee1d64863172383347a5e5e2eeb8256ab4d1400d05883a779fb12d21fa99cdbdaf75ce765314adc5bdb26b4c8a8e8f237d02e44b5a13df4e6f276faffd2f59cf046f5204ea39feaf40b6634964547307e43504249ffa54013977b5a7409d310a7e4c3a3491cc9632e9605423c7f0ad5d7c22caf695401b3bcf903bf180c6096915828c68879dabb69dab2a27d21d112b2fb6a726c80fb51b1bae16938503f61c30ca185871ae86bb9cfd1b67cbb4809f92950742b9a9ca2329658adc4df4f72acf0a36efde85c77977c7b89444061f41cfa1e76e59aa11c9dc50fca1006a4f7292b332b88c2da244b23633014964f324e1192e25c987044fe8cbe906b21b3523ef445d808c70ff76a042af8d2d502c89f77be08e9d2816fb8ab25cdde1cc3a2b725a247bf8f5930bca2df8ebe6b0d31e3dbae4e9c3118112aece6597d56c3eea7696748d9df619ccd1c642f24738580338ec6db352e403a6c76ba6b04c6ce15893cbbfd7551f9c37d5a8bdcaa18bd04b8afba6e162af1173f22c1b01b6dbaa3c31c19137c48afcb29ec08b397f303fadc025fa166aca9302171de6c925a633a98401ee137cb011fb191c27c643f23842d8928ce1955833f51b339711a2b8ff2d1f9c024086002fa1b9bea2fd60e57beb3b50fb20273a154914482525857a3c26d16ba3813e2cacece81c0f50b6cff2f540809d77bd3feaf5f8b2ab6e8a5542c0e0fc71b3b2c809a31c2067edb8e43640d56d85da77ffe713f6ca8cf3650ee68a02df02b10acfbbfead1b16b599317bffd72ae51d350cc9141335b7e8bad790213aba5d56ffe64a6edd4f9e0245c01145718fb037aea77e0b142146841540ea1c8745ec0dc22f45b3af822e21831376eb1244bde5f660a40bb1a9ebca0dbcd0f9ec5f1579e5ee7584c23509bc603f35478d961d913c260ebcf2d97420e37e9ded0434cb740e3255900abf7e76b4b17d6ef625bcbe9eed330e5658d8ad2af4142c36f2999e334ec55b42a58709d109fe883aae1564c78141274800e20b4abbe611d66492f4f1c5e8743dfcb85d2856092628b4a7954574532f7f4cd7b8870380707864934ac36996c055e3dd27496f7f7f467d598597e33f9dd8eee95f5fb6397c466c343a647aa84d5c6cbc70c5dc258eb3c6a91c2250126cb35741ddaba0f489;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4983a2e8e63fc0020ef46f15f63cfffaa7a451b134d4cbed4fe8eae14939dc02c5fc57783165c993ea7826bddfc5cf209f8bcfd32624935b8394b890ce2448b830feafa50e8cb405f720968de99c31796839cab497be101516c7ac3ba91f0bcf260198631d718dd865353ad4ac996202112a07ac896ce51ee799f30af74dab222f95c0e1a30ef4fc0b89c86e4d0574076443c84a6c3fa50a7efe836714015b38e54b08cdb1ff83c48d53af22bfa1bc0ca8859beab6dfbeb50853603157b4a1e2f22a0178c90d5cdedcb56e3fbb9f7041efe44b23ef1f9068eb8d32a446d09103e3d3a54987fbd61d894b086b24ef1875c6123724ac0d744feed77a74bd24ecc358953e4207643e7fb189a26a3ef96360bded9559383ddad3ee1ef7964912f9897d17e13f07cc1f207d8c4862b3ffdbed43d79570ed5ea74b248e9401bac3243b22e8985e1c1ba9a573b736fd0757f63ede405ce3be7834c616710ca256e101cf451b6d9538149362b27b64894d830c5a5ee48ffa7f591a8921be0269d68006cc8d6f66df77e2cdbf84a3560050c93873339895ba26ae08f29fea32177f58320da223a86142271103cf8d212c0aaa81c44595a97115f4a625d2d91a8934f39afa6bd99d2978b152721a4dd5f61eff5b9aa6894683539a54acaff328ef08121d173cebe57b26059578e70f9005d02e954f3a545ca7a16565633458088ba2b9c836c1a8721aadfb5bd82fdffe59fbfdd7569a4defa06b78f4f963feb84692db63d4922dc109f745fc4c0abc9238f228700e56111c5e71a07ef5cb477725ca0ebbc92def80b23001380c300bbf3ddd82762b0964ad6d6a5b65968ac20f209870a8d1c73f32b055ba504964e9c13a1b00383e0d3986694e9b1b6548351193b2abc587932121c6bf695181d8e7b230a3b52e306b2c4240fd23616e35fe72d6ef8516f1ae5f5070e82de383b7041312a242a3b463ce8407c152ec7591ef7712032137c506f6026cdac756b29e51c0aaf36feba767e336668fddb38f5b882d87c44f8b3237f34e7b21baa00d995c48e6e184b9a4568360c3e90d77e3188d7f1e88d7eebf41d67b67eb5ad45169c4b45fcfc81d06bcc182762cfef5b93c75dd42df4bc82a0d78b3870a277d52f2e320343a5877b7733cb3a269e8f91ec331d0b7dfe7477fc24f2708748b175d5af4f094f043b30e775b001e6ad9f875e567c18be735609c29bfa44566a64f00d4238e181269c3ab4e4bed3e135f528e5bff91d8e4cb34b41fabb9ca780bd243a19f7394ab01a23b1e97339435468897593c76b3363c998c5c5124af56bc3006f0a81334a33ef4b2ddd0262f965a9efdc6356651470e2ef11748fd540ed7eff5c591630f602d69548329b77981e94d21a726e0e41029208694f212060a83bf0d32178b479d760210b4fa433d4ec0d19cbdb37cb1b3622481;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3160ba2b98fa075280e5399605fbe627f94a75f681492b3e1659e2bdbe2547beba8ec22668a317a0f80fdbee3a71742cd412807316849041e04d2cc2df9bd46d67827e1343e5781cbf6449abda94be7bddb102f15fc58d36a8ee846f4cd56b1160393c6161f39e7ec40d03b4075a5e6cce3fc136246092b9595a7fb786784f5c05eb3a9bca4407fb74b9daef9e6c56f262cbdb1746d89fa0b4e2f529f79cfd778c8af87298eab6dee25004ca74a086264dcded098d5a3551592331305f2d6b2a3419c82f6584a37b086d9b50f9e117bc142c4a05691430f2560272180114776985b1e97f28a7c2e30fc5e71d42303d4920fade2e5a13bac4b5a423f75120601e0aa0158e3be6559e03b46d8bc97d7f84a68602c21ea4684e802cdac27c6f0429905e0165eb9c4c3e53af27e9483ec9033e258938d8edb990f754cccab42247dbf93f107b2ba09bcc29fa49fa99e4aac40342a7215f1f8ed83eadd00b848e52f1ded0571a6096b2f222b138bf9c8090507be3df9ef821ad89e02a1d1fd631c0276000c52b039bda1b7f5f18fa4216cbfb61b7323c75027c00f794ff579bc24cdaa5c995c730866629fdb2cd2caacbf59e5142ac6eeadbbe08f0109f6e5b26518412b2671997f67a4bce4fb21f24d1b8d1747e0fd76fc03e19d41ed709a5b07450d96fdb09aca7a0d86d148ddb9ca8ed8cf4891626a92fe134f2cb8c6f347bf00d2f7791163a75ff46822d2298e15db923629e5b79f5ea1d21e9d8ce700cb92b145a1c76695ea757c23b3d7280a243361c13e88b943e184c4166eaeffdad8fb7a0c03718f8bf99d90c79f15d73ba843ee3f3f021242f1204dbfd34e73564b751c2aff6de4d69f0dc6e9239cce712d59e800a78c5228ffcffb0fd505fd05585ac8522aba10ca12ac23c58396cc38bb30b219e5d10671233c71f739d61f4394453a11077c0aa4c2b57847d9b14f0b207b99552199f122e9ed0db5d6c1ff3e1da7083f188accef37475e9d00436f81b29a806ceadc690be2e229d38f69b32e6236f19675d2dfe2d7c7f7e392d5b9c69b6e328a789527b0b0f993aa7c18015068787f433475d830e674462ffe1571ba1050456a6cfa211263de150d725512485a7aee1d1af75f1f6dd2455795f19875ec11e94d2328fa9cadf9d7de4d98e467e325fc2d7f57035732776a9565ad7598ba66184adcd09e25ceb3615030912131d1a385bf697bc4e44b26e7816ac44a842ffcf448c371ab7d7302f359cc400af2bbdd4f3db794b10adb068b788ad1f196ac4bafc620ac9c5509b3fd8db1b88370f7b948ca814f8dd0fe357da8892aa8abc6a1e21212e9cd8f517a7a5eb155daf7375cd7124060b467bc255b567039ea05977c6347915a2c7257ecbe900746666207d323cc15dc3b685f440555e88591b1c551fcd85366432afd7a80144c30a704c99ce71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8fa7baed5aeaa09d21e871ed64d30b3819729682f659e8555be6e8a8d3bca02f431e055a73f25d7664ed04b6659118a5c35d4f710e557ad656a530ece28bc811b01aae138687c81f42120eb0bb5d09b1961adcf6250146bb7c8d27a019a7b0151962d229f096ba6af8728d2ed15f45c5f5aeac503bf4b2a196a2e33489dd4e0cdd279a7acc7dee13a8efce16a5c51e40769e12ae3443e183e16f524279be24ec08fb97bd97312c618881826e43c90875184291ae6c6607c83a3828b932de8a23c3bc7078fed476f612ccbcda95c949587eae6866aa1fe65b55490773608095a3a7ed3934c5f1b9829aeed77164362dbb55ac3812cdd0f424d23b6f8aba2984ec52fc8a8a37fe610f3544e86075ee2c1247e52f4662628e2536330176bc9d366b30027d8513a7594c9ddd97a1a2f0f11ee325399e3ae5d8d113ce671d88cba3063a986dd467ea69ecf3b7029502ef1879ad7b39986f27be4eecfadd3464a6ba32cb4eff2bd989bebd9f74828df54aaf4576f6920a34bcb56b2423ea089e3d78a8e51e7e49042ec521155792d30c8efa9080f64d3e35385b425b23f7aa0e4ffcb8ebf652c51cf263f051309e08705002217bf0a7c413124efb227aeecd1d88c231a439a1ecb12ed870e415f98810cee4c2f8f5b7302a506d4fde0def960088501d4223c4ebbc3f9484a904c8711828a1b5688d8d386666c13df438093f78af840a2ff4a608743fdc360788b342832224c80977a714edddb6df7ddcc1d000dd479773c400881da14f18bf7121d24ac3ffc07b779179f86837118aefadf383853936802af711974238065dd7e5f0713d16fb3b450e46b722ad8263eeefd9332b3506be4d4be142dd7a4f1cd2ce91187490a7462559996cd92290d6745231647bb829210a1e93caf772e251daf812ea97b055f5d3ec94322bbe9c153dd876cf15514b8d59dc138b6aeb194ed7b37079ee31bb0a4837fecd8e9d45cf098e67274c1602e72332af1acc9359866109fda4e2030cf8c0ae629bbb7ed13d19a23aa15fda92a730fccf17087c436363c9e03de3132917c5fe90a24ea2cb6f9311a9e278aae1febca3b84dc69ff0c796c7eb98bf67fd2eff47a02a960bd1cbd3ffcf0a725fabe13c8668032560de176510edcf37fa4eae75b4adeeab6867d870c601120080ceec9fb049b9922147cfe2b2abd3a383cf2112303688a4ca670befcacf461e08977538cb740cfdec9b94399868ac3bdd0597911e14d5024203ceb5b7b68bc08d64b64b4f7ac16aacf83b74fec16b79221f5105c97f03b39fb16cb2879bd7a2085ad0d90f5e08d66f16a3e14ab0eb2a8aca2c6a572b9b15fdbc86fe228518da0ca870108acff6a8031c98848997a702c83d5d207a3a1ca73512af9fdead8621789a1fa62a3e02110bc3af09e70e349e543d91d86ca49af62518e68a18035e34fe4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd3c6d9825276930b20697de9c0fd955a1378e43a0bfcdeaf39ba9668cb6ea39d9d1767b54d98f2b8f2fb349018b28b1381fb0b848b37131b1b701641b4dcad4f14429c6ece2b358ed0a1c8883308521afcaf2a9dcdc36c7441b333435c3134baf0b145aee9b0c9830be196742b1b171a729cd15e76ea5013ca2d13c33392dbd3665c38c23ec72c01b8421dcbcc78470476117eb2bbdc1a1382c50c8ef4cfa196b932143257b53124e2713868247ace8dcf0f3583b808a14794eb1ccbd28d06b8d489ab2ce71f139352e88bd65e87d5cd8b63db69176a0c44c55d1eb46460f8c9784a022d37b4df74fb8ebd7161b1279786b28b70a341622bd623075fc142e5ca741a63f590b3ea2b96b640bfbfc404bf14a0a33477dfc6258285fc7844b69e34f21d00d6296f42c8f704d0b70bcc186daee70829b9823c577108aab6a8fd6369cea77ba91659867aae37fb602776833f9032f5dcf717315418f0a5bb85a66f3c6ca47d70948264eab7f32ebc874e90c6f34b56c145ed8c7520dca598078e46f63443f12b1749517a0a79393261bc9ac5576e24e5438a99e8798d6138bb9a66e11b751d7e15988d43bbf5589c9b106aa8731a882523aea4de909c1882af5956445bd83fad1ebe47b37a9474ea28ae716d814012552d5ea987ff5e8c6d1cbbe0f12f20c2f8659aced7519eaf6c60f91629382c6010c44c6a0b66636df00e123e8f8bab7b6d1c0d457ec039532825136ffcc21065c17f6c93ffa6c0e52c5e58f85e2996e449fbbda86c3f9d167bb956f29c6927342210fc9c6177122d7ff4715d9a147d56bf36095495feccaf7233e717a4acda11a859b1222078fb3179e4496481b1db2cc89d216b26c43331f8fb6a7106bbbafb5e9d370fad40ad1c4f339a0c01f7656ae26ad8a5b02ec58d33485c68507aa6d227fe893bd47288f1664d73aafb7713414e9754f7aaaa1121276f7f579f008c03f760f58be375700e3b13e2729f7e5cdd440671f87417cc01a1dc90c5c037d14946931877b54fff8c3b82ff15f9d6aed1a74c48cf1c5000f168a6002d33739ab1f4a38c9369e5f002239ba19d84077d98bfc56a128153e9b414a5badc217b1a6e68c4a1a179d64195e73a72c9853d40f7c4a57b652219e3cdcecd97f007cff0562348ac5299675a64cb3d68794e411d9a177dc40a974e6bc3fd566119f8fd30214c14f7f60b53bd8d578d20ca3d2199903b2fdaa487e842b70fe7bc7c52a0d2300d7e693ba6ffb59144fde5f9a3508cd8eb3ba7fee383ec56fa4e88f60e87afe1946c56adc6cbbb6b7aa9944915b9e7132f18d62742b8b0cfe505d4f3e170b934ba9d65ffe11bd48c72dcb1549a86816d6e282904889c79dd62096d0b3ec6bcd4ba2e4c126380fd755dce837f83ea80c1bd80a2010768329b5e9dda2569c505a43dbaa771f5f770c7359bc58679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4f2542b78d1be7e1de2c33fec585b811829ed84ffd9175ec0c9f419e734988e521f3cc8e5ae03ed46e7d433cf950fed2d646afd782324c40e5e0f4483efce30fe287c12f36829f95b4aa91910816919d7b8c963e87a3d631b08b130b117265a607ab8627c979572edcefa2cf4e1a3dcf2d4bdf97e48ca0ec9016d17bb119be2011c9195083a439c0bba33c14a520793aa93c97b453c7b15f40f786681165d755d60c0e45fb1e92c0d52fabf858d728fd6655eaec489cae12f65dd34816e75d6d3624b7840ec9adcdeb07181a43bce9413118056c49e3e1bd656508af931bc17b468eafde99c40190c51b21742f5e310a7664815942790184d338960f2e18373b93c0d1c0eec9e7c4ea0f26b0de101b2133cbd0597ab14b4a9b6a3134987b4f13c84e44c78aa21be9f617592618fd6ff197fcbde8cec5c283ac5d3a20301bce59a806b089b1b169b6f5950bb4f4ff6193be1d6580e3f1515c28cb86bde96a641a15ea125f26d7beb1c955aefd7c8e2cafa11291b3c92f8b163ea536e323ebe9d0c2bd4078e82b8042ec499aa4eea8dd43f30f00884dd509e15a0700e571a1c0c595f86d31c43b042d0678c8b91bce1f244a419b20831021f6b01e4dcf78f3dcb1e050e1175135673b0f5e35628a5055071f4da04eee4e085c3f5ee934d5ce0d419f3ecf6f1f032fec54fb39083c8524bab2a37d652b24474f765c7c9f9426dd040450f1dba36d2cb216664e652f8451f869ef8f1322b9937497a795ab53bb11464ded8607b9d2f05eea6703c374f7db8c8f81e29d67f3bba652b1cec624ab181f80ecb96833f45942092577a0d240ea3a4b9c25f2b3f9fc384ab9111beeda54550fad2da991a47396feeebc14e1de7b6714127b6060b7cccd8fea03e12ed9666a16b48663aec712bb2c44f5f06fd790240ef6da4f4dc4ba0b18f151ce9c5b388bbb1c281f937ccf0b19c4bc4de8a69c275077b82fe54f8bd6c3788fda142ad0e9a704749bf327fbf1e91ae3d608e73db7e9e8ab9a74cdbc66905c1a970dfa7815cee700bfe9d82f2fc14aeb0c39dd0cfda87658df4be2517724c8a0f4a5f2012c531919172c17cdf537833c2a6734ba01223ccc720c430be53d0f94311ea6890b1f74d7877ff82d17830bc881f60474ed0706b9503da5a2743e3da4e11081f38da04582feedb2bb315c0780935f047f50c212bdfb531c73b6528e39ec0278cf3f89549d26a2b8d6ef07d2bf0ae5e98f2d748770f08568ba28ec6573a9bcfd430f7b9bd220a6fd1a9c614095c0cfecbbd3d51c21a3dcd20a8398aa0831269214e47af62bec7c5619008eac1296a9cba1107e4b351377c7f2dc714687415947c4811d7de09728388ab1391ab64a9a21f0d93e3df47dbc7b51188e310267fdc55d67a6c108cac3144b7bbbb9ee628336c2cc3d8a643263dcc330ba84f49ae072c98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h53929dc879c83cce35abe139b162d9c553bdb2b8f53367fa8aedf7a554779101de6acdd0e1ef380d4c1f10ff76f2ae69b306cf51492a837d187b09f78264d85b74b09f3a62c8061083defe0c81eb4a13e43b4fba9fc48caaa16cf287d060b9ebe82b99e9938e440233ff53793564f4c7a600dd43eddf27f6419448ebb6f1d5865a260d8429c1127b0ac1551583515b9287563e948399edc5cac173f784ebf92d6acd71ad66c5e735ab2e3dd8a33857e08e99fec3ba9b736040367a1dd67f8738704340051a82faa026e91b5a1b123776310655379cb2a02b494b8316d533c197a3c9b24b271ba876eeab8c7698811f2ff1cdd35eba265a27c0bb4fbff74eea785df593edb1d7a5bcb951e1526a5f865ef72ef9934c7a81dbbad729e5e30e38eef4bdeac87ebb1d490a2d01b4fca813039cd448e07da9dc423e9de4081b91c13017d2359f0ebfadc1851ec5fd16b0295c00a9f00b2a2944dd3cfc388cfb54723462af1173179c65a52e46db85d69e491bb02d8dee5140516a8e40ab1b16b10f5cb9f8f67a5378c3f623f798518b4282d7ae4ac0570244e73d0cc75fee5f9e7b4293bb994844fcd1907eff442801699958651d0fc5c2987a7fd2b26f365005afdaa099f4501e0673c14930dbdf4bc65d727397757cadd448f0f680340a0f7baaafa6738cb15ac7b5da7c18d9fe5b8ded99caed38a9806f0af30781912125bef47637d05a847eb79f430de4aca2a307af9c489858f74b7540c04aaf97084a69ccc5e8b347a7b134e3f6617ae3e52cbeb68e0b9a0e84f30e218f3f7eb5f58a765e5990d371ee334af7748aaf60635fccab59a61eb15a9f2e4e46cb32c69600fdb53fc27a03cb9b6e604df9f580582dbf55b3ae7ce9e952ffee772459038fabeddb491f0ecd21450fcf2f64c413d127c469702baba3ea193bf19d70bad75dd7afcc62c112841cc424c7560b897dfe01883d715607e49fa835d6b3a84f21d9a83dbbac58c9cffa754bd1a4b69fdfdc2aead57d2039ae4b6f83b7b0d7877cdae7cc27483a24cc04dc8154d49ac4c945d7027ea187d34aa31f4a9cb8f5325e800b3747ddbeeda0fed9bb04d3e66fe178fee9bc49d85ee3cd18f3af35a62f9d3aa8ce4885e1e20758ec0e4e3f34fba8248d6a7e31c1a0ab783f6dcba77849020bff418266021a59a79b55012ca5d91d106575c51cc2754714076a5508570ca02d994545d07ddcd5a28a174f16a8cbb4be643e3722d02b411909129a26894ea7c8a8fcfd0682660ceba02833379cea94dcef41c37c6ae017430ee467fe0c5616405cf37930f8b42ea773a93208a4a1f2488e2ff95f096ef49aad7ec4ef185eb54eb41b3c1e1eda92697e3cf0330fe965ffaed260879144c3fb49d7854e92ca805d554cd90d1680956484bf4e2ad74f544280b304519ca833499d1377262eeee74e9221e573;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hee2c15c7bcfcbdc8aa1742e4357df4c7cc5697371483850517b6e220641404d408c9f195ba83b2a4b72336b2c1f75e7faa933ad7b7c3c4d6a1b5cf098394588f2d322d79cd34a12888fe48cd725254f0f00334e683f958b40bca1b4f85f73081d62821b0d1aed516070259b540721bce523ccc1f4541868f667f5c8598365e42544ce280762767d76b22d0f8dfb47e2c97b35ee60051f76279b3242cc0e4c2c8e4538db6054e96e65ff4bee181a3f7713a5fd94815321ba32a8bfd4c37f5af4442ed367bc24541cba20573ca8c82751d7ec980d32e404053a1afa8dfacca22b45b08da1a1a92ad3793269985409feb8cf27a373a145b21ec9c109b5e0359ab2b49b3dca9b73cd35a5fb3c685b28302067db5a224fd7ea332b23a827f4e94bf4ce37884eb9724e1cc1b9458a73637facb9688bfc47e7e13f684430dabc9c2cf6291f0cf93feb7c382d47053a923c30493f8dfeb6c97ef8946b716e701c54fb4aa2794fa1ea181923a769234b14be1c3c7d13e2188941ae39c1304f3d47526b8c4e522518f41e7a55a9cd8f04b744639f843ad6a6b7e79af8f40146439308a3474a89084e006c7127a7db42be72c0fc66a4599b62a8ce7e482c426c30f7e23b647c0b16c17c1f9d4c0db8fb8e4ffd041cbe7d3ea4df97f7fff3548ff921aaa774196882b744f1252714049c296434e3ea1503f1e360078bbf233a40713411e4cdc1f10c80ab4b67095f22c55bed35836bb1d0476e54472f9b0f19063134db9598d5dbf2c908c08b525a98a3a834891d512b6372440155cb7cf19fdb0e4827c0aa7e7882bea206f8ebd9919590ae35504658b494227c80507ae376e1a4f0e29eca47a96390e7d2dc1c23f3cd6380434521545fd23cf2b5c321101d53f479edbf850ec5a271f04cd097df0eeeeec0a80e3ea7f00f7a02ef558a531020cfc50ecd4d5421c4f5e1e4b40cb91ec7fab8d9702627d9af550d38b2a617dfd36faf85504b039d99726b7741e76d4945fd4f1d41fbe371f98b4d643ccbc59e39de83211365f8cb56813c4b2707927174617d8fb5c643357d7b60f6f52207b74310b865f70acf44aaa75f4a2f7ece02c37bba0810ebebb124c3e6e08188da91944ada8e081774f4bb071bc8713cddc5a5c209c4b29f5808223aed39934313fe66378a8fe40b7e297c28eee5eca367e8038ea56dc6def0996d6c75c52d57b850182dc24d1bf982c9b2cce9572932d3cca23f60fb6743af392ef57e10c1b3af50d755fc87dffd4407f4f1c299cc5ee3422c577fdc9f55bb14bf7e849c42674c6d1eede10cd8a31adda5e13c2a7b065ccfe0b2b1d85510d77b1edbd3dbf69a4e97fef8bb1089544b85c4d04c79aa2f672ace54816285b8214f44f78a18f585dfd31d5d9eb161e9d264572f6ca6348825212e119b397b49145317a2056c64262a046088f5167329d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h51e1515348210718711f911ac94f5532148f403e91ca4208af5c2415bc8933047469f4586cab45a7da96e49878ac7dc5c4363ca529f4c6502ab23697e6870ecdcaf5267351b72dcaf6a2c561c8cf09fbd73dd1ca8b86c5e7fbd043a89e8e7529680d41ad654d8505547eea410fafd9e7a2d858b4d2977092650b39164e3460e2e090df7781402a45925f9b88d6ce3f6ab7119a4137440370ca93bbe153346ab0925a64e2020ba4672caff2ccb68ab552d1aea3fc70a640a916b13c795840822f5a60bd4e86c2ee0ef12519bed96e9555264ee9734c41b2d033942e0322ebaad4f23c6e348cf53838ea589175cd6a24367186985d7a2a8d6c6baff379500eca33fe234f26327e3d0db7eceab68c1d3ea2b9fb41c5af6155f2d6688cbedfb77265de3d0c93b3a3409410284536c4cca25904d1afc6c754644af64204d55c7f84ef1360f47aee6f8f0d2fa42da1e1b0d99f63af0c6ba87ad9677edd67a83c63f8fe2103ab119fa94d6b873f4486eb02c83d04ee5d037e9953333eeeabf3fefdca3baa30a9c6abf7f4df3f5c0e4a2fb50b0e65ad29709cba94ca81aea5edab3423cc5ad0ac3a7a3b64d7d5b3b70be96213b9d4234b1451ced2b1fe43f00ade4030a28ff37b6da81a1ff1a2e1cc13649f6722e9dfaa8afb609f851d693a05ff9b94877994be787cf205c56ca68102c636589f52eea999c8ebbd0db8d347500ce7bc0a6c53f60a0f7e3594479948f07f8dea86a898bfbf37aa44398e027d297972c0e7092034e236510238afc58d66e3317b892370d66bc9fa98a13c7351ad01fbc6ec846a9df1503dc300ec487a3202102ffc04b52b32e97377e9d9bbfa5110a9af58567df4b97a38b02709ab72154671b8375c6b714590bb3047793cf934d5ddb12c7abcb71b6dafe9143d9ba1762d957a610da5189581309837858e6921f6e0f3a2e9ad69990e9230b68719a52c94228da99d2818e0ce033188740b1400390d44e38c4936ff951897f628e0670a590bd370bde6542bf204aa2335501d241bd6345f3c9a7c78309ad16f0cd4e0e6d05110501decc8468d2df7a6a48e8f2a1195af750c8946077e2e21a27f1a13e774944be7763343333c8864859f58c97f97a1c3a14d27ecebdda8e167df09911fb8cede1dec17d39c2bd359c0c386d216116fcab73fce2e9d1ab1e3f9826b9b28a5a32618b40d40db87708fa3f566d0647c178074c43408f30cd8e4072b2fd34944eebcdf2e7b967b21ebc1f2299ea41606ecf52b9c794a04ab65a5d33398074277525d78b72863d450cba483b9970652e6e92f2e3cb161031018980ac90fb39df00102e7330f90ae34604731ce9e71cf88bec0d0d39f9a1f65bfda638afcb298ce34489a1cc6c9afd4ca7543f9f1f8c2082ac5b898742e7bf49550246c06731d7cefd619c30bcf8d84cd50268df794751c424498;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h85faecd1cdc6c81466435593539fd7d15d88937c78db86d7a478b8198dd07b9ad9e1b7b97e73ec188e84f2ae5f8ef1aff055b6d6db5ac8d936059408b2874b2633bca318e53cb2b2818f90e2d2ba0e1e819106ab71f9cb8364842e4fed23e9feeb155b0bd0b0436b7d1798adcb0e9451988f9808f8a9293c7300650ba0632e1b05b459f1294d1cbe01fb20370c65eb69e9e06add542b8b518a0f727aec0baa1b366ad0c4a6f4ea64cc196e65693a1faca0a87091550132be84bc92e2c64152af65c4d2712916483ea725ce82e716097a876bcc6fccf933e0e11f2f2101f1d2254e2fb17438043a06880872805c0be0c6ee14ee3452a7b3caab9107cef0dcc59f3869ac473e12d1094fa523ab362988e3ed934b26d49127cbfb1991b9b4fccacede9c3e5bf41ec2ee40ec0e86fa59314f22470b79c3c247da9011a5e7000e8a7e2ec8fa1b95cf7a3803796c3ea9b2830eaa60ebf826f3cfef673b838f91df90173d50c267903d2d20e93ef10644622a9dc89b83902f6d061dbba10a42653abffecfc267ec1cdc232f52cf05ec0b0aed38ad82c47611f55446b0233b877002ad57ec02068abf9176ac8653f46b6dc76a64cc0485af513332bfb1fbb7e3ee44be0fd9c91d56e6fdd7801c259373b14504ab2ec92aa2e93a0d153cb4ac113039991f9358acc407ea3ad00bd522610472ed9a087df71517864966e9e4ffcba5d2a2d5d14aad62e20c2c01ed20f65d8e6dd78e0835ba210ab5a4ac65dd93de56fb6a7aeaba65290905c821277f4d2909f92b982faee48fc60c558a624e625811879f6a32ae8a0b09629fe1b9ffd5369cde9a2932d7717990858d664ba997812ba03659d96f056bd6ae37e363a88ae130420e6de6f2fb90974f769878b15019ea9fa5603d5ddba1666c9bb6b36fa7c791225e32080243daf5e2d3c7e4a0e80d3d709b869858a7dbd1a3efc26c0cb1c93e58ca857f208b371b74bea2348ead93dfbfdb6fd5ebbc0f0a59fca40df6e70b84a922cb593dd8e35be1c4ffe492454d3c82725e53740126f06849de912727d4fb25e2e320c0f3d084f0b41284657174efbc1ef4303d13dfa5f808b93c191940d82b888408b9c36e266274e0864d48a33d786ff0eaddf1ed3ab9d71715badb996ffca0d0f473cf5150e26a4f226ce7ff602dbe9baf1e045ba45858613bcb4e0c02bfaa8bf0c43534a1bc9152ae9547ed595ac42438555854aba5e0907398699c595f960e685869f52195bc929b60465fdf31a02b52a4a2a1017f8fe2bc775dc38920ea8d29ae575b8b409fd508bae2c9a3a4c052e3f6857ac3dda5a49c4cfda851706fa51fdab36f3f480676e07cd4b23cb28f9d27837b71c1d6ddcb4ae60edeacad0f486ee555ca7669d7b2cdc07ad52152f73e8acb28a7ebe92f3cf67c8e3b877220c9dc5555dbab216755af8f181ff6c70c24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfb9012168147be68ec130b171ed31c0d8c7200d0fdb05d3b57ccf79e5aef4e8cb64e99bc46ed33c0957b90bca1a7b491345a36c565d023a45e0328fcdb5b107a4e93ccea2859f366a21661be8c725edc08e2ada5f04639853a392790333718cde80710afd2729f96c6dfa83f53e3f6692f5b345422dda46242b7904b9c961ba2962367807bf4a1c8418d3bceec288bdf112bc78202c2661dc5985ec90321e43b9c4469f1a12a31d996ab3ce3585b394d9d8a8aa6a87c3a25ec9ed7e01bf632de2e8dd8a55d09f3ac4cfe3a038538a9311422ad480b123d4e1a524b5aa6801a14b4b6f41d058dc22025c92df106d4de302e6738ee29ed11021b37dbf3cda607503847d26450da53af77a24bbd2f1b663b4598ce63f0526e8013ea78c8dfdbc0c2087a25133a1e1a5f059209be2370d68ae0e0800a20063f955785fcfa149f4d83bee700e6f8a23e9adb9c3f31b09ee22b9c8d37ae1e0337c9d412ceb00361a36a432843c246a95f1276dee686beb96b719e2e54f011782a1da5a44a9d8c509cc666fefa8d978ab7b12393cc105b8331149021e964044492b52c4e711a11577b45a1d0eb56d08c74badce9530f7e6cecce81462f5856a13ec9d8977c64c096c394c0da92ac2f33251b66d7496dff3cca4bcb69e0749b057d67ebbc0bfceac530a62bc26b22ad63ebcfbddc52b1260e80eb4e0f84a88c1ba1870406b294841ed3850a2a452bb74c0c7dceff837da5892c73819141b47fae9d236dc51761aeace1a3184abe72cbd307e5b37be19c431ff66afd2d6761fd213d71b47e7193ffd5610bcbf8dab11fd174a85b1cfdf7f83b2eeb7fa4bee9e9e682373ce5f208e82c0d96ce964352509fc4b0ae54e5d28c0b5c8780118a876db8c3045b36e6dbbdba2ec4a420cd371cc42ced5b9e0a225f753387d1fd031add436316ce3f4f4c0447c23638e599c6e6a39f01f34e9e0fef2789282c376fc00999184b71c0a828073b2c7baa138084e78b043653a9df6e2964abbff6c990eaa841e24b13333562c644591adf476e8d2f56f2dbb98d4a3702f1af28ae9a6a4eb0329f428d68c9cdab715929f3362264b106b77df07b68c2e6d7eed4e4c2bec089095c9d006f230a16b408088e177ed284fc8549bdc01d7ef252958c21d390ea946a163919a0c968eef0626b23ee1bd152426fd95ce8e07b211deb38022a7321d2727b7910f515a6ca289a550ddb874af20c8253a2f8e8073cabdc0b3619ac5c4b862c9eb98862a361795f0881edb927dfb2b2ed3d19304b17b9b2b5439b26db19783a73c2eb7434d5c697b8f10a04538e0bb59bbab8b4ba4ff643657395ef5f5da85fd059765902522d813a8f2fd89e982231d1683f53cea5dcbd8c8dfe025c6c5898bde1b531f67c54c6d5ff0a85250393001fc80ec0a0d51393bd9d5eecf2f5d00d73bde3e8fea24f9c7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd447d3c8c3655cdc6d606e68c1a25b9d9193d79a52e12f9308c21711b8f2c9955637daafa90ffe80a6d6a08fb7580d646ac57df87169d93ed7e61b8e485854bfa862bba3e88d2ecd8246539b2a04ca88bba90ec8c6754d38267e6f6f1138ac27b3b6d688a8ea76c234acaeda34d5d51253a8fa501c9819a0b031924213261eb5e893f905ab6128c903769517543148006960069a9504b87b18fb54c8a0dbba39c93a1f7dad35dc7a5708d09c16ac154ea3cd01f1add88548d39ddebc5143cc44df0ec84cbf660dacb82a523a5f8b9c73d10aa37c42e28289e0c4684ed2c1324502c7aa8d5918efd4660f9918f08dd60c4859ddcae18e39cf0d993548eca4ae13e19412badcb37007b356c2f7ff113f1707bc4525d86d8a0dcaa10b5a18d6775d20e2f11e44830f3f81843abc5754765bf777e3ea2fdde8f29189d3bf61576272c009dcd26c46b9f5842451b2cd8175b3096c09d62098bd66fe3a4f6931f8058c44d32fbd86c4bc438942bd38c20eb28a42efce08a01f0d43e250b70379cd3b31009364fdee6ac34d83c5c5ece318f29b570c1a3e42e3cc9de14eb0ef50754c27dd095242c7bcbbe52f4f38100a17e87f97eaae48ba03a382971a8e3d5fcc7fded72b1c71c453161fb22ed64d0f14337c758ecd1d097e8f7a42592c8d7d235b42058ac9ddc761184b08163e834720ba4bf07b3b708dae31d751d499def3073f9a3ab7fb74e7899e9efd9180b5acebc91b0aa4735328ca8f88984e9ce32498dc4c17ddc1694e0faa3365cee0bd4ed6acd616d1423aafbeeeb4e31e399661fc1e2babed9186d741dcde1a1260d3660eaa30c612edf024a021fa7aa65c9b640f9874d394adc5bdafca1b1d73f382b33c323ec617f6e228cc8be72c27ab684bd828322e9c5f72c4e89418196aeb88e6da561fd94755b92621ca56faa06f89db5c9948a0bc82b4c3b20d795711e6d15e7ac56f9e8af4dc31fe3d65d16b3cf8a01d4eb4e085159987814089ac0bc40b17c49cd4e0c10590f88f3ca2269930b42811c8de8654c918236bb53311e119b78502530ebcb61d915eadd4f2079ab21701471a9c5c1a790969cd2acf2db3512a193bc3ab68e5014208c98af99313b7ede7b739187e00c8a12dd018063e5bdef6c42cc8ac1cdca667780c99204181207d6b9b21b755f87cc01441eb7846cfc536041739c359ef1f2eb5716807ec971ad1ac185d5f33aa6624dbc555586d0b4b7ec8741642154525cd76c2f877fce84c26ad4abc1158fb552acbf8b1e9b5fcce21180d0d2a73a4e58ca2b768052813143c2f7aafc27d26b80e20c2d39a8a0705ff3bde0586c91a4f853f74f365d45d51cc90367386e17b671057d4f27f73302c7938e75e8293032ca4f31ec345cfa99873cc766a68e0d2ac706a394fffcd4b8a9a6c6e45534c0ecdf30a571129ab52b6c38edd33c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h517bba6665c8b2066a5b9a52fb34253be947ae241bed592d3910eb7329b779f1e83be82a18f4b484c3935462fa9e2be3b259a0780df15eb462bf758d925c4b215828445c218d8cacd517ee6d92401a9e99b7218fc1a2b9a41a4a2355077c3fa60b42aa7e8397511331c14ae25672b0704f9d5ec351f129b755a610d4ce611af852ccaa3ccdd05b87ea54ff10875ace0603d2ed7a880981a214cd4b315102ac9ab9d8fc508696960e4808ea7601b7db947ad4b31c3f5dba7101dd31d77f9e1c18d116ec8268a28e96f0e8a2ad8a3ed7d32e680dac398b4e8ce09d32c459cdac6d2aa553f660ba6a37a980ffa174221f0adaa3e3585c97a1d0e4dd3afe4bac217c30cfb6668549686d8067955c0375d446e1f79cb5ff900898033a349ba55a71a63804af79bf0709815618795d1b6843ed1238b634950659446eb7f743f1921232db43649bd680d5abae48561296a7598683715065cc48a76e168c94909cbd763912a9772b554c94d174f92d69c731a865416232fb8326b403dbaf5f4d2ee55dbc69426bbcf177892f6e576c4756a69de521fa6f65f41390ea57bd6c5a3fb6a1225e230965ea3a1fd47091f86f78f46042b3361c47d76128d464ba75b2521be7494c18ee9ef5885859f18696d44f077245ec236da5fec61d4db46e993e5bded9a05011b5fe815dc0c391214c49b5f08a4e58f103cc5f7e190904e19ecb5747eea3a6dab05abd576008eaea8cff1f5e5b1fb9b3e742ae54f47da3028cd8304eb6a6db3e55368140896aa38def33e4557e3eca53f9d3dbe25957ed21a3e69f4c72864e256b4736aa204b3c4b79bed4dfd0d44b3b54c667d0c337d8ab83789d7d5adc1b7984331edbcd6553bfef5430f7d6325bd8f57047d4400f896b38af6b81bc949ae0d26fda1f9d9d21afc22398b014a0eb1f800652f90824df44d5482d527a2b75b85f95c5fe5f6b1f4cb355aee074a2759bdd3e22a0d26508b7c9ae3d71d374d54ed54520f019423b0ba039bf3ec7c46f5a3a40c5000981fe3cb9126ebab772559077c87772ea23384baa222da165fed8f881b33136704fb2780ecf798c8c181c0cba7bd185d0622729b18be1ef68173214e389c39b8763e7131faa7a63e377fa16f90d4798fc350c628c18004c4fe11ca8e0e7473b6152c5cc8dfcc6bc7360dbb888863de556d12271053b2f1afbdac58f7fe13ba715737a17177d991885453a6628d9ea9666e2c66e5b034cf02e6a720b01a8e48765e7f62f95cd668f3318a48b52b6901c1f893f83256b41b139eb7f0c0c191ddeb212217c0fae18c4c04d04e603945117c46a707a6b16a860d5e2ea10e5e134a5221da832836f60843a058fbbb1210f0172439903cab0f3952b7c798f62f85e46da522af6b2d108f1327f71bee66847bb1ed3a33ee1e51eff4973029bd94f84e397ae7dfbbd8fc5adadc6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h597eb6d5445a2806fec9497af67d19a2d4a0ddd855cdaaca8204721b6fab8b8bd44064bfd3498bb74a38ae38729e3c48af7bb955ed5013594f0b8582dcac14a7163881823a6e5d7b70c2ba87d951639739d192c1c6035a9310bbbae22fdcbb76d311a60fd2990443238fbaa5eca46a1445184ca3b252c886a8fb2905536bca98552e00f12c320f26f2900f648f7bb3d59bbedc48f79f435eda73362668b6175ef9d54404684750123a965986de535d699dc3f0d22c11e1301148ce91089fdb04b0a2d521b21a8162361e51ed9ca779daf707a9e2ccae45aeba56fc75867085bca2d2eb157242fe942e9b03f4d18c51be0d8d4e80f89ce7052da871609bb59ea1743bda8b2702ad39b69d61037d43d5389fb877a974405da4dda82f5ee1468c62b42d5b7659558c57fc6ea4b8697aac8cf3df7e024db0996575e47758498cdbed9473225761e05578ccd73b0ebc29b534b58ff2b7873eac524a6fcf62fe2626c2fd3f2e89c67ee28d366906686f93eda7f443863a99d99e3472a14a7ac17a5efc88b90e8e689456cebc543b963c5c2789434792992a8e3f78156c803ae9e37785a86a5af9f386194d2f4af35c0ce8806e1397f15d02e5bd5e437b0586c052d288e52f87a3fa3eaf5405c2a32d74cc870a04b73bffa972a124c3e1bc9c5eb8f1362394902c6a91f70677f7359c9c40f6b6ec3a282d8e8ee6e66dbbf933f6af66079a4da4932ca790f4a4b4c922359486a3735380305304cc09b6345b39172d2dd6a3d043a75d49244e5d4bdd61279272c8ab59ad1d8b3c5a63ce9365fceae5c6325aef54abef7f998db863bf3b33acff7c41d9a5f476db9a675d5b5f6c08d286f7658b9c68b52ac92d28d6e95ef628965398b8f097943dd0eda4a12c1cff291de7709812b6ba3db030b631dbe88b50e26c22363b5b02d043397f49cb52ed92f412a02d8427c1c5570be469bbf07fc6fb380d4e9994544ef56f7c61cd1b2adaf5359b0237a792db7bdeeb21193d86dc1537a3c441279ae75ab0ff2050d6d73485a56e49249c9387a788d29f890c81d89e949256f8c4ada0e71a19466cb03886fad404a43e6b5c229eecec40144dfda73858836f62712285ec97118055e52f72cbba486006bb084bdb07698bc8e31c989b2f9cba2bd698397cc610c363690ceb98af93374f66619fe2b8a08c254fe39de8373ac0f5f77b3c4863fe9878a19673a93bf74f8dc2c16fa5c370632d3cebc7247e0d2064ed5a56621f46e7100c51d3d7d49bb8593b7e534dad367ff9b70ee17c139213131047abe131bf48326f153bd185a7fe2cb638272b9dd4d88297b9610c3f9edeceed214e1dc85fb63c834501fff3296eca326467ebfe4866d0a92a1bf52a7be674761b750107c212543342fa481dd781fce3a5ad2d1773351f78cf898648999ce6086fb81dba9e1491db75047b54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h253d78b226e88178766b11efa381e57e7b1c94d940d4145134919a2d38e9c659542dca82ed6e7ed69137eafcfc4cd0e2dbfd3649dfa3475f1f76edf440b3f3b0fe48b58b26b93facf21cea74cdf0f30e2481f16dc311d3b6ea7f07ecca65b9f0794f842be505fa11373ce5a9e69d844a4c80e798966af2989aaec14776cc173c33d330e85846f86d702daa5df67e710b5f22bc21f9d3371fe69f2496b7f136daf1f05de50829f10d17b2316302c45c53347b5509aa2d9a92b5c4f2c3e4d2ef468d7d34edfb11adb91e890c68e6d9bb2b8bc2fff2a7499448948d44228f263da5954e097e1cf3956a4cd0a53c9d70be8d67a74b9adbb6ef3cc2fd036cee74bf13796690ad108b2f5d972a86081b0f7cd37a16191aa4f4eff675691b9e7f3b7e35fc4d42fda8acf031db05eee6f54f2e3e835889fe26fce42c61961c391f25698dc5c423d136512e8e0d7baaddb82ed2137392ea890aea7dcef31d3815b96e547217c0787a73770a678a8d36972ca834b4ed80c0a08d1a9cd96d367bb74b777b41827631a4532c307a83853d2f2f755b928a2f79902e648f8c330a54c6aa3c083877144c33e6e128f5fbb2f10e78e4df838b3dc9d538b32465fef4489371d1f5baf2bfe9a46f1f3107fdccd8429f2959c102692aedfef82d5f3df5176628d658012361e577beca5bc5c0fbe67256a499795f9d1119ceacf53094ca49fc83e3eca4d2b3e29bd03db56e07c4f0e0d7e0c25100f8c46252ca53de34fc3677bbd76f4df088f9b7c0baa192d8a41a0dd260ebc7a4d8bac4130f0bfaaceef631f9cc31d710c3c645d05f8c3452aa134e17f348b2aab23facf744a1b00a228f958520d227b9b611dac2a16e1c162cb639b74e486c0f1d1bc95877d0648608a9fd7e085d82b54416e49f2ee4904a4df73aa637dc9967f8bec0eb50118d0241dad27e2f531833049e884be74a7a47512cec2c7e149064bc304eee17bcdd4c4e5e9a0f7388b39322e48e4bf8a6070fa12425dc9fbb0ad47f5f697caa1976d4726e927cd79dcf57b53c69a44f86ae9a3990d500dba003275a003dd50f3a86c1f816824d495dbdb5aff802dc9a12e24433e769c2022d1e3beeac4d77cdeae4b649bd0fc0a98218978e7b975979c1a93a220aa1d4485a5f9c8400a77185109442a3471eb1237b94cd4588db9a08e9d2b4803fbaed38c19bac93d52cf9070ca72b29213e4091a093fb7808dd076bd294be273c994b6714b23a11c69fb31b677d3fa548b4fa5296ded2272e8caf3115a714434df3c981d0d1295cbca5f4bbde3c912e563973b933d39524a8ad82bee8cd0022207d0c8864e1cf414ad22cf6e0de0bc2ac48005c1278c9ec2aeb2c2e63a54c1b15f5a40dfaed4f05a8c031c553cec7a27d7b7bb77d174cee7cadda1ef503fca207b8b0a7619a94b0c00b08ad0230c488b711b2e0a3b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb6324c36c29933f1bf93041f23c4caa708334d52469f702f7c3477718cfb93163d8fb031df10abf115c752e56fcd8a26babbf0f8eb3ddc47ca2e482cba634111c57121dfc917d108a25ff43f2731236d4d5c846f8d264678a3644ac1d6db1bd02ec167eee524d5b6d03b87c7e769212930a5694ff6a8e34192f36124f1d20899f72e1c149bb6a211f6fa795c031fdbffb6f64b480359f4ab1c736a00da6c325e36729beb8360ae51e5e2afea0e973c08b0f8dec800d0674ee0162ee88327ef41b58087b5d6062f9e5dade489e9f6b87dfe1b30945936ba38a2a66613e3fe4b4dac378b05f2ea97a79ebe2625ba70ed2793b4cca937459fe1f69c7f48e499dcff7ce0892d20fb898cbab4bc1b27459c1154a4d9e8749272fbb2b8077a478ddf06a3d941a47929cc6da91478bf9f52ec1e52e47843957986387b7d63670248008ede6afdc01e2fd4c92250cf426367402cd440ff00f01993184dff2e4c572e2e2930086138735b620cd157c06fabc38d526e39ade850100fc471c2c1dfa342da8ba6e6bb61734b045661af5ee5ce70c15a77770cbad6b8069e3173d73cd43efdfcd4a43c3544eaf4bf8d99e0afaa3f7a716f10546f2c620c61d28b7ddff8cb04182a3659487d212bb6d8b2634a1471f07661e0035f65462dcca8e9d0b23e51befaf96c197fedbeea6d4d22b2d182c5ad5b37afab347c8e58343eb86f8963c7777547f8e8fd7c3894a9726f1a624e4bae53a6bfe5b7d6d2ade925d9fb0afd2f2ea6c2b46163738356a2c0a389ad765358e3f0083e4f9a6c09ba8f1edb4b04e902888608e9e2725ab422094526104bb8a8cc71517d167524200a21c23d2197e16bc7f8a649de551e6b6133007aaef637b3396f2e91a3f4a849940610a2d33be6c4b8430ab9b530a0e3bf9cde843d80f29299ae0ed3016a455a2593df6e0d14e003d4da0a399fa1636319982a13f91abc7b408627e3c51c5714b0760e6db66d943718ede1e5fd09755892d1d094120906fbf43620113abd2c1118a85f8aad3a325c972deb71f0fb1b22eb76c6071468503f54df376fb0d4c891d1d67d98efdecc6f98e1a9b677c2194737acb5225293da33f764ab8a8db50d0a25d76b8f14752ff17071a2295d2563b2e8d1fb06b4b0291e149a8d7d4bcc811cf354f928fcded2a65a9ce321644f5d8d7af29fb1032d6521cfba9731bc77095fd91bd6f8a1e113114dd4c0720dd01c097860bd2b9eb39d39cf2f5c2fc7b28768f7a12dc30d5dfdc9ee36d6ff03823ec8a84f0e74145e7df95dbd758c91990bb83453f2550315d15e3bf5bc5ebb50b94f4300db5496b100a5d976d0b76a22b37045636eb672bb347ac38baf7b0d2cbcdf1c04de96a5a4d5ed3c0fd02291dfb841277d04747b5cef3d513bfad17a64683fa82c413a7244c504ab2069cfb04966148411f050477476c00f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5cfadc11b676aa583392d287879720dfc6a71efa6143c7315aa798da4ca3dd89c81f20177c63e58de164b65b57595d6451e1fbedd832808b401a6182973de498d40dc892e0c0dc047bb36d14afdb934df7dc71eeca7434fa70c5f54a7e9c7a93ad4e8fde2a3b737853abd2247182131f327e3fdd7864c8c12f3f1293bcb054ec6ef9b65bc3dda5d1b7357a06cee4ce0056f9b3230ace89e054b14b483728eb240cd829f58e9dea2105fc4ad368e142d211352723122330254caf9c38e32d8967af542f26ac40ce772b58465dfddae45d39ca5897f091456a8ce2b62f0a781d940dfb6c39a3579687b634c19fff34d388ce569da08050500345306315cbeb2e8f7b6cffc51e4e7a7243ab7270026bf10bc564c58b68df50781c43176e000590c36b153a446d6d865c9a1b06ff8236e79861aa05e98a859d30f877aa20de56f5b5b0f305fc20b3b73f383b7dae4599b2930d5f271b2827d4df146f69b72da76e284a14ca108e7468f5c48302e484af65c9034a0b9b60ff59d6f80c71c2f4ee5573de9a2e0da3a0961e04a4ce3703fe85fb792ba17de25cb1777460f8261407486e12185b091e65ff0bc1a548de78bda5dde2090c72e033abbe4cd021a93a0a61bd8252269adba4ac4b78250d106b772a8f20359e9966baa843cdd6be1ca66d5281c4710b33b419f03302d62806e1e3b31f180fd74fff9a9b0ef0df353759c62505b47b9b053bc05637b7d6cb475d12f456956062f9eaf6ed9eecb3de28880068c2c205a2c449de26849413b867ea3e2c909d4969244dbe159861aa0da59d53f753a9026792d02d318a00f8b0f15f18e41daa7f5f03c010888f8dcb0c72810721157f8cc69da56dc312d11f3e9db6d82e66774996e6852073023394590b35a87a01c78bbda9afc3505a94096ba81d9c11aac3f9c8d9d64ef657925e72f8249c07e94cd389cdd9991b24dde49cbf3bb364334d0daeeaba3961c2d355a8cd700c0106e1ee52c4ac721ebe8efafb9b9f1dbc012864be84808bdb387d1258308e79b4fc5be451b413181d9b74170f3a850c62f8270c558af09c49dd5ea82c5e5515d77d1307f42efd9fbf908dd89a4c7dc94d9c0d477c01b50de263c959d31a00dd8db7f56813cde325d6972fa23911c23b0931b042a819d11681bc545d31476c0dee4b9f452f1c843bf1a4f7f71719c9e4b35faadcf883d20c584cbd1dede1657657ef4eb787a9b5322a9cb7aea5c7d0e6886beb0637537d6f613dff2508d2a62267e8f8a5eac743d9c080faa1dec6775fa90461b4465695356ebb793d67d711dd5992b1cb80200b70fbd37797625ecc86eb76ca82c03875b2c710ec79fc77d2c6f325452fb34094b53f959c2720f1e51857d55d423ffe8c6c5368dfd24647c61ca4c4c7787dccf2625b4302e252c9e40f31a94775595c1795129d842ea25aacfa7894;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfd79179335b887e539f4f3df403fbe9ca0ed9ce2e9feb98fd8851299bf6619ecc5acd23c429b6e41ed92ca283b0699f6a13dbf2a8f9937929eb2af4225b9f7ab7405265bab6d67a64ab4570a7b73ea7411b3cf72c769d97a15b398dd1d4fa40f77382d88ae75bead87667c32662e2397b285e01f860a0794e6918bc67698c6ebda5601c16ea165323e33b54b0a0e1c48973c4d183813cd1038a144e4e097f9372b0accb316d5b57574ab13ff2e6cd8af8bd5508718ae4d0e25bbc0904417d7a0a9fad6609cc9cfd0be6919756adc348cb964d99ee2fde1d3f3f6db21118389b7a14658330877c582bd2f1773d80ad30351a530d388d6272196fd978b4022b4ac647bd1d041b77ab866a8762ff7ff5794a0085536a798716cac072680640d5db604e7037a55554c47a5ea4676177f60ffbfcf5eb53a202fd0269169dc6f68f78a70733600cb94adc8bb199f2883db1e4a378f5cacb396ba1b9ea9595585c729e20e9a4dff4dc91311349d6d18022bcc0ac7506ab339828c8b4f000d3de2de15c1df0a6d2e880d8a7f14d47f0524df36c8e4af3d582646816e562f6b4da64eca20f49f57b600e193c86eee92c8a2179bee3b8c352ff16e188dd1d876eacd6139a5d3828d67c8a2280657a3104d840c15434de09032322a2586cae84a9464ca6496c335da93a157b2029b14727eb069963090fdd8fcac548f24fa48cc0fbc5d8f4944ddb602c58929697a99823fbdcd1408e208ae20428d59375eb3b45607df94c506e2c27e62b2214eb94d2f5d538e966ca620e36ded914892b9e8d7573c5a353322b77cdbccbc1e01dfeb6838b79e3ecd0843847efac373f7abc838a1d5b3ca41f6fcbc46bc3fc0439f6c76b8e26dd7c376dbda6132926d9074745e6a9163ce5e2f93ebee67b1ab32d24525d239f61b494c2c3e02b0b7c121d260a971344f8ee14b7009f9e679410136e50c43f41c3acbffa4b3d886ae21926b920fdaea2bf99d70d4a2635fa822a35149b72862fad01191769e9c23c863851d3136f228fbf3e4d792906422e1374d0134ce572b9769988edbfd382275e574a9073ea51dab735166245ecc3937f82ff13e19e0565197f8f16ec9e9199cd3abab95e70608834dbba019da2b44ce20238b2f084180301569cd97ada50c96303473ebe7d502bd0c2236667b4c30d52db9eaf5c637609cc6427959b0b77c11b246b9a2ddad188ba0aaa3c3173eea1da01e861156412f962413f3b9677bc98ac4cf165e3dca662485250b7292345811b4db9d4c5b11c523699520624bd41e36a070ea4843cf1d65d6510f67b8ac02657dc104f60c0b0570e3bde555ac0f11f20c3d7ffae9578e16373a86142d686b2ffb1f110f432060c79c566588909faf4dff873ab205c91720f3750546b628c1c698c91f581a53e3ab0bfd60953e978a046a8bf28a2b9529191508;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd21790a2cf49762f6353313307cf6da22f3ba06ec504db47fe708b36f4d7c291abba4e029af49f92fffe197a94c12cedeb40b2d25e5be22b0428e55a5bb4a292a6beb0ef69835e18a3d2cecb4dc73cf9ff392de7a023859527f1fafb25ad5d68e05dfb754590ec7459a8370d5e106216a4efe13e8daa8e120fd6ae2d3ade67869649d2b559c223ee83e7cf5343f46ac6196691c7b3c4f88d4233119092e0c734ccacfe6df68c3baf78a4020531a77cea42fa635f3fe1cffe8ce338d66bff1980b1dc49ac7d158948dbf59dd91fb98bd30b0c9c511a80c54ef1d649cd4c58d293cf90f478ecf8febd92892d9832046593239b5ebfe4e69056bd25f2062f79205ef1864c2352d7f9ab5b09cec312a388a9fbab70921794c941e25705522a8b7758bce15b8d479c226613092efde1efdb6afaa00f9b09addf2b341f25c9ed75a91ade48532ada8308939746b9f2b4a5336aea1fa5aae8fd4c37d1b5920f52e6ac5035594cdbbde9284f7ab9b5cf7cf36ffe551e2bb9cfaa3b85f70c4fceb3ed32ebdb34a54e625b9f2b76dd112e987f11c6348a65a6df691041e3cc986c1e9bbba547c90fef164a83c8449435012718b1d9c11e67057ec969383a12a6aee128efba71e998d1e1d02c5753fd9b20ff36c66f382fcd8fc4b9f89654a6723617e1c73f2ef448b506e9a74a9a8220cb274c9efefcd1351c76631f58eae2e0cc241b0b107df3181ac0603e2185bffe33d9f076238cf767cf0ae18c8d96dd155c1e5b15a71793425fb67ca857759fe42fd62668b427c8a1fb261234ccaff13041f91d4686221ac9e14ed5a49e9387b3ba03d5d4b79dca17e3ed50a67ca1fd1767d1f9861e0df7562aa0a184e30b23dfe2bf22e40f7e2cb3da2b48c90b52ecfdaa0f4aae4113f22c84f59a6a1a87bac16d0327e906e3f284be78d47d3634efe8003b093e82aa129eb8d3f580aba4769580c56b9d638c0641f9023609ab7b1dd7b7ef8b8a7ac440d8955af5a97641540b45477d094621f0a2ba787712e21159fb1dbeec1304dfc8546240da1a24772f49e58005985d8b30e2098cccbd511c4f6a8a6d85814dfabb3874c84d848fd7b300ca6044be974235e94518cd4e1f09ffc0e053c106a7298a0f4a1cec84122c008f18136aa4356007c99402b34aa0a47085bf9468f21a3d0ee191c7b0abc741076ee9f20ad697f446c25857262300a78d14a6bd983cd000fbe9d8027dbf39c87a70b6da3c0561384e5681e7460e8a2940f792296f868518e7fb481b40de7e6d1978a96b5d991b32884d118dcc92aa6b52becff13e4631dc7c168b7976a0d715d03ebce6b3dd8fb1dba0cec8af96351cbb3b155d8bb2c211add74b467e205ac7986b386da8fc72f12dd174d306c21850948577ddaf898735f6bfa5b2deeb84fc6edd80e5343be5a182ad441134767aa5a04c99a4448565;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he162cc712808e03d950631a2956a8f6f90d2ea6862219ab5bba2c496039902b088aaffe490d50716f4f181c443554a8e96063d01fd96ae1fb359782b7a29bd39c8073a906f9939c1734bb2ce5f71fdf54f6fc12c0587412b534f7d5451d2689d56936c9da859ae3a7580ff9e60463cacc84c0789bc7ac4655c6206ab819894746295eb65fb5a4e880dd37602f2773d4df684a3f16cdce163d5a45bd580ded765898382a58426995ff98c3d0ebc97c3db82148fa03ae6cb7b9161981d42d16ff245860f5e767740e55d7bb317a2d2211acdcf0e167400d0c6d3d31be0d32c55043d77739db79b5aa093ccca322e09347be7b43219fcb64bab7d157565901934299fdbae2523fb2f910b1bc23622a06d7f70fb23b4d7978c938275b7ba5d2a6d638e77decced85eed0219d0721990b5da1b82c34bff79320815802557243d6464ccc3cc5d32340b14173bae703b31cbf3472f61d83a1f04ca2e24b8cc68df31a3a8135cc21d4fd370dbdbeff6253c2a8fd0469c0dfa410bda7ffb8b1dc57cf5ae79a754aed1528d3bb7ab403924ec5f6d05ebf36af676fcb7a852cc4567499bf660af135d85f64182f16fa76fe5f53628e0b978ea80ed48a07382e83ba47bcb9d8c595e1abfd92c3512bf9c7382ded9f26226a0ad8cd8a44d3c12418dc91d557aeb0dc770a82348c2fd5cc6a9bcd8e6014a18798315e0ec43a40f03b33252b53158aceffd8f93fab0b006be1f68c7a770646eefb0e89019dd2a9b420ebbdb164a0fb521398e1b570f42d65c0487577640301a0eea065a7a9a516061bae56c1d610c8702613950eae09c37567da012199cc05a5320130b14050ad68cdd1f40a815a3c0e8cb02ce92aa7787d04b52e67100cad2c53999253b32612e4624ac495ba71d84948384ed1678e339ce57a1e019d3526cfc63c54d6b32deb73a9286573c8f50d1d55f6a457ca8cbcd89e283ad8d829adcd44c06bf6d53e03ab7d8375714371bf8cbb9c341053c1a68d1cb812d3edff973b20ae1c52a681926addb6d967bc85ce6ea3ae3745a7d728b4f99869c795f56ffc5c5e1dbb03e1a4b224c8ef3075ebbc341c0cea0efcd873725c9e8e2ebe86d4c37d647b615de04f21fbc0e991970d4c37ceceba8df6f8a022f4119d02ff1f797119c039068f75c5fb37a24b72023af89968d42731b2e5410882e6716556e87521cb6714394f9121217c81dc34e698ebaf98377199e422785ce116429fb3d649529f796d43bdef5682de291f64c9b8799b120ff3a3cd687362462fc3665f35857c42bcf309ea909649907b346ae197e69029b6acfbd5118298777b88f8772cfad49e901dcf9e610ea0ed3e9766d221c1904fa256ce639852433a37bf8e9612d55f674a658b33f565d6fc2605de2d9546703e31b4f251544a4df0837c4b5938dfc0e6202a314d2aca73f93cb9622926;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8d73c07dcaf2dd214e576e73ce8359cd73c8329ba6fa6b9703f49de312f3220df7af2a6cbf4a9356ad784251aad52edf5321021472498255c0c659a5b260270b5a9e9875425dff793970595f500e2ba54a3e55af3646ac49923e1a88707265c4bbcdf7a3634bbbb1ca9ce789d88632e2ef9d6168419f45dbef8d2b2d692b898dfde978c56edacf75fadcffd5398f0cd7d1643d7d3eae434d6a3359f5d7c82107a30cd4ff83c66ceb8836957e0b6e4d2ab1fb2a5ccfdb978e3078b6e30bd66d2282afffe51568e672ec3c9e39f1a6027ba24224e4f9e88b156ad0065ab2576b080301a78501e61b3e3ebe9fe6f49105295b132401255a0a11d91d9f313d3cd55472e072b2b61930337438adb1a9712a01217dad55e2874375f6e8cbd8cb31f1c978039bf84d65de2e8baa62d01e59458ddfec82a618965b3a60ca5e2ca23203455d40a6c5c4510845f0766ee0d9b6119dfec478a656c5a1465bb94a4a5d729d7dd16e218010eef4ac398ac44557b7f21deeaea0e870f294f505fae4f3327914d43d054f6703587915e2421f20cbff79465cfd7c731e217f0b724e681d2b60ebf5eac29bd50e7c41443c04d91bcfb1f0b216311e70da5bed6c6d97f109270db80298d76ea2ed3c771a9921ada3c8ef80d59cadee98efe849a0426708729d1c51f6df2acf2d80b1db5fb5347c8a275f34899db06fdf4bf213af120ef05c90c06f6ae00f0076d60f8ce3914cad1d82df427ed992f8b0e9e10ec0ec69d22f89b068bad2cf14da51db4abd6ad91958b0963e08cecc5210f28bd793c652a160dfdb1416c3a83df1e00211764641ebea998ed3906129098e76af6a5e8cebb5c020ac6631097aa9451709c518e5662a7dae481d6efd81337f59f7ed5639ab17c875210ece219fbd68e6c6994b43e84ed56cb7fdd71e7a534c41eca9cad0f58904cfae41bfa8d1c3aeeae87635094d325ffa11b38c15e55d1802bd073b24b4751b0d33d028a4391f6682471d6c70ca68a8590df0ef0d2591b72ac6d8b2eb4f8693c538f64779abb6186b7c4e5068594206325b06789a2fbd42c1a23a77adf8d54d110926c1dab797631646298a95cb600d3a01ad158e9cbb996f9aba2de8e8f7df229d49ba961c8b873c6b253a3544b6653ea228339b5898d51db1b1ee3121495124c2a6e9c3cc4de29373cd165135c3f951e5ba98b300e3752755aae1b924e887f7819a1c805739164e535627caad18d39a2b745ee1ab4a5e26725615887c3416c6caf87dbe0407388b0f84b21225a5392e5ebd22c090cbd01e24a21823295db5b15900a25ed0442c10132521ceff1223d5cc764a0926508c78d40e4af52fef52170fecbf3e505eae2f4c8475433fa60f038e2657ffcab2732469e2cbee6bc12dee4ad80dae56f8dbb0ebaab9b1d7ab5684e6304566359e4bd633fbe686dc42e4bb4f4745;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2bba645f34a62e644069cebdf1b8a381b91bedb05b548a7c737a8f1f39b2e9c3d479d3b4241f82f4495ba7a732e710b34ae4749ad7ebd3664755ff99f2d9b4e4c083f42402d6c1e05e710482b7d2604cc14a16620f2f15ede7811227ee14c60bf9011abab52224321b369de379915b905ac26f177915e4ce0951fda3f141f36008145a67dc1467d3091e85b4b0b5ae6f7f5091cf40b4f36e2fc665cde38ec03e0d1ad9675d48dba7eadf033089cd14454f6362e268899dbf92c62ca2aca7d7366a1b4f8a2eb5562e15f02f53f3b6ec96d72a47cf19e0fe8075e3c3d120e3cbfa15fc6a73891059b2eba713dd9dfd9803b52e042a4694c53bdde060d3c72e9610e64057e5ef0bc15bd733c1649bf3536a1ea0927b7efae34a16a5d78b9ed857b648d196c9c8d4c72cd3454f4b65733da818c1a8117b22630e5feeffcaea747e2ac88c73bd6e807839aad25c4a8b933a8a0077e0150ff5c16eeaa5aa48780dad44379ae7f12a28785cbaaf8a651e02b10a7e86d27f42127309fc2dc4ed99b02226426189ee0ca62db293241a36151f7f1f98f07d900c9d080a43bde75d15e5c2925a970f4856c70ed19da1b274fa2e0297e8eb81eb97b752a48acc71f0d4263718ba7781d3b973656ee77d481437489e2a37b3826ef4207f721da9a41fc0cdfafcdeb970ff6dd98b6cb2e606f05741a46930f4f7616d8fede70d0a134089fdebed18bb556caf68d6be1291726e64e6be0691a8955eb84bc96b748be5cd7326bf7992c8d387d7a822c4d84e0f0cde947d691319dc510d1befa559b4a633078942b8dcbbfbc3d1ff74d5bc87eb75f7ccdafbbb3c14b388dc06cc68395920b590f604b4749daf42c4f381ecdd143b325c76ae047de996b00deb576fb2e7077e630283db7aea9418d569a5fe420cdd58de6923f6ced2d586bb5101e08a25cad8d6f8939d59159c6ad1d1419372c57035a60cf5016de29c5519ad6d6bdf8feb9b7d1cd5612f5ab383909c0df8cc9444ae35ee9a10e4dc67fd64b46a5e1596f6a78e9a986b6b1ca08ffe2364209c37b6b536464b8227327f8b4a784504a8892c9365f19047bbcecd1fd3babfef6c92a2d8c6a2afc2aeb77cf9ee169d1c43b0e30ee876f0db0aba7828a5b753f0473642efc59a04828c3acc89aa4b495caa151043b8d8864faee324bea067fa805e5b4a834c64af332ea0f6dfc93951859a612ca98e035c50db8f0e65068f1b40ec89fd0d9c1e46f4cd21084ff6cb259cd9e01472a747b9b6f1158b62613304342ef014d5e5327af320e7dff437201e66431a7a7f4ffb1d04421b4b39f90e973d50ba61c9dee73805b428f650ce67c107a0903976d02c727f30c02b2e93ba66f3687a3681078ef7725ba89e38e7916e6bc17a8b86a44ca01fc1514b6085a6bdd44ee69371ff19b543e3df47675a12d1f998eb4160aa6307;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha59947b3f21e47255d37e9c320645261deaa1b3bcbda9ebf483f2010f0c41706fb4f7231df5b55cc0ceb77afdf8a39209cd5b6b52a9e6223add6eda69e58cc6febe53f3dc7dff71a7d46f7b65121484f2c43b008bbd3c1c042d755773a862b9704a4eea51e5a84b43d20f718646fccb1f653bfccd177bd285138bc7a201a3d3cc60c8d7895a12e7077ea5768fc5cd87b0df38c285decf5869ba80aff12662d0fbb7478b6d631cd4b82b8956930e7fc6026da1acece0d336cd428a6ba041492c203e9ef5735d692dd2a239435ca94141817bd6510add44ac6bdeed51ed4f96c6eacd113492a526035cedc84cd2d979d9a1d2910b175102cfdf9b30848736aa13a5b8701c21fcfc2539165bf4f7f351b8cc77d79bd42e1181a24fd360fd49256cf4730b79a5fd9001cd6dfd4b5e9d2b70a6861e86389c6781d9f53a4c972c59b2d444737ebcebc39936837ceb460d7d8d2d0171082cedeafd975e503957225211a43928ba7d85a20c9fa8efe527abb6b772874cf494f061e1206b8c216999aa945d7c5a272989dca47a7ef1db031d40bc964ee8362bd445adb97a4aa67c4fee9be8925e41a94469ea1caa438b302663a4eaa0ad0f01184e9d1f51e973a8d231532fee24248e6b036edfb79a6aea54f4b5c5ecbf51bc5a1a114a7cd0492ec4b864747c33e2ebcfbc3d10d6017ee663282a7ef30bb262df9c06c8276100262f4ae10223e10e825be936d8e27c6a6f4c10b62273a76248c6828f91240461f24ec72a5cb577f9f63626c41b34c1452e3820c731648cc35079d9177f038137ff81d2778633328667616725cc69c5ec8eef38d38c5d3c499e89020581f628205fd840be484f58f2d98e61c4333617cd12ae6e429b64ccacd0f026163677ce95fcb469eaba5f7949f82098e4f5f4256af93e62baac1d10b4263c4fad9750df03ed062048255b9ad081ef03f0e0f679d3f83ccf6d0f2eca47732a3f8a6708a62235f974e69eff9b76592d0c32029196231b1b8defdb91d34a8c239b3de712a56fe166e0c31c21b370a5329a75fb258ca66e894c68f5badcae8a711e5fb4fac0f7b8a72ae7e22a18c9aeb6203d179fe7e00f9439acfbc072f352cc0fae0ee7261dd8d3cd420ac8e95c5ea46c54c52001d7babd52f292d132cc2c5927b8488dbe5eb088d3f90b4a5415e516008c65c33de9672504a0059d7c016651031263ffc406cc171cc9c5436db0f3a9e972d2b43cebc8edcce18334c17cc27060dd2b92423407731984d5182c3dea6cfd2957ad23649c6b99b5987091834d5c0d55c9f57df0d427124bf94f283f2dda4a8ceea0ae3c04d54565a304f0396d178a3f84437a70ce6b6136fc0f82974a86ad5b20824db312dee0e8beb024de8025fab1f92775fa86cc245d2864aec5042edb46978404408bbf7fb3f183e4aaa46263851007523eaba5a38bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3118e8437b3381ae2221d3bbe5260ee7738e1e187a057bf0d110402db9c732bd6b2dd1b6e12589fa1d66a4d2bfc2c607e36f4afc019f8f5bb6706ff34eff068a91cce64fbe1cf8e61d3930767443ce8ac85d5a8145405075b2d8fac00464f9df059967e260ff3445a25d7dcd763610ee978af10273a198be631e3e3aaaea6da568852ad55645c42bb047867c877e892aed7412108e9c6001decc60e4253238e3e8a791007fb0a917b83bcdf26728bd70e64b8b4d89240c5ff4902758205f42ce7080b8a8466967bcadc9aafb635a936b32a816047673f6e71b970410c3f4aa5b5379c70e425654d30a27b449b9c65cf2f969a179f3a55833e671bf3b4221af7066923b9ff64ca4e53c40781c46800f30e36b843ffe96013362feca5723bdafc4c888d6f304c215374b4585cf3f16053592cb79e9d1db49e7a17d20c76101397adadc79742b7cb1067a70f667e702ba8937e031737bf4be13fc77741c311e2203d00821281c8fef9ad32ff37b52be5eb0104922c0d328874ca8cb639b516e8efa306403b81e27cea6724aa4aa4cfd0ce037ccf71cdbeb37df9fe660642d0541d9202b32bef563144a6489407f90958bebb7ab4f48f120ec2d024c89b2255a02271ee70e228063a03ef1fa3fb7db75412efdfbdcdf8b065775c6cb63808d1606b1dedc337f6af95cff8978f1dfe4a8828d57f18976a3ba30d12a998ea66828d5548ee1e0f472db53ba39c5f1401593a70da634a731804ab973c112202fb8d6e07ac353db7d0826dc6a30201200460fbd1dc0b996ede7256d6d0aeec146066f457f77e865506faefa651e881f1c40d5cf0cbcc4b96210f8af05932ce8e0da6a79488dcd6cf243ceb790425152b84e07916fa8b77d1c09e8272ec4d213f744b984bf13cdec18a7686964ee332f0c80613246a589f6e86492b833305d7069e312117b54e473def7d12003647758448ecd034ebb86dac0fb5616ffd37fccfbbb079067808fe34f3183875d4a55a0eaf509d03a79b5370bb6f04391b9cd2da1f819351499ea06a3175bea55bf8549fbaa9faa08ea5a1eb5ee90de3bc8c45d2be20d7164998b299a8936e9c018bcbd7fe46587a1ca38c88b48bd1946d2fe124ca6a03c06b0e2b106f7a74e31a548fa6ff8e913a9bbabb912b8f33485486fd291739c1dd858eb46f0f5a43ac528d6969d3808ff0895698d915b165e1600bc2ed7ce32f294fb905ada22f09cc13228e1847442ab8327b2627afa682122a66d7d79aed1fd9ad30b688b63de7403e45c663dd5d4cba80603f69c67744553936e84c42dcc7e689e9792eccd76d7f331a53cf8c2d02ef77c46951b6263c5b00443dfc129c997e2015aa8b1a19b4f5c5ca8afa3a6464aa4cd552cf25edda7d0af87cd88a0ffd86186252eb2e663b50eb51b92f52ecf30068639f83af5d3e528ba4fd5d5c1100fe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7ca536ba49cf1bd4ad1f8dda0cdd60f770269013a5f479d0638ad2c9a96f0d14f2de6099b2e874a22e3d86557c315e7964a2db25431f84f2bf69b7b595b1e683e3f29a2eba7526d4ffd587e22260ed8bf7c3cb9516d7eb3fd26a8418ea5806a1da3c115e3da3fb18b9d0821180d3ee034ca9bbd99ade11169e2927d26833a88f6d17341fd7b94d6b05aff57c99f14174b72709916e26abd729e716b18fa56feca4f873753c38bd33b8416292ce3c7043fb44b46f8590d772256437c7a3b38aa96f5dd9b9be76cfce0cfd3764439dbbd247631b017629e0005f38c235e7c4fd7f6a558009c39af287fbe93b80060b14df8e330091bc22352d2c861d22262d5de79f469ec86e15a554c8c095a8a0d0a438aebfefd29696c904b4bfc0fe1cece6e9de23a0caefac5656524952ecaa3f5018869a4df055247b32fd05e86ea85d4d99034b2d1533ad8e07f57ae049015643d478acab322cac9f5fcabee7ab5f474ee1ee54c7da917442f31932115b3537939e528c4c5f1ca2d0b6c089fcb5329fb1496cfa151e0d8e376680a6f1109a8ac25427227294cfcf68e32e6198530e35ff4369e5f396f03145e24c89086f60b17f997d8312f0a89108d970f87d46ec559047aabb1356d6cea26982b33d94bb6c708d59e6d9450c0e7fc2d6ed8456910df1384ed876975ad2920508c315526796371da954d639e5d2b4bceefd0b720ebff00cd8e79c73a709fb2eaa449c3066ca3e2d0b5cbfb2118820a8879b1ab909ef8a7baa93b8ab1d5671c32986f2fb197269e660a884db6536c7af552cc404c0744d9766780cedfc3591cf746b69fe8ce8899f4a091438d1d5a3f6d045efd3a73d3e76a6ac936d53027aa5e329fa3f3857ee9095b9bb107b7b3c1832d897aadca5b411cabe61e02c25d72ec530bb8a17a257aafec05a0b8704608b4d820da96cec314c0ef7b537a14ae2b8a2cd818eb8cbc988290f02383f661ffabf5bbcae20f95123d4d1588135784a775e7007be6a2c3aee1f002f6cfc19761eac860da7cbf2225c30f7b72e4fc482d0cc201640696e9843d6cf9244fb517d667f34746bc26d4ee6431b2ddd005d1c522d6c57a9ffe3bc1afc13f20a7037504e5f024039dfe79d26dfb9c673516b44d6d5e3408d5bb74644887294190c40ac59e7bab9438de40c8e0785ece08fc8fc71777aa7a12ccdb507380e16ac105e76b404827344554c47e028174fddde900dd11530696c3bc157d39a0ae0405b373a3251a3c94d2885e78644f145f982269cdbf9a97d67baaed2320833f8b78af0d0bd789add5e4b884d478fd0bcb3c5c19ddc8d9471e5beba2654005e3e71a76f943db32df9aea0be81d84d6463dc4f4f1903463146e6d6e458bf0303e3222a20e4be6a78a7a7268d1b8dfd48d49aabb76b3838b81c6c7aa08805a72c75cc9593d32669ad3695b72c68c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ba081ef6d1f660d61f8711dfe111ffeec14d525470cd573ef8027c324d9734ccfc8576f439e0347617e6a6131b745118a0f909bc0ba7ee18950594ee74224dcb0108d6b0852bf35c519de78d1e5e783a6cf293720e0ace3ee057030161d3f5bd6e6f03d5550d95e694ba61ddf1ea62d4296bcf0ec1d116c5850a0655739c0b5ff912d54ab73945c7e6ec2bbf191742882b0d895e592a69c14bd79522635cecd758fda5a9c64c663f56f7950521415ddbb13fca93cfd42765feeab1c66a06c7125f81cf924743418dd231ddc2b625df5fb6472de787ac1e11c0a839517daaf1fe2348193d4e7a6ef23dc82ae5e3a55c660781f96a26f0115392f39a6a6e608a77073620f1ad48495ca779a9c76f08e4a1ef474417a6ea3333934767e6c8976d619e13814d3e5a116a5db046549b97adc7b261b7948fb64513dd1428deb69a68cf85e747f7ec0df7ceb3266ff0d1e3e71c3927eba87a8b771d0a7d62ff4145ad6d53a04740c2d3504b0e1d9e18d15c9168a2dc173114b42a3ab0ff4901cc577b025601f0d66838b38348752f38eff303bd200234dab22b698372d19967d4dbd28c8488bfbe4c8dcda10cb2fe568b17cd81cc85568515586de3aa661a93f04c969586f2f395ec753331d37ddc975d8af3048bffc5e247f136a7e22285b389f995facfacb9508bc6915cdae4d1caad2984104d2d5cfad4f17aac70178a3cc164b613dc1b0f1b22b0fe8d176b675500ecc8ca4cc1cd022d23a88ff571ca0ff229264805dd0ff5644e7c9aab54583a059c22685536f2e2a3cec9c675557535dbb921dae831653f9e53d72aaa888f2caeae1e6bf60d0dd39103ce24b3ccd58530ee28af2a298d4632e0a5cd2ffa282d10114e9f31e6c3c6dc1df717e30649392de548a42d54813d383e2aecfca8c2d1badeec4d7a210f093d20697ec209d5db19abbf0da94d9c49059b4cd6e25cdb1c21806b0a1ac00e7b038a41d7c4af48a98e875472a811a1bea28a0b8bbdbd16e1b6c02409d1f5ce5c582946b30b371b94007367580b69ecc6348e6da72e31a1a87c14281fdc956abd5865413e22e095ef283730c473e6fafd1a445a82bf88ec58a80e0e2f3fa8182d7c183b1aa754de3538a88ce1dff02829417490d3dfcacf5489cb328cc7600cb3a4c3635dde17d85a730784573217f72aea30754737e265fda8428674d59547fa06ea98c8ba546e5fb80277e13c31fe339cb50dfe14dbdca66d088f23129e481981bded32a5e00bd4ec2c9a30fbed553a23bca64fcb945eac47c055aee9a7c9e2f6582f2bbc6d03219f1af0e8061b227dabb37046fde57a2f72c204fca76fe39e60eec465b094c87ea6116e928fed02e71643270dbe061c02540c7ddc5406354194e1e9f60d2b5d1206c1e746fb86835aef07b23495d8d202d3d208e21b94191c1e91ce0a0fbf99bb5d50a8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf90e6b57fe7245d48fcbe979b70bd7ddde3f17ee35068059e59c42715c2739408236a32ecb8785fb00fe8c37b12b51bbee81cb8398f4d28259668efc5e0e61500af9644f5634e8c75fa0361256bd22d5fd75827b0e0d3631873b9bbb499061aaf59eb92331da82c98ebfe0b71dcae4636e9bc31f905b9c73cedef34e51509b06c6331a167de2b15b466617f35b91b57b792ea4d49c42c9acc9ae6cc8dc4695c3c8fc1d2d2312a19962e6cd22b6614c05101d802468e016748cafd66aef56f12ef9d0f63b614ecbb774b5ff8bfdec9380af9985ebfe5a510cf1b43d7db47af7a329dfe35be84875d0258796bea9eeb608ef61bd2ecdd76eacc0a2630d65f7a1682cf1c3ee7a8b0c5d3be5f51e9aeafde54b5fcf0c82631596fd1332da7071d5f9202909a9c44a694bfeb423bff18982cd938aeecd4c7d2891c55c1075e82aba913d404312ed8cb1083fcaca51d87ceb670883b90f29e4662384778c85978e699f4ccf29a9769740859a6c80478bc328881210f5125adac1bf555236cf63364a558e57282b75d002d99333f734e69a14a8831d246c772364efa46cc0b447f426228103f1943fe7094653be75129042867750fa6e77e2a1eabb18a2331da830ab056170cfc68c25856a6aae2df818afa40f66a2d55574b2cc0b68ee6ba9cd426de90805ac9ae106898795d379ffec855898a2c2cfd7502cd170911f7325e6c7469258d85d69533946c2e215a08dfa70230bfc736ba4145c89186cb68fbd4c9c60dbcb078b5d2f6dfa6c18ef7256c6399b745250e8b74f65adb300ff103bb872149e519b03f5583d4801e7ebb5523086418bc850911f5e4680a22dc103cd958ad3af4491f3cd13a7a719095a346a82ea24cfd492a60f35284a3a37f08e4862d8a8696c83017681435f45868160185ce70ab52ad1fbde052fae74de56a8e8ca26f44c5d6ef245d88ee44c3f048c2b29c5338b335cddc23a837884cb8dd7b4645ef242b4f0f878e24946c0baf7e0d0fbabc153b6529d6c489897369d75a834aae4fbbd36401628f4642c8b7334e997cf6fd60f088c545067d6d987de751447b58eed344482168e89182a968a638e087eb947d98e9dfafe40b565895d617429734f86111e147c8beef8f39a646f728285a337ac77458abdea9df442c14e8de4b2d7486098af62f1cf1c6549606b115ecd01e34d236b2f18f1319b6ea21f87712da5f9c22f5c6be52fbf72723f7278aace9ee912e4399ad112e7015a463c26e811a512019162c99be291316092d4d5d7324a2ad5da825bbe8e1869272e4caf43cc456c772bdbea5d68b7d6c59fb2e95a080f5b5b5d2a972228628f8beda95b3d2487905c4e149b9d691968c12d2d0cc8973c09b80ffad68346ee77f03d6fb6be523cd219b66d873d8b9cb3574b7a2cd991037383c99d80de4c7e722c475eb9d9cd1f1fc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3ed103a9e2596ecbbfadf48b424cad24f0d6028f4d6b0dae35e8d8d1a917d2d0629fd71cf8a358106c4414056d1667a58980f4008000d6b8529db1f6f1776ce43c520d0c65c81149993a2e7bb6bf6f8e64d4d62783e8489be6571f3da7e5de265936fff333df5bab8cd12a0a911055cbb860db872b3abca8e61c958bf00dfdf679265642ee5d9202208143712f3691a5a93eb01cc85f5972f26156dcc5834df13e9866348875a0aee9395440a0009381bf1cbbe963c4887c3d51f1b16747d026a960c9e215e26a4d7c9fb75f8593444cb1036c920cba7acfe52360dbb58ff550d586df88977075ee3e1c2c3c8b3b955b7321d5d5747e75512b7237ddb60fb6e65b04706267a57ef3985fc8765a6e7cbac343faa385b2cd3b7bb9e23883775cd1d7480745bd186018b19b267f86aebf9ef139b60b14df641d5a34133a6f9428adabaaa4753f56ee84b07b4cc5b1c0b093be564625b2fa98deb4efb5b6e51a753a5c5f63a8e2169f803a981a0f971272ea69ac2a0315598c0658593aca394570c5962f3ef66c257868bfff9aa0ac00161afaf5985dffe31e14d7180a8647e6827435d9c126684a17bb9a3585ed8ed5243b4f0a94f6861ff2d9ced6b39d49d5a9f28ecfda73d891e6c9d093138bd429ca472e35baa968f9da203be01f00f2460e2d843bfece04fa64e76b86634ec99701b3b368325de2c9ac0945f27500f8ffbb898dadcb31921d95eb1da47cf31f6de2fdb95b2de4f387b9eb87b8963c25c9f286ac35a2df07a0ac3d5e9d5f197601a2bee038f5fd4a76f4a6bb53e9a7cc19b91378bb4ef980d4f6ca22fbdeb669d62cd2fd74956a0da5eed0f5853a4b572712f9760f2cc31eda6a9457b83c8214db9dfff1e181a875862e513523f6445da86f12ec6269e5e20dd69f01a01c915c4b534bf59bb66631b3032be2258257b6adb468eaaf2fb0b95f0ce1ab4e5d800d9d76ba2ad28328de741a63635b9bb1bf15a7ae8021a51be1eec2bda85a6d3720ab8b6f4112332a8e79ed6b73d3430af9a636c36c4e6b45e59ceffa255b0168adb579e468257b2b7f2614986a7f243158dedc8aeb3f4efb953b7f0e4b0ed73be9028c703dac48daf7313c11eb5aed8b71b86d8dbb29f273d0ebf0b4f7836f176a51f4bbeba3cba81ff381fd3c96fd578afa0972ab749aa3e3368b297a389d1d4e9c56c27dbf5302b56b7981112ab1395fd272157a000c752fdc629739da9f041ff9280d8617d52f790a7df917f6f9486cc4d0552051649e5a8b7dd1ddebf6b8aea43b78b907dad558b8535390b14d8a4a5daeec4173c2ea21fa403fdfee0416d2a09e20335625c418a79e815c2cc6370c1779313610f9c77be62adb1655f6d82b538af0f90aea08153dfd01475dcc7619090061c364c4e5751c8321ac7c4bb82d4d23baf9e985dc8ddb159e833e9134e9e17782;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf1ba4444d8947c2a10c389800fff8a6ed7847f6430245de30c4c34cd69d34fea25bb1e390a9d245bdafdc8fed4f7cee56412661143f92587caaa507e8cfcc375125c7981e9d87d8ed89f246744d3795e8eb778ebd7025269b1297e5fa05decbfc064464cb812213f77e52fac68f742eb27d0ba01416090d5875ef3162adef086f17261c59b033cd84f389c574e4026f5f373c0f1316afa9648a46cff120b7b35ac47979cdb58218885b25005381fc6b198a5ca9608849433a04b797af4d5119faf9104d192b9adb06894a2c4d2e6b518fdd977b01a820ba0bb807f06670071c8f296906601b57191ef178546ee068bc9909683689f54304eec8af6d4990b860e4a86898ec79a5f49197d953836611e50cb0f0c4b1d4e92c9c3086e4fbc697e0d335fb7b412cb1310d307efbebceb5aaa10d9126e8482107e13bcbf8a5b5072643ac086ae6c69cce858b72bab27872b26ccd112233b6622c0f9dea54f21bb97ed881ff2d956cdf746c77d159d6bff86ff90d90c3c4da644d9baa213004dc4b52f521fdc17867919448c7d736375c7dfa733e4607ad794598907216c2d6d55d6d0a78adb270140363353ef5a2db4ac4ef3423a538dbe8f883d848e3ae342fe2eee30291b9e5cccaaf9bda1713c0591ef85492efd912d6c1874b3550e7dfda96d998bdb2f3e6c5c76bb1b35791248c4e95497b56f61f10b8c89431604e1e42c33cb5c8f55c0d182a77c9bb5c457e0a2aab4c990539a10b560a59fb35ca4bac25854a93250ebcad1409a4060e5e05e043ed7867d1fe7611484d3aa4cc15daba016044f839728ba014c2e09bded6df04039bc346e4214543ffb0f0a760966d4e23a701af0878f5e6fde9a4f202c35cff3aaa502d9cebc6a69793daae63477d39cb8fa5c3222370eadb7b8743787ec33c6597d6dc646671a26b5f6c1c35a14934656a2ba945a44c316cb91810c2321d4efc7f9feafc5632fcd6ad789feb290193be935116f8c4604802d42de038c19a1afb9b6fe5732255f636fdbd8835caa80e7d30d8fe705faa2e1a22899d9bddd93dfefee966a55c88c53618d02ee71f39c75f9abde3ab6c8839fc38d1e7c7c776f9943e6764d197fe012f296186998cad25117d46a4bcaf1e96a468074287189b450a2a3794d7854b95f6085fe6f5134e7a53f852405d548a1ae1735624104acd496c22b5cbf31b40c89c8e7ee27942007e873f24bde6aa468d60d1829f39b12b4d82e45b261b8884d8292093e1febecdd3e88bff891de03909068a8d83a1f3fcbf253027e4a6c32da1d540823327e4c9ab9f8ce276d04731d231cbf04da1bdf48484d8e18d99ee40a31d9e5f2e10d1884cf17057a77fc0994c2b4a2cea757fe5a2cc07a47e73c04fe0c452959c33d9cdf12365e31cba5d49612f0cc047083dc0cdaa96c6d4e2f7d9f3f2d71ebb33338f11e96e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbad7b2c1d05828aa97a0f4d22411006a98a930c9453d889030caaabca3a554e7651c10ee5e7170cbc7579ef9830271e5583936eff8ae3cdea56fd67ecd7468973d9b1dee9cee76c3e2a279c4651c7f034e46a1fdde75f946c6bca8f58dfa819d2b5181544e31339c740b1ccb6de482f78eed98f81a36cb8c673f7b87aeb63f9da8130441cf953c2ff4fcced7292b267413e506162e9197175bff16c20fbdf85adb01b7245cf8dad11922f4db979be359ba6d2bf8404fa9ab816bc44ceb92cc23a66b64485f8fb67d4c584573c9fb1324269b53c837a65b25099e353b993e13c226c6f3657332a067f3aed79fdd507250d23719321d6910b6739b202c2c9d2e90111182f2d8d4e690cc640ccdc3dd01ca03eaef7d7aae9df90fae4ff754eda888464113892ed62e380cd3c9d711fe00818138480cdd2daa228bfea216ded992f1c4e2075f2e472c5f0a6e71e367c4ec1b0732dd374137e0ef31b2db2dfd85c910aa621a6486d3078ada66e95bea038861c755bdb93af95a06e73442784c8f92719c4e57d67fcf77b8457a004d319217fd25433b871093d3b7d6a7f77022c8998cbe500ca4551ba208ff7c2efb0210d33f29fe5c7f1db5e60f5c7464b6791c5ece3e0d983fbb95770ae5bf986dcd23b9f106123ba092df434f48ce342bd20eebe14abedadf355a5b3fa4e7c3d73a937929499bbeb50e1b4a2a86507808a32abfe9944da89ed7ee7122f469775ccc10ba40a795279b3857de2d59c48a4f327de9b980a2612570f003156cfb36f963df55ff3b345ae1b4f0fab3981ea4a6df41b14a2635aad03bed0a3ae62db719935998989082566030cb0060c753fb57fdf8c7ea929f6cff771502becb6ef180ba96f1fb1cb2331609323de8957f7a8cda964383ae5192ec642ab0c905246df465d45371c5f7ea1b90cd07e2bac843098d1576267eef24aaf05ec66f2ef433d0e16f51afc692133b996ebbc8fef4d2b9618796f48ac56b937ba449a0906ba5d02f75f2964683e6c6575f1ece5b5489afd7450de88f2b9074482e59efb40f7b035f4cfa13a39588accc64a0cf5f3876b8a96374944449eba4a25a1da19c7bbb44f24cbde7b539992538634c58476763db3ff77e993060854a390d0c2f30b135d4fbf3ef7d9f7d35af1b7489c4677ddf20b45aa1719d0922e07d1bfbfb7c5f5ff2169824249b7af576b228503b364f5154b58198f07f56758a5e15a5ca2db83afc2bec5a7436421c7f502c6e030813ce863aa54a9dbf70c44d18d4b445f01943e063dae7846ea57af59ede08acb4af1fc6ad0ac68dbc6dd9a74b8f8e14e6fc46dcc1f3598289e3fc7bb5f737e8d6c24738a9a38016eadc07249fb909708385ff6d90defe1abcec7dd18e8e57afc6abee5f432aae28e174fe125de73724b2c8166755b4d9e0c9ed2a8639cb0dc98e195bd2184bd88f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb887f1796688bd6b95395cadb3bbfa7965eeaa96ef4bc7697efb6e26d7602f559afa583003da413c1b83f9323831dba2d0504984652add1ccec9030d48160bf0feb54935fd7e4dc17d0d215bc964f061a1da115f60f46512c5cc726e3a1fc3b8a20f7a684e7554c6958fbb658a49f8fba9f6d9307a57aea511e1cb7c8a981f60fd982adafa59461f3f9efc09c0d6f4b3ba3a7b016ae430d724d7f983e90316fe9451fbf6d342bdb7a156b8ed57d86235ca5ddde57886c888df0f0bae1ab70e4292493b5ed6eb309890ed250350d6b1d370eb746663d582cb67d6b0259fd896ebd3eafd022f00676b9f79a96dc1e924a7794a051a0dd0f75a38c48006faa8bb35b711a99a0ce1094ba972b41f7d87b79e796207c3048d0a0448fb918b4a9ed62976354c682cbf1645b9e59728cf75e3620d553b049199cebb27423fa71f8593ab3215529823c0b0e664fca19f3a4bb5bb9c002b28946c6e2160f92358fa04e792cc4d05000595a4e5fed53c4d1f468dcba1c4bd2caf4920a485ca59739c6110163e3e1da8442aac1b740b6691deb7651f640917ab592e0806261b28203dcf5baffcedbdfd4284b66220516ed0491e3b604d358e83afe9bb01b1799d42c9f5a89b1e5f817b3e9731757ccb6f57dbf07ce59a2b2890117e9de11cb08811de5f640efe1d81d414a1d524521e6099cac493320e9055224afe5247bd1b3d5d00be455f67f5182a53757189354690a018a14b2c3bd0621d56a79fd5c042fad26de841e63018238c63c6200a27e29b5f4577f03a64d0f320c52eed885ee68a3a9586c9dd821ea1c3deb3f832269240b170b61e18505ed3d36b0fc1669dd69094562bc36b718107c5f076ceac6dc0d9cc8f1fa524c0cf428dcecedfa703869745b68435dd7be70e7598f04984b8f2f16182c64565bab5c998bdbd95b5656dc176d04b878e6bec1e56a3ee1e670b3a0fe134d610eef921b283e396d52208d20d03e9e6721a29575534cc7f1b1e742ac3239395aca68f5c83d84a60b6493f9a917ba42c558244e3d07c33aa99d2388f30f2935f3c2148d792e0f6e0c3f8a79705207ee27fa0fabe7cc4a0f22db1c0ddceacdf427f9d001f97661eb10689a0388266003a27af71e464bef33bc6f349a4b4ccc86b4ec4edea459639e7905b9d1b64ac4e0f0cee820656e4be2c4c849f01cbdd5873dc239be49dd402ecd35c7ce41cf4fc268d094c3afa4a733fdf42b8bd7529341d539a8af233f242fead22d6255f40c28bdb5df58ceb5c91c0e82bdadca62e49e74e614c682097b18fca7ea6c05fa1bb27ac06e88cf690834916561634166184fcf46e9328ea9376b6a8b9536846909c4e0dae6a71cefced70884f7e99bada7c38f0595fc68b7ece5cfba30bea08d27f3379686c301c1f29aaa09a6c7e300b5695c82f9f478371ea555d5034ffa10cdc3915db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4fabad704222f81c3069d65b37884ebb352b40e02b0394d0d1ca6a61ed8942e47888086ca8563280db7a2012e0ef4294fd5d1b1c9e6566f8ba46e9691acbb6ef4b91d3d0e47ee19818c64ae132a5075e2f9b84033bdc55d19db603559aba91845b01ffc5f9bc233a28753cf45c044bdd06c91cf6ed9367366ef22260ab0bad1d0287860c2e3c94084d12476464f3942092b2125db028d54e0735b0e49d0b4fa81e286af10a4a32bdcb34c35e8b6483ea9e1de44545451dc9609681dbf8e35a3b802768c3f92d075ab540676ac5faccedbe8cbdd68f2d00a314fe73d64475e27542529e73e9539a20ecabcf5f8129bcfbec709524366ec062411f194806f56dbb15e7fc9e139ff7e3a2e16a7489d4e40a999a587d0eee9f609e16a04b84fa0a6a05f8a543011c64b9c47ebb783851b9abd3b354731528a6a53172c039b98e1e6c1b823bb34917da980466226a222997260a26dc02cf0b58726f761ad64c73480bb147c68b57156dd07dbf30dc2e86efa6ac4b3d1390c6415206eff82c20cc42316969729c2af389b5402ba32b04e63506fde343d3d39f9c123996fa88528a081c13585ad6cca15c341516569597621aa3f4a636f0c9ba0f24c90590922f9f378faf6f7b367f806208104fa72170ca668081208b5fe16b273a5c56023f04d2411af6f3984057b01fc0eb0d5df0ed72e674025d7e6433caa9c4d4bf3b3ef9a699f06a5fe90eea76716b8ea830f5062e45cfb1b8bf07db06ecdb0db610b4069ab6907f8f4221b94b6086ff72c5e39732e7d0891f3635d7b6a721cb010663d7469a3f3d556764757c2b250091e430a7ff5db60025a9e804b15833289ff7339b0af5f532cf622b10f791beca97bfdb25e2ff744e9a6c88db2f4b2672e185f92ea0455cc8df109d8d29a2bd0183fe7cea54c3479f42b04274e21f85cb73585b3187c8cb6275ad2675422c90d4bd4b0572c7e6688a71709bb3e0ce87c7374df86d2c0d90206db7088eba5f01f2a986400074bcdfdf3347318859945e119526ff6c0c775fea432a38346910ad6a29cfcb5b510d8220349bf0c3083466cf1c178ab3755e088306334d3b51dd5fdb809a7db260d23576c8b6a9baf4effbc6dbcbc31d87d42c0583d3f322da7749fcddadd204922c654685c992b9602178221757779e88fb25d233b2b98a714a9e932b8868f6c89edb6c5a54dcc72bd582492d24342e319593a5e0bb7b269b2eee96b3bfe14b03c786a1decd5d8cac19e3e30e4f0507b16b2130f47452154b6ed2bb73431f72010a2beef777754ed7e9f02604394fbb054315b63c239e9d4a651499949eb8874bf8602e22d158f218c8326591cebaa8701d232142508f88be1f51d15f93eaac3727ef29e64e79153cbf871b808a9166477511cabbdd2ba802ced3bea8d7767f09c792c2396e4466ad4118d343fc833434a2d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he9862f207d4e33893408cdb8fff85e1aed4b924e843ff91807ddb549a47ef8bb5d5f816b5f8af3c99c2d3f837ead1539dcee5643d56caf56f5d37505ea3934741d21cffdbaad623fe5248504aa81c3faedd902ac27180fb0b71e0f2d5d00419650150dc7914635189eb25e3cd32ef31de452bb2ba1de391a84b48a6177546f74df19f4543bb9f55f94aa5be5cd7c23b9cef4869d3123eb1f61dfd1686a0877b1b72171375b845c25481ccf987b8c333132b74cc6d1003fa7ac2aeba4cec48d7492b13c79c6207298af6b13ae9dd66f00569648c73fd202f1335c9da5e0643fde081896f7630ace7038790c39fccb304c5012b5eecd0f488acb29fdbe283f906ed7d6349cd355461474e87159f8d5c3e16e30f0d374ad849fc823ac4a1a9969daac4777bc5a3f5a764dbff5b299d9d4c465715a957446dae5119ec965dc813dbbf39117a4594227bf100a8d868435843edce7c14a228645e8bf0d0ff20ecd8b9b8289dc6e3f75cae0dde159dedb31fc6a40ad481bf11bd11ebae6394b3f37dd25ea70411363b98e367462b7c1f4cff34a3961db2510d5f64baca08d00829e5de7c6f714d08d86f099c7be4146bdd06eb5069b40bb0b956d4d1d6eabc15b9c3f359097ad245bb1f10934631a3a1f2381eef9adb9a2e2adcd2ddc5fd7f0893b66a489c24435ce2f7d052ff7a676bf2972bfccd6edb99059236ef5991fba03a359006ce1307652492da7ea8ad2d2f63007da1f4bdb50a375c96e64c8dedbe1dffa6d5ae262422ae70f68505e2ae7c2204034423976fd89edb4b9bba5eb1046113437a11d9374a06421299e2511bbad83f09d1ed86ae5266d7e4f743dfe2627ebb909a0401b1be20c68e3addf209f3c79e7aba137b256e72c64e9eeb1892d6a2123919639bd9690d4c50b9fa9de4876f8aea36ee9422f7c9dcce95654262db75966c44151fe395f07a2c08b63600da2ef720508e7725f3f7e1775b7136687ee55a92c595cd50826a8426232d5aafe332626e4d9f62243a0cd9387177d674b9a1686c131eceb7ee08fd41a365190d9020977112da1edbb2f9ca9542341c9d7364e45423c8591dd495a6f4f319e7c137ae9840c39a3f6df5d46546982e650a891074bec4e96f512e4109acaf53873a7e7e628d420dc26e5992c234bf16f03f67ae6e2b576263d1d2c242bd5fef6a6274df5fe4fc4c7c3dda5574f3b487a85dbf114d2e2a9381263c88e448938164bf75edaa511eb00b54da16ebb5683ba2d7a9c904f2ba8c39a1008f1fc519913cc1208e430f27e52855bb6f4b11c2b31844bc64c9d70096162ab5fddaeed3e589c1b78e1743bc9420f06a0ed9e4a0825ab53b0d8fe34b05962cfee452c4eb6765fbb359b5bb40f1dc37cb99be637f9baefcb475c99ee7fb4a614df0ab8b23667cca8a5b22f3c65474ca78022df544594e00e0caa48ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1aaf9ffdbd77f9c35f0ac2eb769dc516a55f7236ded695086b6fd126f44898124d269fd0f1fbdb7aafb5ae6dcd4411220734acc1c5f52c61d542d8ab16c47e4b633ef807c1fbe2df378cbce7e0393d33b3cf85d379c173cedcef019d2729d7ce644abc14a175a3152ca29c0f20ce4672d1d06e6ff595b8f0176a1c3ebfa27fddd5922dc45eb875c7afa47aef9678e91e42471f0b525798328a62a2d469cb5ecbc97afc0a99f7237303e9cea37f5e562db00f04bc1aa63bcfe2aef0181f6f96ba4e084a9fb3602c87cbd7e547b0d508b74091cf2cf9030d8f0ea52ace7a702c6ecf26ba94371df77c322ac87bb6107fe8d0e79d7b413aa2b6d1531debb6d883a80c4589b9ef50ff1aed11c510f0f0649f5e9b1555d38e60d3d0c0ac676534cce491cbbf2a5260d1ae19c8ae80f10e86bdbc05360764606683541443a39104c907ffcd49c3dcf6acdf0f38211322b562cc3b54125c72db6cb999a6e0920599ea2824c4dba6ce82ea3f0cf9cc3ace64cafbdf849a98b879a0cf776dd3efd10f931b899031b19ee06dd148aa44daade29bc2bf0eb9f2e78391c41c418a176f3614b3be9708f6885ade4eeec98fea833c3f56b01f540cb27ce60842d888017c4a578b37e9322e7a963ba7a0d92f366a28d55c7cb75b14a7f49b253b9c75bbcb0044836bf5e249f2e0d9b7e26d69d5950cbc78d4b4312729992b7cbf36b5de51a316396fa2ddaaae9c24060f16c898d7e789553d2c01bc07580c726c81ee7fdef359851ccde06dd715b276ec32774859ebd98cc1312cc96b329c0d1dbaac0313832c2a73e11bf104134603bbbe78898cb4a87ee5750701359261502a4738346b19c0d8f9ed0ab609d8a4987c8ed695535a4099a52f936893e6756be95a554121b06f8667bfa36c03b436c8b38413d4f06a0875fc5a12b238e9648c09787d729496779e6a0398de56d1eb615e75b51bdd16ecd499763135bd24228a28a5c934b34c2d9178b46c02a9e72f46e053d6219059b9f7cebe16d070b529ded25db13bea1b4adf5e740361a9ee192dbaaca888aaf7bb8abc11ba287a70fb9705f84d3cda9f025f981e6d7f41b147c31ddb6bca43193a6feb38b58c3d649a826b6af83de51f5dee46f7f4770074fa101c0baf09c3dae8ee013215d21167ddd9d1a967a2b34051d3833c1c09c9ab75e6f95a676a97a26d18fa5d848f5a7c00afc027eab4d15ae249f54be61e8e2b9611f7ee6dfe1212afcafb175ec9fd97622b48a8b5b1d746d3236193e15f987db45886dca3f1bc2c7993b6c4126d0e868aa266e4676931d058f2a9b4051557fc6cd2ec5105cfc13125a6afb1ceb1054cfb40d41c4884b8186c1a366613d52b8cba1056a8af93e762e6548229fb63448d9f8f3019b9dea964dfe555a6f79f7b164af780ba4ba0d4346c2c1c3a324623943c48023ac3384b8f0d9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd40e8af28fd2b64dc86be5d37e2cace9a9b45a5afaae700901f26858eebfba4fc1e66d67c3433dba008af660155269547fd1e3a2e2c9ba591cd2e6dd9b077204ae2e34d2e4584a5548b6b5f517f6a1a36593f10223d282db33b49ddebbf823a8b8951daf7b340209dd05ca9a73abd159eee01a3f913cb092ca056bc034b08102d6a41b61475b77dbfe33baf4e62e2a6f0f5b80b3b01e1e9ecbe7db97654669754ba6598331ed6295aa929658aa854ef83b54d31e17065686e6152057149e3e4b88d720694d69cf676ac94b5e4e6c6360c267ee69c3bf7aba640b80caa13e4a8d443acb07a1d013e92b2ab1d8298994c829ce7c1eda3907d8af9566d3e58d2ff00d76a3c7b43334ed0dfe1cb0969cbd6f371cd86f20d9af6a5f72e5dedd5ee08f0107ab8b69c5c7c17cad76b6697935fa894f30bc00e3fbf66178be4a63e4ff0f075d8bfc811485840300efe0bc5eeea6ba19886437221a004d9aafa9de8ce9ca42826c84beef619f8d40a1cd2bacc688ec95e7b4fae97ad9cf2fd8b585df13194287ac7527ec87ce685367e1c9bf865cae7043ec850e09ee1f47269020820d607725cac5872d54de304bbecebee76574c02ca0311e7c61e9a4f6dad7e3ea70d72b3600d612df0d1ce95f331904857477236add1ee070e6b09c4929693b688be217898cf6b020c6a0fce0dcf01622f2a9a3ed7ec211b57efa023d53d24f8612a3cde082f03001e9de1d8d2d9a239113ec3d9189050743eb74102969f9498002a52ba26ed8dd780955ba10eb9ac0372f6f3c6c595d02ddc4f62fb42311b7d0df8daae8d25d86153b6f63cfec03b343bfe0b5b8c69ac13c67f791b559c7f3ef21a63c0de34e154e83d48ee790a6852fdc857859970d5b4e48dad9682d58c4e12c8853c1b1d37e9753dfa0186febc295c5d4aa5db735f5bc6755b008e892154afbd0bee08055415efe16ca05e9b10e0517970b8cb5c653caf064b0f270188bd82b628b22f25e05be3f3d4c07d13435cd6f1a19f2bb015d7ca0d6fe23aa090f12f70a15a25448695fd5c056fa25f5b990514142b9d54e59f680bdc23a008ee93c329481b0ccf43b626e66e264156a63aae4e75588bbe4628848bdae94ac0372f21eb27480ae4c4abae8b4d83cbf9f7f9639475d9095a5a4f8b1f7bea05a4377c68895e49640de309ac01aed5cc317432bb033869753faba6192fdb8d5c10964c5da26e79ce49aac0d7b9d47642e5d9a5384fd341b1e0a185ba717758ed034f08de5faf43d8aa41b00397670bb7fd0bae64e9c32243eb415dbb2d692dd3315267dd31a2ac852484c8ab1956c61095ce3662bcd46222018f3688524d13a5a2c5b256c5818f012d2fe410d839470ead6e7912c48b13e2e2b65c56a5dd5c55508cf3fff3abbb619b3b774610cdb08201ceae460634ad7e08c9389e9fdcd3ef801eea019ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had584f06a8e2fcec2bbebc930d42aa5d8fc8e0f9ed5863f60b0460ece3dd8832e55a00e7afa92c804506d553baf018cece50203cc07b9161da7fc1de9e0a20212e6567cce8fbc0ccac48a201f40ad2f2bea8ebd88cd59ba17624ac09570d92290f11a3b799d65af2bb3d79b649d6e6ac9d8132262df99a6cfda3cfab46f6de4f617a9cb710429b84b08ff8f1b64680f749a56d47e8b9897da9c24607e0f6bf797d430741334f2588e6bdf83f2489d5a6196f8d45c78f6c7dce42372e7835989f30a1e7b9700b3f5e2cb47d77f258be7145e86752482d6d87577905a35635a3d2a089986b190cbd6666571d8f2bd04a867072af7756db695ba62efb8289f7c28de25c3e87fac67cd2532a12c7aa92dda36bc11cc1625f67a0e880e7fa8ef8f76625a473ac27bac661e342bc3ef60959bb3bb08e5cf22fb97f2e51ac93324853393a914d0d87c267aa85038c858ab9c40e21a273b7cbe31e2d070b939601b9f99b674369a676723ecc57f9d987098ab151da13f2bd657afb086e2dd31dbbc88d150d50451229ff9e1abf69717ab534a5f26691fc29816c961d4770a26ecfc5374dfa00854cb06a36e9260f55a316fd42d799a91e739d9ac9d210285f4f24061dc6788fdb6d254edfef407ef904fd0db8d6dcdd731b3c1c5484642fbf2aba25df0aeaf19c60f26f2ed9a214ffd7b1a2f6fe714577b03399b52565f082943d8ed3f1da04c7f4f55c222c636954a4c5be07e4dfcd520bc7e845e6c8803ea3d6bc2047071e5d4deb600bb0ee9bbc42cff5cc390ea9d6d98d543f3f752e538039424d5f20b412751dcaab3691b5f65e0413c7f47985bfb3faa64c35b0563c95fbf59da7b6e25ffe02d23e5e2c5eaaf1740b664702a840a0033c8e1192c4397ddf2173df6bf189f06683bba77061d7482c295a53653948eed4f1a6b31e030cd680d96b595015ec3f59f617a48984889b9aaf29483dccdbee01eb8ae7c817922a7cd8c6fe4413892bd935d48bec56010e993995afe4e21492f9b247e00c3c14acfc8188542a227e4e95cc8b9fd7c6e8ec51041011b6105070a1002192ea0f61e6772733da19140c14efe947f1071e00fb10d5102d1ae88e49c046ab1b78d230e3f9ad1c19e30b408a9ee8812711d17221b0064ffd6cf21120800ebb07034f7896851cc52a6d4124594c67499d7dc6cdffc7d1730def50d6a10b178a6210038e98dfa5a6dd538d24c777d1c30b97d5eafd583abf3901aa977cb10a4bec63fa12482fcabe95177b0cc0e004daf6d52a6884e4313dd7ccc9a47d8125b6394f16856b5b4b87d8f5ab730397575593339de73736bc59723fefb576cc5929ac2b9a38871a41067f638395f1b187fb7d3018092053e5aca1f796aedef492d4165f238b996353467f74f1b546aedbb829ad63634057190f2e206c2ebae25521f9dd52b0eb8747bb8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2424d4ad237bbeaf43b55508dccc6b8b5ee704ce0db6d8ba4aac3c62c58b1c89edb019ddb5dfb7a9b97448f082588e615a00a98593500d9e1ac0accd1ea397e46fcee99ce18db8ce9e3f2ef4a1e699532859384f5a0f53cd5d4e9edd7f5d213ff8fe7bc2aca143af68e42751b6361665600b396d341f67258fcf5ddfe0b76ec69d095fe02f8afe5e65264dbb20b56a55ae8a5615b9d3788b1f492ee5bd0d40f7b824244c393d0fbc8c6890d7be92e84c00d9d5e6862b029d680818cb733953aa3a920da60f788e0dc0be7b4b0d7c8a965617a7922c48442c5dd0568ff8f8d5c697501dcfb966e249ece82dcbc54d15a674085852f50b3d18b6385abee9b5412aad733a3f1ade14cca62075ccebd29bf536b9d79ee4024aae771312f38ddcbd5ee3640d2fb3c90125133e2f0a5d1c583f5fa45629cc0fc2285ab08227215ef3138231422fdcb1bc125a5aa4ad94cea8b4101f307944163c0ba6b0def4468be8a61bde8637c5a2b5c9e11f174fc65fa48fb9b8d2e8ac41211ad0192984838fa9ce66ea6908ccff23d71f81fb1b249139ad0fc2f564c2130ca5f0d3a9bc7f16c0921a1c4376ac46f78ca310ddfe0873da3f41c4012af162e078c81620e59c6055427631aa518cb86caabcae241f6e94089f3c15252795ff4deaab2501fbf3bc2623e59a2790a3401864ddbf26b556fabefabd25643a3e8fa200e5a893f0bafc290fe628b1f770b071ba7c11b039af44090a47bd3f261335760dc8a758064e4d7d018e78993c4c03f02f5fcd059e263dcd6b696c72c56fe06dd31b052f360ff33f2cf06858e76e06c65cedfcdf1b22721a587b9aa7b6e6bd62cab899d985c0fa1b74614c3a9768b9947b2f0152bdfbbeb02f433425523c529d157aa6cc7e1514e9cfe22b762d7ddba839375c9e40cd03a56b02a028727bd024f70e5a1f3d83624742a4d60f985ba2067654a20b3ac12870a6bf43be11b9082a535b49d7ebf4a6e2dab5b63be706e7fdc6ada67c1da432f6ae171c9bfee8cb94e24522f241869206a4bad1a4f5f581c675dd6c5d6360e33c021900ba76e73148afaff0181a959963699e325405853a97b31833df6ca2c1519063eaf761c61aacda139505d856f3814306ee7f9b85e653f5c400a198b8d82912677d31c2dcdf1a4e173a9edf570725a32bc11d26af29296e4f03d9e84af36b91e8a6a13fa849c59994eab9981e96aba949861ca3338754f13ec13b5d69d02d245ae7021de003656e9d322d5b11392259bd2ff79db500f7bd3ed1b998f5a447947fe33cee4e9af164a7901a9efbf787af435399d75f6c96f2531468e95e235598c8838025386838542e3f07a5949aaa9250150592d243759c6d5fb5143a6d7ffb4f6e3df442f12b7c51bf558e746e27a17a416e3866efcbe4a4012c1503f1d700affba459cdedca7a67f4c32af12268e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h596fb9c5dc2d8b1223b5bbd713f0f8d36feaf33f0d412bf8068007c322289a0a0fb0adafdb123a8a3cf6dbacfea60fe383969c0e50f1a1b26377f34a7c21d7a29bb9f19142945a10d1d3f7fb7ccd8ebb4ace1cff67d6e3ae0077d6293994b94f60f0515260677f187ad045a9e81a15312d3ae1ce3a62fb77dda7f1c378b415510c2430cd5cea23fab61d47b99b9dfdf64e622a9a74154b3398b13bc29518e07b1313db69e386cfb44b39f1a2b24eac84ea287d67b728d9809a732d60f6b747c5d47019cfcb4c5beb9f7b8664b04f34e75b017fe1942503a2d395234155945e34d04244a851566bd92020791e4160c93224549afb654ebec68b8e9ce41838cd88eacc50804776353db15515f78661064d251d2839d66949bf1887ba2dca3e64679e006eee3c5c199436c36a941a2cd90a5785e72bc8d0491db1bc406c0836edd79ae2c10bcff0c85b72e724f749411d9e3a42ec2356204a1a33b7fd51446833b4d7b880a24442f024c8597ed56d39ef9cc8c1bb2c1dd55f40eba5df023ead4c533fe005446eac1358a2427d7ead6a3cbb982277edb43d16e712f8a5f615647f4a1277fdd591148bd69dbdae7659ff47e11e0fd93ec627e2dadcc26b40e0d5ef64c6a79743d08e9844b78241c2f929f34acfc09889c6d4fc9c5f6333a5d3789b0917381e1acf1157627dc18cf5b60b71a3fd39f268c30dd5b9a435948ba40a7f8550143b464eeb1c8435c83c34723c6d1db8d6ca8d0b80c4d3914dc054b177642e2399beeb1d719e397309f975efd517aba6b17bc9b1c3e77e972fc92615ae3d9c0d326bcad20bcc7d694d6461926ce9bdb4176bfe2a5bbf2aa5a7dabc2341de71d9b67d02cc1cc631a3f7ad0607bafee5d866dd79f90b02ab277f4894743b463c27a76f643031e2d5bedc2f93eac371e050905f2faf676fc1ebd34cc2190fc10d2a7ab0b828b7877fa3b881a96bcbe00b497ccec0729a0f4c5803fcc007bfa78a7e089d39438a7024aa89a8e63260d3ab39e71b9d144e07e91d248e3f3d47ae049bb3607dd6d88d685c4e4e3c0e42271001ca782650d5a16cb4af9ccb35f4ad7ecb6791cb6cd2a9e93e489a514e1413fd086da7f64a0bed696aad487e83b27519e3918185fa9c80ac5efb8f1e5ce2046fb1d1f5dbf02a24153f467275dd3dede264c112f897799a6436539bd5b61d9e9039d29df803f4aa8ec33a1619b99e94da4110f3be10640f81bd78f7d3b7714a492da54a619104484c2141c8486012f1fe27ab8e9006f21267c23a243d10c1b65ea1b8e34e75565d1941a313e7d9b27749f9e040b17a1ffe1010f26f2f4755a3df00c28526be8b18745b456e5c9f362f84a2a619ee1c27477152430e8bfd057ce26bd5564a122fae9e72d797db87c4794972110da6ee6bb9ff4735c255bc71446fcecba2c6e0c878b670985a4d471455f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfdd7e44fa21bb8832a0773fcd05130e7e478c258a8b07767ad24289227de147d7d4f7ea0642fbe273c90b231e05537998bbdd0223ef03662bbcdbfc69619279724ede203c0b26f5d58baf07b71bf1b306b2958db4739f8a837dc1bea537424c82cbb7952bccbfe03b9b78c64f4e3e9e6803e85ac107ad8d716a48fb8674b9e09065ece5a8815d42b81bab206f0c9e125ad211dfdcd8200b3d697811a866eb677179d7bb5440e07f31d4b9e056d32c045d07e76c3ee961ef39e928077e18e873336604efdcf579229be262de7269c710c4d8464694c52f2f7f48e607dfa22f937f2a31e36c9c28e170dd8dc2fe2c1c751bdc5c9b4b9cc738f3c7e4ecce363b30aef10081c71540bea5a7ac121473870a8c98370eb208b09aff16aea29bdf05fd5d5f2f14fff0c665d770aa1d5dacb88eeeb50266d68189fa2d6dbad39cb31f6c51158f233feffcb87cce13faa5f2039e03465eb8c3aba862acdf39cd5b77d5a82ea2ff53a66549f0ff078758839467f1d6f3a9bf0052c497bc6b6d4f9bda6ddb3dabac0135b3e3cee71a8266dd89ba50cfdbd818728af65420ab9bee1a898467a2ef2a361bc95fdede2432ef16c4c8053d2c9e730bc93adc8b92eb90ae50ca140a99a038f198f6809d0426df7a6999c33bc3a2342698c507bf483972f09511b7036da78c1f9936ee67313261e7b71437b8cec23588a68e67d556e1f80e651e5cb9c71bdf1596d2913e7b4cc9e4987c0fe3be2fb35111fb302c14f09630d89c4e42a528a5b7269cc652c2dcf5cb1a055dc0f1d86e7de3337fc85432750655076a2265189e71de34fbdd1aebbb14cbd94a5e2d37f5dfae839b4d9a815b39c6a41e0117af110678addbdb8c83160dc138ddf2c99b98a55641d07e9b45f32034b0654a3c36d0dd4b087ea871f09770b569348a3c8a4b4f520b053c5a978a7ce1c5ff51061935d35f1bd5cd2bb443fac5cbcf804079be2c30c727d82b943b1b82dfe5423244991e90fe6b9dbd1398fa9688bbf61e6e6b176b9af3b0690083d6c824add7cb292706ca02e5538599e9270d8e5485380757044b7c263fde5df3f397b5e5f1155eed96607fd0c78bd6b0782e2ff89263cddd9748db3b0de12847709ec5ae0e55c1bfec0e6a74ba871a51f2910d5d8b5ad800cfb84d9f15b44693c0ab8cb55697422d2f3b65f1495d89f4bd5a581c8c52bc102e398ac641e5518d5ebe5de9b0acab52139177c7b443e2323ab23a42a6a4763e5c39a5763cb0e0cf6eb805be559c7a7065c122d88d1e6b1a059b78577c7e493c4f741db459f451d9e08c49684923c921cdc1547170a97e39a83989a881e030fd2f06b8324d4f6425b9ccb9b65588e723673420bb567696191331749c0acfbcb0c8e46ef47fde75f473a9b86a8130371cc5b3989d353937aadc388d80eff043d33935dcb6e9689de73cd22f650;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'haa2792e58aa5446a35fa858572a867f5fe327d12aabef4ed7b66f570ba4379c51f3e96b03e1077123da916b00bf68d6f2362f1b6906c7272b044357d1e5bd6b48eed269facb7a6e9269bcec8b36b5877ef0ac45b24bacfa65ee9ca5463bdea3ca3477e007c7ae7970fa527ea2e8b2ec118b039b148c8c0a1e392f6d4ed653b9aeee4c4ad6c6ed7abd521c2345ca3453fbc223ec6a13ad2f7701a7a2d4eca11685066e16dcc572dd523cd17f6e0f599fe59b9e97b1b06059e29844adc63f7bc47d6bb2b29c68035cf1c436a331ebc385dfb59ca9591f3b75b3cd98b0448127033f00ad4eecad78c499c48a5253a505f59fa506a137a8f742d6f3353f73c71d7c99d585cea5f4c273c78c9ae0bfed4b7a816ca4d80cb087eb408cc07828c7d1a7d92b7b11b6f07ec94b60d1769579aa2e5161b35cd7fdac48e2ef7ae01179f20a9fc753ecc588f404f75ca44e4ba5b6d1afc43f9b6a191157dcea39fb7d382ba296793756153b48fda397365b8ec6425acae134e0cc80e3d0e449b9b9956ffe189e708db262354592a34677c853ad6a86437454ceb48038ac22de16b7202e392a36b6d4665d0353dad9372aeb49183faa1447dd45c9fc927d88816b186d3c07687cb5d938fbafefb7bc2cfccf4a718e3ed0148e5bbf1035c4bc74da035bfa82e5c574adc538ffeee0c0e1042df18930557604d5e21543e271c9584ef0f8a4f3af2470829b01528da701c6e61d9df9dce6ac5d94ccb3c954c14acf7decedae5a9eeada472e80ab9d114bfea33824d3b155b82976a292b5f707e4a7a8391554c5d6f4278361463d6fbb65acd4786967b2304cb74ffd4a871c974cd64d333c69fe3bbd3756b25897416e73f6be101f1f3449253cc79c9798400d069013bec20fe3fd2892a44c54eae7a73b08669e7294d71c3cb6948dcd6630f4dc9f5c7fc6c1f633c52c9c6c3793afb5e3604bbf22a9919c35b686ded38e3b20ec5a92c9ec239021048b1c8b6deca4646705f45629522afb1d61cabf5b6af6131abbcb277dc6a7a8de4337a5ff14c20131cb242f7d65ae75f3a39180ef9bae34bb76ec0901c62d0151b3254ca45b2ea54b8d98fc7217ef53968f7515944a405c7700037189ff6f3ee4439bd4f382602732263a5e0d3c027a635347a0e91b27fbccb690e89e1c5d0be65aa266688dd401168d29a3fd9e680af432fd5c28c8958aff2fd90fb37222b568c9a7e9d2a70b1f92aff616015971016762955b25caa99e3de32f2dbf59423216ba8736e741742a9a4a8ebbd1750a82a95207ceb574779590becadf572a2a8f413132317276e9d0ebc6cc2eb10c1dbf7d5b94125fab31f84962aaba4bdf95727039f3b54a3dfc84592a97ed7a875b62aff0ddd94f84a17802202ec64bb9dda20249e4ab9c20f5b952e84a7383ff1a4f9e587abf0e7d39eb132271d320208f741;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2a2105cb1c6863bb1bf94435d48311561212fc24787988090cb3368fd83357c7238a167a19a38048804b76e760271a9898227a464e73e6c858835fbf90ec7ad94955e89d3a88265bb4e86caab5de3b1e972b899e7c32b3304c55e040978f506227610a26576824a58ffd7e4aab89cce64197b39d1d47175e612f202696e8a8138ba62bd7c94d573b27dff2eadbfa153d0ff4a64fa702856ce3d6ed8dd65c4a5cfbfee68b5ed00dc37e3c9f73b6b78076c9cfe759b9a625fd8f2f37a88e854d9383d56445a6fbb26935d4fe75d27aeb9ef56967106844cb43c94481d3bbaef7d9d83af8ff21825651df5334eee1053c4cdb5233fbbc9f9bc833ce05cc5725853b09cc1eb13802cd509631b480983ecec5095839fb9348081ad80b2be6e2b0b005bff538828668d401a6692cad8205e5ac0a7b330deb87de8f30783c8ec9b93551a7e8a1c72df789aa349daaba43c401257a0384f36708f2332509942e525beb6d5d964a9e5e5e572c2ee1024eddce49b9251b471fdf2ec721cf6f3e8c8aee74210e3058c28a0d68e8b9d745aad129a307b7ef1aadd6474cdc902b5717311bc12e1f6d48c21a40f947cc3296abbf4909726fac7b0f47669889c43152903da9576628187864fc8c24daa3a3d3c65967caf7b08278b3730500ac3fd5602b172a0f3620a048098ed14b10ae4650596ef6cf3ea6694cda6831bc5ea4e063504583284d842c6e827fc79bf4fd5032da35df356307138b02db1b245edfb322f306221d710b3ebfcf95dc4e71a0ecf9bd6135b522c4ecb21f61e2433c5f3f0c550e277f6dde8a58b09dc0a47f702deaa0fda8e089ff985558b6ca6bbf75757ae74b10ea7ff0ac28c8ebfbfde24953d4d146e28f7f10f9dd9a3529a586352488f6d80a0a2d028410bea5b1a23d8a67ec505e33eddb9d348a661c06c9e2dff627793f60e684d7b221a9187e344c3ed996ea8b6affe0946205e696a3e572f858b9519872455b11ad30d45a641bb26859e4d28215be0f5f90a437ceff8045dd094a04f04d6b708044ef243fd0ac8df6aeb95d692ba12eb6d3070e326b44970eedaf8e6963a9d753f9391667cc03635447cba654db9863b247e8b2612163c7e13fb6db7e81ff0fb382f102662c4181dfc56431de0547bfa2050621ce026d92f5e388d7828482411698e29d3727d6e51e76e04b74438936e508fe3e9c017fe5edca2ee72b1f4416cb5cf620acf74f30e94b62d74bbaa279dfef590eb3eb9d2ff9c81977a16728930bb57450b7c879c1bf88480a74a9dcc5455ed7aff42204e1ddc496c4cf56061e916def53a58d1d38b690654a16a474a71ce24495f7d2e0f50678ae9cd87ce85568cd9503648c59fe8ad43f853b14a21dcec8664626acb2bda6dc8edf69ada36372af3e125140da25ccd3f3c979e4e0d5760cf1ef9060f5956ff34b1d1b600ea2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5693e2b522f7dbb1c7401a95e9979ff1a9fa4eac2f979019289aa079db079bc3ca76de0a922ce3bf4481ea25f8c94c8617aba14c275b80174bdd0d0578282487895f0c637da1fd2ce935b24a09a8da9ee283318ba2e962a4c5ed97c4ceff722f5c3ca62c8d593b9ace2d5310bbac9f9fc2b98740e58236d0d3d67c191ba2d778f7feb6f4330d083a1f43949f369daf5ef0d7cf2064b7f95a35b8448a62ca3b980c9160e0a3e04fcc702ccef06123fce04c0245af7c2241eeab694fcd652c0c07bb20fd1564068645e28fd9ac7abfc18586786d31ff6a594a4030a3a93c240fe2872325b95b30e77c0167d03067fbaa37233551820617e76d73965db7587e537f9cf03cbeeecd0952d35099fd30fb4461c80cc1bc9f5908a5295af85eda0afbb08c91d45eaa41befe6286fa0f5a7b3daefd1936878889a3a711d04d32c1099f3f77dafd25d56efde8553f27bef515442689ff83550c58eea547822c16034e3f79f5a35a7f34ca8ef3d36b21da22d06f40ae823959778f593cf2bac2e73b27f8499ee1b7c5795fcaa772918d24082d2c964301f70cd04e75a47dbaea956a7956f64d1004bf593fa6c5a9874e426ed63e41bb1326e91bf55574d68bd49cc4398d01783548600daca60b55a731bd5657adce2798740af2e6a01bc2f4a3988e760601ac4a90c6d79d658dc508d054676d05f7fad887e92530a78e1ec4ee4b47fa426afef22ada5074d90dc809221d87ba0e2f45afefdd27f8b2e0586e8b88489d73ca000218014c6e9605a1302263779c7e96935231ef8e6467b009ec2a0a1775db8be4e029e442fa63dd363f4a2222bbc570c9283a8f43055628bc8e8ca32ed940a33030fbeca98a3acfaf0af6461f9ec7606bb7910f9b45bcc74e6011e959293b5f08110895c714585bc7330b612702bf3a79110394342c1b4ec1a9da7c720201b79aede66af053fc4dbe2e7b71d391a41e3015d037c221798737c4daabe94504c7bb6cfb8beb33b6c1f4a09b84f72db92f0f392b9cd2474a685909d03eea75355562a424e024407c828151a3c0d8ca8d0ba2364f78da6db762b505c2d72c9575b7a8578cf0ee6af1410654505ed6fe3bf193429a3d1f9ac8768e434df85bba3a0bcfecdecccdc51e875cf27549d4bb6ae110a7c48017ba856f94b7c8e43e9d5fbd3402bb794c821646924346bf8c423387a6c62e4bf6c072521fa59c68babdef9c74d6762801b2c1b6f29e431a43be83d4a75950edf3a494e57295fcd849fb8632c103423b6b0b1822cb2d85341501c5b85dede72449cc661914e9135033fd40a80c6e730884f0c4dab820f79f2ca29518a2d697e886f4c16ece22ea369facbb6e35951f56ac052a40e8accc27767d3afd035d9ada4567a01d21819afd103041f0fd1df284109d47cadc3493ab9460e735a6a3149c2157e14748cbfadf8c25e6ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5d2247bcdb075846e93d1a12a0119493e004b523c62a63ab17d96279251143a8ce6b33f449a7362379d50faa6f77b66e1a3f2c236dba638b4a3f93d78501c3d77f94e46a7c00cb51e0b694a3c73a8b15b989e40a823fb34b95ee86dc5727465de324f04651d0c3c61c5152483d90c4d9e853e4692840408b3a44b0e13abc0c93dc775329627a02dad1df9fc58fbe55dc9d48ad4130b5bbcc3594253a88a4c316d9374a7d062848fd60fcc730ce10fb2dd4629c2c6459da55c08a9bb93329fc6d7f301ce6bd0203e81fcda0b66b959af8d4099647efa11a0067f8e29585c36de1148a4fc526d5188087b8b0e7af20be06391356b4e6a754a4ef91ad6d40e4cd6c630830364ea74dedaec064480d38c193a97b5b73a1595e07dbf673f24fabc82a2a0ac439218da5e9f9c555147709d544c85ea7383651c6b2d54711dd1b2d46135563b53a8681c55a90261faa1e9f726cf4a7e04930d4d0e9a0624fe3df752cd00f3c87f0354b6468ab8e2322c3d2239085813847f3b5f47baff5b2b0add48ea0ad88480af0c7191a9c04284162fbe5f8cd2b421283db8b0d660e4d79203ba7ae030ec224411b3910f2ef649d089c166853f2cdde5e3875ee979b768adc31aa222fd78e3d12a9b1fb19d4ea0b7ce2e3b921eca9bf10f47faf0d541ab087d9576881cc814114a7228d3b3b6ba1746117e4109215b2e2ffd3d8060158c49c209cc43b7f3bd54dc8ac56223b9ba0e8f25283128681312670220aca6c7fec3046228449802f04298490eac00712ab0c52ba3d2b9f2d30c757014c93d3159da0d50bf8945745eca8d91dc375a01d4d02014914b750cd4174da129a8a28455a5f7a1823a356b5822fb6cbbe1e7e12d5f1e806b9dd534219c8927432ea94b0269906f3f098f2248a9e974530d7dcb557cb8150eb9644d4aa14498f3444f80faeec1ac959ca4185fa75b5c4a44a4c5f8279765d889125b8a510da08e67b92949c72d64e9c0c4142738c656a269c10a824a3d28eb521c99ccecb3bd4042bdbebf3f265fff03898dfe2b804b631d2c81c3639b6b32d81d81bfa446b3a85341ab37041ceaea22746f0b2f48fd3d940fb7e4b57bd64d7e488a15af70fedbcb89de5f2bed31360b6da48ac319b72e7fd6861ab8ed9d1e72bcb170152aee61157474cda711ff7fdf3b7db18ae9f685da0607c4771ad77c8e6f25ce2e63097edde3a78837a719bc143414a687df3d816ac7924c6bf14fd8530eb040a8df7960453fff594439a22eee07deb1262dfdb6b7bd5076188dbf90193972fe82185ae2371bc09afd0a28a4e8e080186f95ae4f2f29969ff7887c02979d346b7f2427a79bde460580dca1ee5c538bbb5b6245cb52d27e2e989fa3dc89734ff40b063c48c257dd5374ca9a75e9ddf5d7db41a030578268fd9b3b9ecc362b60809ce951f877e4e6802c1703494;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcbf7988760424a1cccc7cc9bf02f98334491adda36fbee94ef8a97ae3960bc4d5bed584b4b23fe8bdce87e6c90cbfb19dedd9871c4e2dafdc15fb219cc154921f409b1beac8010708ad7cd5a9fc932cf5971c05a8bbd4352f8ec916e719671fc19964bddc24705fdfdd6db9edf0000924a51fc853b7468919e79012959255023426ea90d8ec41d01740e0a534b1edfe056bc5eefe6886b10f59f835bedc5274c59798abd5be6a5b97cd5cac38101fcb26571d56648bd935640ea258ec294dcb558c4e3abe89d8621d76b8cdf5e0f4bf4502085aec2935c2a086fd6b31578035cb0e333948f512c4f4de188bda1f9aed03773a61a9795637601639d58c5f0ffd5a9dafb238bc57302eb66527f55fa36330ad89c250485812b3c81cb0485e762ee32d90946d2ddefa327038b73ec6e4e912dcdedc8a9a39aa715465c746e1e27106d809d97feb05b3ae5dd633d1907f8eb594b7939fe02a51497420ab9bc23e86ecea4e78b96c265a5df3260aa1f0ffc9e3a1feb9c75be0c503ff8c2153224ed48ee9975ae16c784e89ab26d7201480563679e9d5c8bf8791533788c869ca96c657af7d9997fdd4a5a35db5f6735968c18e63b95776da98da09ddab8fb1434c2a5c42c2fccb3a918b8cbe4e8238bb3692c9e4e0b633378c24bd113e3404d1c2d92cae4fb24fa6165ee86ad65d9d9c950ad9a262e8e76e9a7912c71bb79b8ce36fed74ebba5af8305ceac8bf87fc16fab74123b2f38f8564296a08a4085313529bbc39dbb080890a21f505a6c374c3fb4154ef37804b223f4a1975afaa621508f70cb7fc79d5923c0d336f84ab81dbffdfd7898883e13c7b2dea0f74f10b4a184757fbc39455ce9a4b7c77265aac06bd0cc814d0c69dbe2ddf64f12179a1f7b5484cc468f09b573e2745ccfc0ba4d00bd7383ce71ec5f293c38c1879601c208c45462d5a184ef08c452fc86ced49bc834d3b3890257abf3ce2b58bbb129c891c87333811570019cb9d69d6f0e99ba1c3f662d135261899dc84791e81a22e1ba5c3545770d9646e9d98fdf21bd67a9120c9058e55814fc8f89f1d008c2ee2445e3ed2c0cf64e101ec489615af9955b5fc24709741ab0c64bd6ea049505d33e1b67d0e818684b72762e6e5e4c0494690346d1f630e6b0cb649f24f4991227a006bf852815d05c586dc18030ecedff6b706a3803e4bb9863328408d7864d745585b14a7f0bdecd3b70cd7d74d6caad17b96cce45f928f44ee198427ae73c41d1810edf35cf04d89d67d07957b5195d34e990d6b658ac8fb6d06a6f012bad1ece5c09f72e3ff3bd764df326fb00c347bf28346dbe5c5363b1bcbeb21b2eda6e25a6433f496ebe8dab292b16549618e57d6265322e5b6c69e41818fd9f32bf701f48f0d39b673e5dc8d79cf872e2f5942d36d9bb6efe7ea98714083d199b35600f737d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfc752da1d903c966bf78a0b1191cf72992d10462a1c5956118f576565a59f2047044baadcb308bd309e491d3880691115d86fcfaf8c543783e9a9c5a39b686e26a0526cedf8eacf3a017b785cdadce4aeadfc2f614dad81d63acea9f0b43d3742042e74fac076728723b8454108c15c00f3cefd0bec6a59758a65a7067f8f430c5b4a184c474d19c428571524f03d205aa0a4561bfa76d78acfe0c18f88a26d54132802789238f63c50751341d522481f96aef76db1b8f61591b5d9ebee88673a86533a1bce06dded829fb395b6c7c01c4d71e55e17bed01661d40572da2eaf2cd43f2fa23e83ffb615bf83573130441c598f7e88793655eea11143e3abbc53bcc79fcd50e0d3c8bde8a1b70e54cc66d5c4e32da6301186b2abecfb22a14d9d7f9546db71e2aa27a0bb5640f2b3ce2e9be3ccd52e1de3e436aeed901d3ee5767d0c7b3fa4b252cfebca68eef1fd0ed6036e25e8fd065b85f6205e16985105211083cb7d3906852e4431a948f444fa4a1efa056d5a9856ffe647f69d51691fbcfb313ea3bb092ce1caf86621d8d98a213abc4b86ae01595a1084effadacf33d0ee77b682142b221ad4b30f9cdaa3ee149e0d71c90fe7fc5f7cda7a5f1b306dc46f34a11a9ebe15d64e3449afe4d7b4472f99ae16dd2e1141fccd4df345728d435083dea47d398f3fb58345590e35fa2673d000734cc2cb090023d0ae295c2f371575e7e8780147616621afce1f1398c916506599d020cb0c4481a1a1fca9dda44848a6bc998b37a261e05d1310d87ebe50fd67a6771a8442d2f520d71c1dbce300bec36c51f3bb01ed2b751fa44b627ad54cb368ed3acb98245a2612d517d8adc73b9ef455c045fdc4c0d98775ed0181fe4c5aa626c668afbb5dc4bf90eb69047d702e3c503f8713b8373d7590ef2ace2340ea37d58dc62b3fcc21a61110683527b6116b7f678bfc1a3630bbafabee6247670200feb53fdc68b3d3046ff7e15607dff834e45457585eaea6f3e5713ae2469b30a215d5f957b71fc6ae9adf53e6eb32e0797200c4618e8a1758e62a3c90cc90a653325100fb5242cf611ada2c1b92bd7f1ce50f847a461420f54c074abffc020e14a64648d0ad53bbfed1f41b7a4323c60472199aab735accc1f6dcfc70476b0e8871452e6709cff8c63849d255317e370c35a1e6400e183bdab897b14c4f0ac87b59839d7f04b4e9d3318ddb2f0650340207ed0b33d9a322e65a9e82e64a0140c0511314fc1a03a2c087cff785f647082e6fda6ff9e481f99f8a785c43cbe5925455509ae66b13aeb10212ac377d26a1625f255125266f513036b9d489d47e81090e79995856b3525436bdd6ab7b944b94a5623398ed75cb4fc053becf1774f45e2f0c56c90b10c6b67e6ff707545d5d6f83b4eac6256a119a15d711522f263f5e4a94b14b9d6b5f28f199aeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h330be0c449818ab398409cec7888e5300d1d725f511058c76db12693cb5ef0d57f5b7274084a0fb065e5df5ebb5af0f3d0e8851c0fb8e05f8847fb6633cbe84daf50f3f731fc87df4580c34d29c97f5566c30810fbd146f97003c377425917b48603ebe3c506a40cd288e4a2793f0e9cd506dc1b169347fbffa1cececd627bbb6954eb77d3c4e9303773fdda57bfb3e17061d01fe0afd993cb6661c2c7909202fc011b48a740434274999734675bd9b19f12a1bc2b36829047b474ce4f7945956291f3512e3f31b1837f57700146535d5b833a20a9ea43729f4479e7c47353b0add8d2ead38187f3ebbe8223f125fb37f99005531f5ec299543c77f9a644ece6bc53683691b46ba20304099bc703085148386a153fd1e14a5ca0e40bc83c692b084472127b275e8393ef704ea67b8873f875bb3b4741287e73663fe2e7afef2e2d13df121ab5417f98ef23f3d57cdabc4288b8e98669b5bd40d5d75406223690bc26074d29be980761ffe09e86113c8fb173a44cc72b7e05517fef7d5cf77f3dc14d6ff10301bf14d8260df45ced5ab96226a869e70b93dacdfd931f14b03557395f9a7f90cdbf4de3a129810d25b518502b7315eda9ef9cdc9405246bd3e51fc411ffecfca67437730215f4d562691ec3dec9cfe8462c0606fa2fe041ef36032ead67a872b1bf4f8807a59963ff997d8a1ce713049632f7fac937ad09baa0280051f8ca0ce78b5e2968fa507b65af0dbbc18799f1ccd6240abe1028c78af0625bfadfeff8411569c719da84fc86e6556c3041b3109f8d43961bd49aca7839947d14e0a048503cd101a122327b87e6c3a9ff98895dc8b36a529faa3b782d19a4368a084fae2f42c1bfcd8f109200a19a3a0d7f3c1cea1047673f0aee595819b9f30c34905efefb5857cb0da9af0ad16381aa55c74781db5201b519d8118f785ffb5dfa317fbe4f8a7d5d8c54a454f6e88697c64e2486b8b452be483cba6f91df95a806bf0a063a05fd572cc390c38a8eb2ca99ce49c8d2d037f68cf4e7d73d5d4c74e6cc48873ef2af124ca60d78136ee8a57de89dd9187695e12a486662898e59d724aac131c42137c512b28f7c4bcbe6348e84a0ca685ccac9a9bb305d6c76f97bf07952d433894acd51ab09e28c4f636fbd7d903602d2b4afb56918374b15f579935c52765b9b19490de398170a7b7808457e42bc96b5f0021e6e3d20e4dcf8b603d62554af043ffadb411d8e05f9c5cdd123c02f3839bd4be43cb685c7ded8f2dd974b91eab0059b9377209302ddef75ea6930e71ee4f3806b174583c47733a8fd1072b79a25a3b9bde0153267d498a67aea93b75020f5b4daaa1b20dba99582a4c4eac0e70f724fa78ef209d574f52fadb4c2abe494271db9807e0ab7c761c6e7dc43bc83bd4b80f08608f48c25023e773b5f6993d9866f3559551c15cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h17c6a1eaca633b6898c8e85d12619fc9336940707276c6ee08ff2223d90a213f892aa5a679a7084a3d66bd365ccc7ce5f2a26f27bd1a6f1d1bb55a42527f4f4702eda9367c1380e932c69734f4568dc6d67f05b8b5e4aa434b4fff1380ff56dc05ddc9670ceeef5d4ae3f97a00c94d29445d2d1fb42a68c897174ec2b98a3f50310c17db57f3f2139cc95aa05338e0e7264f2b44337e2c41134590692f945086cc064e312fec9d255d17b1c1b1221842eb4205e67976234359664a5cad94c29e139e2bf3e11b4ee216eddf4b34adbe7411985ddc5aa16b9fbbe68141df7156844a28923e5070d48a14f05d7d64b3e45b005685fc0f7ea9916bd12e7a0dc87b3f6b76f810069e4ffe86dadf1904d013e72701e5b246d6b8add681af9ee13bc9e4a3815ff80304180d152de9a5393e0c94231eb023143bb0766c00d67d3ca784348bf3693c2c96a1f2be6fe0f6f2c6b12ea1739fb7e772942ebb273610576785b5e3597698e9cfda65a833fc32ec256c48faeacd2a2b026353dbdef0a0b96291ccce9df313c0b64eb3f07fcab3bb838f048383153fc5d84b74ae0c2406782aa741f2d96fa9de4f656cc1c030de8556c20dba8ad657df2c9b01203a30c632fc23cd69dc45fbd5608533091fa5a711385ef5883346b75d0e22d0cb7e2d250fba9d4fe5f0ca54337bec1d6aea2bb6e07659d7e58ea942ba283ab178fb53796b23f1a4351e38d1224472967cd614761015f671484d413d83160f154744ca075f620e44a96c7d58dc9a0c8736f3dbfaee0f403d614c788e86c0940af8f41575101da91ca38eb053455878fd3367549df1046cca1edcd54c99b2479e3f3a639c2b2fb6f280721a198b55adb5fa781dda6fba5c99e9e0518925dc25b6ca26624bd0823eedbcf3dc91c4fb7af329b49d52e5fad388ba618711d873eaa346cfbf1485cff9df8e14d86b34e0efeac90629c862624cfd501185b33eba2a12618ed904e47c419257dde66fa387cd5f32a2994a40c227224014f766ed2ae5bd893f368236306b3f8309b3652fbf0d68886b9dcf0859cf2810a37967e8756c4b903405cbbb0e6420cdc9af9cf539438cd0df98f7950c491a63c8114fe462d3fd4b179347f11b6eab68751e7a26d76dc668de395759cbf0554e125d0ac8f41085fcd66bd5ec6f9c50a9f5fc55454afae4e84f758ec99cc9b67f67c96358b00db38fc602767e06d1704ae51d6dc0ea84042e8b778da71cf5a83b17303e8b6f73014a6c6171b6151a1ea902640950b983ff536a169d93c0825911a6e1901df36e26fa637abd8472d8f014ef439bed9524dad15313b568d4b3126e1d0f0bf182d47a15d8f8613db2d5d271122e9a4d92ef8a08e38b630bc5135ccbbf990434f2d61a9eae8bde3068148716bf2f5957e055d291ba2b3007cb5c40d850d2f1b1391205b60db519f6fc3d02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2014b017f019f6994942acd6b7db59f7be4a5afb324be4bb7f75680e2c0892ea9772c31a9022ac6448b60a137dc62374a254e54bb51c25a45e52a7b90cef245efcb0f3d6cb85f2f6b5e118bdae23b643140bef2ce07972109b3b99286ab17f66ca57a1bc3b10453a020489fa76c2fdbce41c711c4af4da124b4b7f4a800b2c4153aab9a57202afe1924b52c68f14cd35014b21c5fd4228979f28b85ef4eb6a26310a584e4e28f8c6d587a008ea4daf0398ba8bb9425ba3e77888e64ce7f6f893daa550681c0e32eae6be261115e5889ae5246ff6420d460c4bbf09e05518f721694b8eb215a2a5f3574872f01fd3f2a73363220565ab840dc6c8a1dea1059c11ed836cb80f70a46842866a647cee55d791ef5a56f424209fd813029c2a883f3881107bfe8d9e8f209bc9bd118d098a26c8c9f1451a015a28c41b31b71a9520a5fba09be04105bd8690d2855e8f3eb2c1fa3d0b660fbe73925384e7a3a572a2bccf3ef944829753e2c3fdab70d0358941fa3aec5862a99f52706efd4a214ff6ff4f474be6debb055ef2b3b186b899f233e41b9c2826624aef8c18e4375458f8b66b76f42c4a658442c062789275ad77c7aa558d0b76f252b9cd06af127b977990df18214dcb232eb1880581a84fe3f6f8e4c937f91c109a944530494a708ed2e253b690ebb20c278270c42b0dda68ad75af884bcff529ae0123497b5bb9670fee3d9059b52a2ca168b7366b3804f94088714bb8d6405bc1ead073015349c0d7f78b4be5e16db6423ea492c082e68e1dc92493ee3cd17936e043859bf1ca331ad9e9076e4c75b53acaa4473e51ea086fb0aa1f254764ffe4accabe36bae86dda9cc4727f20abca2abb31c1a48d67063381749ed9d27525fab262f8411611d3a5e64352a134a34074581bc3e0ba8f14f0d94af44e57a0eb611feb67e61a7dd99d31227dc9058d22801535fc0d19da8ea54a577a544aa682179821384c9c06493cae1a7e98e4d6f44944523bc199ffc3aa237a07f8963dba709afc7efecbbbab8de88c89bd667b757631ee8136994f50c25d8cd321fd9c8bbaaea014825490ddd3799afaa96b5a0bb3b4aa9a3116c24582bca034c911375b383fa485552ddaba31d2096bedfa57eaaefe191f7fa2d4762a18f120117891ba1361165f4b4293db49ef3b9ffd0a03616230e5281ec391a890337cfe69b3d906aba3fd3ed6c96ef4319bd42ae83d86b5e27580ee2d35ecb0f3c2f8ab14526ec9753cf314ebf3d4ec40c4fb3bf2393e2ce21fb736a6703002f52216c4e9aed199d352dd4aec5c09147cd439c20b5fb83625e4f26e142e8671f7d145db77a9b4cc811801d3eeed3ff46eba82c8b993d893e8d6a13385ca8c3582caa8b5c43da3595ac058bb7a3013322bfedf9af6c1f198f2e7c397903a95b4b8685cb9bdab035192d760c0530d66b3484c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9d1628fa460932c9faf6018f92f0b26a9973ee5f9a05e13164f9311bddf3fc3dbec62c43c2b2b9cd995b570b48fad13114ac74018abd491a6b7f2320e8eb9b11b55725917f2ee6ec4342301f2fa3910bd5a892f5eb71a426598cc33a7a95a186bdcc2e2467bab736560b945b0ee8fc2ba0c64c2dbb73f3317bde3f804ce8fbc8f5a780b09d899e3c734e5b47e901c6257b450975d3b5e5a992a3a046e6f1a7ae98799e1937eb000b1ab484efc1c1d878ee982e33b549cccb89eaa98413c23788c0a9abf64b35a8cca5efec22c52d291a1d0454b8b3dd4e580763384a2cc3d55c0cc48a225dd4c6a39c13534e05151efb4fb4869c0370abd7207964ade318e98a0be9d9c3d14dfc6eb7269098292208ebfd7c074483e6f274792155732c3972ed7a43e4384c43093a2765ca7341ade77fa96b78cefee3998126bebfdb09a6980a44be88ffd67c599df3b40f094d427b57f131366b80a5a6126dade4e30e7ea5fb2916505a6b977c12acd1e6f67148d036badecbdc2ce4ca521ffbb01805299773dc9e31dcfd0d71198b9855460979bab5f2c29666b8b09c0ad14f31a4d971d5f21448ad7aa171a5a6cf4317cec467c6c650fadbb913349b06af5586ace6177fe9d3a4702cbbb4c25970b411fd63ca94ac5515bab2ef426b348def25be0402290e6c2d52eeddc297417154393734f45a1a36c169f06da2e32ed08a24519447682799ce2df6d7108b944c6c7ddefbdd20c0c9d7be26f463a2ea4bd8eb5deaaa6e4e99e32ce1d4a7152ab70a9fee37e025afce4e1d527314a827b4adf67a1c4541f82dfaf3ecd582517f18d99446c7245cd01af2334c9ad80f8a046bd3494957a31e497c38fad5c054ddbe5101af4cb6378fbfef2dc164eaa0993ee3fffec438df7c9b5ee10d519c80b7a6fc77fc2894d949c190425f7bb101a2a55455a9c2318fa195ff53ede2412f815a697454ae31d69fba3124babe681df23119a52567057c68e6e6b617da69447f272d0c22927a7ee5b9265168a2916877f345638b454bfbd856ffbb910f4453c2d397526ec63b280a8ff4a0fd834288c30c13a9df4b01c7331d958039054ec29a57c97ced281e4215aeb232c64c1191ca8dcd53a2c0572619f33588062d1835f31c0d2e4a9ea8b1f4923a91c5daaeafcc4463ab97077deb16463d64fbb13859b2fa226fa4f3377a0741828ed73cff30a2109ba6917ffbdf11ba929f93a416f162c4d4e8f4821f6209a0ec36a2752b9098195fbb9147822635db2b2ba187e00508fc2686cc397b926a287c53bd0c272788a814b756367c77e0a00f762715274aa521fd549b01d8294c8dee52d01111d77064c899beafb83f04364de5f1280827ca18b96b1a5c2c73e32925dfa3c8831abdfd579a9eca634d7ff9579e95ad953367cca17f49e46cadb2bc5a6aa9f825499ae9a14aa06ad326c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha89e40b4d83204b396436a83fab0eff394edc562eb1a980ca495f84737477aeeab1d75814898c235826f6b9dc58a9821ea37350ff34b00ec71e0d2e8f938e7c6e9f773692a747c222bb286faaa2abfd0b1433350fbdcdbcab00246d253a24ad2e96ca32ad6628fa430973477e50e5d0f7bc8871e2851cc4ef6eb13b08aa9a99b55537a25dfb26c7312de4360cdc9fc2f235a45b4a0002fbf5ae906f10142fac196ce5017196091f0a34a10b7ea7801acdc4c2ad3fa9cbadd1b0d1c3353b55ca91c2df78fbdb00b0ef80f8327ca280f4288c5bb2b13fa945e8a13783ffe54bda1cb91b483c6f2a413f625b029b1068a47272d10ad237eacd46c3ee21dab9751d463352be8cee854790fe758d946aa68d9447ecd9d20749eb620c226961a8e1c824d6573a0af6ae839177a8e77ae8cbab9bc6fea1fb8924802922ab15d8bb775e2decaa58e18c1dc5cf3c0abbc23256eded795a5a922f6ad363e164f3e162297015cb6cd9659b3f7614aa6d79f6a80b3eb353564c7e7a966a69c6a0f0105ddb28497a931314c8c58dc9fe037ae93721561968f905aa36966dbb77daa7df44324d1c391a8f0924208ba4a0df2babe882a5d4356128bc7abd72b4c86074f526f8a1e580c0174ae0626bd51eaf9c4b9a07735d05e8de1c66bb553918bddfaca211f7ce12b87202ac39e3157f494851cf81294b0a59938b4b443613a35151fa3167582e46761358bbf5f2a5d844fd74f2538b6cce7187c38fbaa1e6cea12b6e0a7b8503d59137c5f8215e938285b48398f49d728f0cf8eda2d8742704d1e09c9bee6f173049e29cce9cce8d0e5bf4e8aeafb2abf01f59c0ca9ea88931223901aaf41998641b47a812b588d1307b00f33dcd6a00c598fa2f225adb09c3feb0a2c65cbdc1ba19a7e9ecfca19d17813b7fa97316c80456789434cd9562008d280f9ef84d3699b9acdbce413e204228597da10d7cd347927f1c6bff4a4ee21b8434df324bf1681f67aa271eae71a6ddf3c974d82ea7cd4a219fa69ba610b3d67a6cc41f8ed1f7a2a109b7b9da70c35754ed7fee0781dc7b9862c428f72e7f38cffd3ffc199fa88377ba0574ba3a2160646e4e01725e74811759bec2313268d59931be9d41f03f88e89f9cf7ce2d3e01caab2c6cc5f7222ae08c0bd410a6439d5c2a384577a4747b71adde523d3818824ab0fd6dacf6135a3b4796a407be59c4bed9d8abbdbe25f0135d11d0f4d6922b859e0d5eab0c4f0fab23df7b19129cf793ece06504048a6cdea6078e52593d2a17020d9a8c904314c06bbd9dbd31a53e4e90130bb4f2d7edb7d899fa0aa97150d88001d4e337b5989ae76329644a530a8f4186a75c0863682cb0ad38e771cd7a9d43642fc6e70728b13814e475ec46ee0c3617a993f8bd9e1e9a3243589d3284d500614fec40dd48d5cb5f4d3146b59ff9626d4f5d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hde1db43d26d9b3d3a49816de71831ccfedffeb49e8a4d8189a71b0592318df69fd0c6afa3326a0f0ed59ed557aa87346d6e01c379d45f46e8d4a262471504a3deac5624169b2a931d3fd3daf8f1d95906cdee85626cc9d6948ca3359c2eabe0363e5ec42dc328e3544a8b1a9c28c62d2e0cc5839d7065a7332e82d21300c0c473ace413da6da28fd2b1bf74ad9dffa1e55fb138920268718ff0d19a41f25f318942dc5a01c03e6b4ebfa9404efdad1835f4cfade55f93eaf6b671914792565be302f92f9bebdf4d5b974afb09bc25a359b007635fa3d2a3ef7be5e1e23f763a31d0b04a38798d313406190cab6a18fc2c8b2ee4ea3f7cb15b2c836ed3d09bd9697f848e285d7979fbc134307cacdf1126c897fe72868d4f1df510d970b64f7a2e816dc19cab8d0fff14d21b9c9419d5652bc7ef20ea6b6dc14ca2d848cfdbafde17f1abce19bb9141e0f52dcaeab8203232b19723ad5fca39abf95506de29439da6f54fe4c9bfb4f9377b12b572672e35a38a156593a774ec9ee2237593c38c55eea1d08e48a7863995470d8a2a02c206c56033722073a8f31a36265cccc07ef31262c81cbda2c478e5cb64c249118c87a6f76a27fe4c8fde2654eee8d6fb83d1d764d192fba08c629409b0594b8765ece64d0c893c72041736e3f075cbfa701a1f756f824f18c25dffa292df0301eb7e9d8891973682cd500528ce9ac8ed53d729bfa88075c3013bc1ae9b6150b53cddc414e047630fca2f1da4fea5bdf688fff8de77cc2b578a740fdf2b75ec530d2dfd0b1a05e69be529312f51f6bf2413fbad2e49b6bccbc1d720350a53922b88dd07852d0b0e235e0229ee4d4afe6c193203098fc8e616ca3e55de45dcd781dbb0caa65c1e9f55bcacb47a713882b5f88698a32c1dad3301858bffc55b1763028806549be21db9d5c678ed127eb0638302bb149a1f8fe5f3f448d1f34cf15355d97fe528e6ef5ac4f658d0f27b083e87af48c5413abc044d6313bbb69c30444d326d85107089319708e43f0b0e0808795cb9464f961377bb8e0469a1bd03b6ebef7efd97498363c70df9bfad1f21d252910196c6527b867e214f0af9287be789fbe434dfc1247437957c003b7d06cb0a8609ce904211084d3a4a92ec51c6d342624a27fe39e540d3d4f584aa9938404c5e81c001194106231f3963b50b2d491e8107035e0995ff1bde4573e331d02b5a8934abf15fa0b564a151172eee3b38df638cfbb2d611c68b41b728650fbbce3d3e4069b884225c1c8b1ba42f353cd64eafe4457493e85ebc5b58416ad683298176c2b9f8bc877e867edfe163b28b4e473257dcd5cd7bae4ce56faf05de8725184380f00bf73ccddbc48110b8e005d6c23d13f5978c0c5ca6c3324b3f293ebdb4569030df330e48e2fbd25eeb5ea0e1c3873c9238b8c7f2fea8a5dbf920c01855d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbdea6063c11d204c9c3f2455089047560b3212e46eaccc97a63ebdf544668e6121a0fd29e295bf8b4da54d7a765dacf27afbee3142405e78586841849a7716e22b6d29a0f890d8a9b6f939d2adbb2f5b97372fe9b1a1afbd207fb8394e64f1ca5985a3c05010312a21cce6cee7b0af4a4d55f8b97371489dfe0afd186e595857986a93de77669b6b57267ecf5a97366b5d4e590098ab8ff71609460ca06b3dfc6477bc319a43d2f286bcc8cb73d4c8536bb703290954ce203d3d5a6d61eb8c9f24c445653a165fd1962d152ba4b518304f06b4bb5e13d3c1d93f1322a3c747a131581c493ca3b42ad366b5a760bbaa5a9fc0149e5d07ebf18799c3d388d83df4433bb8c138759adef7d234070b5cb182759f24c644048d2a5bf76181b4af0f0671dbcc960dbedfec17365efc628a875e8fb4d4652e031e7909e449f369114654b2a1cdf16cbc3366b913c6bc1c8a126da7889341c81be968bf3c61abd5fc03125aff34d74fb1b4c21c8f16b83eb6ca0a504435fc3bf82921c5a23fd1cc11dd399db4eeef6da2971aeaae12b719cd46031db94e09080c37f8c03e50133bbba4a74edd2c84d7070d6f668c092abecbe96ef911b1ec84f0bd0b89b318ecd3763317bf8789e9ac547fe2198787ecac32acef87a4af5449abda5b7d15767444eca3660b21e089fa28cbc71da96ef36e2d96097a0e58257a59e05b66458785e9d14139adf45de7bbbe3f3d38f61ac80f51210b90096ec8025dbe5d9c213c7001234f2207acf03bc222208b26a7c531f6554922762f4464a9dd18c285e4fb304fdb80a4c0f106b79b33af55d3d932c6f43100f39163d84291bd8203779da36b3f9f51cd3ba03210dac40b74a34ca595afed4d7ee8ac295347b05747598b49c5686b105e6b6371d97e27daeb0aabd38de52cf0408fed317e7743ea411d1abe1dc54d35bb1b5ba0fcecb88c34edb7576a35b2c1a56be057b23f5da6ec8aa5ec1461cf2a553d4cda264d4b79ef6a25cf8f3515b3386fe88a1563ea11d1e4bb0ceb1286a28a36e480be99039be4d5e7d001648b2a300fd313d874173a3d605364374e7367233c5ca5965d2b6ce29a50321ad571c6ebfc7fe7f002a3298d392d43ea1b08e28030db6676bf7bd307654d8f4140e763eb6d11d8d44b581cd6f88bd516d1c20577ac858e9904c18764a415c44d4db9bb65ec752cb1a3bdfdd47316a4dd73394cc1a0357fa90e6b44a9e72013400a5c85f36ae619b0195af4bd85ddbb965d2d629ade3233cfffacd385a251673ee9b7c779693eb13a077262aeb4589b4eca09cfd6e4708f49eb48b04e621b04d00300c35386aeaa424f59b260b85a38b4ad1baf57965d7422c8acc0e02560813d3681d82e2e5df98b027c62c19731b0926886feb33bf3109d4c2124d389155aa1bda7af5ab58980ba464e6c7629daf58701b9eb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heffbe9a925b2fe1a1dbfc12e3d7b423769eab7a1ff221e652562c8912d381202907353a0e5904feda2458699e426ee4be03286c0d9a2b750c0f7a8cff126bcc0e3e3881c9f2799db97b2865c939d47e8eaf243fac3af0aee27f039048b771c36907f6e86416dbd785e4065642e5036035144c86421a2183053e45b79334352b3ba7a9f0630d4204f6ab05e8f67ff5d128bdcbd473eccfd16d80a7774a17456c8be82fbe424ccb0dc37a6d754a0b789f25867ad749e73ea9e0121d44d0c2426d4ac7fb60ba0a02a0ad084b6c288aad7cff8df5b6395d873a7992bb323bb48d1937b86af56533770c58cf248ba057935b5f2980146e0fc2ec8f2aff9f2490505d2e554d49cca66e6b7b66113d0f74d2a9fafd39d5fc6fdd7fbfe994b7d9ffe3ca1bb32e5b96e330e1fc36b8a9561425e9916f53c55844a28905bffef62c81065df5ee6f0cda261dcd20a8d8d83a8a7b69c6ecb0eab1480d24b92cb0442f5e55fb61ab59d4e87babc2afc118fe2146187cbe52135a913b05327b21072da022e766291fad4fcc1c163736192faec649685252525cdad132cbc7375d746dc8fdeb3c1f31cfa01bd55a9f0cd75f018b28615ddaf31cf102bee1526d717a5dd4ed69f771e6305ae0de0f36aec06727cf60ad530ef56929ad7a23dc9824d46f92268dbcde9b328472a122a38ec7ee185a72a59b7f797e8b398b57b6c6069c764630ccec5f3c7d6e050ae235445d30d675b305bcddb8ce18561c942937ed46b5c9f289f1be9b2da439d0080709abbb44b8a2adc50cd1bbd2c853f398490135df92da05c92ad08c060814942a74fd0443851767d94d1ffaa2c77bad25476c20d9465087a303b804015ee205bfcbc925f7f62cb4501a12676c2d22aaebe393b8924fe8ce6df526ea695e19799d7ec6115b5d8b3c1048ba6e6d431cadb52ccdb62e946db029b9949b91bcca67fbcfc8dc3540f05363ede499787b163c5736a1d440fd9ad31d4b05d48cb4e883a999ca1836ccf714862c2c1f9e9824044345db783c0b9f02a07b2438a753f9b83915aae5779ed444a33455eeb7fff26b8b99e1fd90c5b981fa9882918b1ad788d73994e46036c227c1a2859a98844c4ffced986e2d8dfede26e3bdfe03aac364f91afde4ff7b76d661b9d846430ba3b1bf25adc6130b5bed14771e87d503c1e1a25b488697c39736b16bc5fbdd05ab3e6a68407a441bf0b6c61c134c5923ca52ec465f8c3e68c9454065a1c6c30e51dfe745cfadc02d4f896892ab4752e6bcf175b881feca289a70ff5d3cd457e65eb4b087f5b669d5fbff3a053b708aa132ab0bba92636ed5c24ceed38921c43c6fb4e216a6e73db0576195d7db985ffe583bc0f72b3bc52c30eb9e01389e1cee49d3551f729a4528c6d33bf65b1b978ac84b15e0c48c473d41e46894625e064b631fc44ac562a445fdbba0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h10b519c031caf3a63f23e1e3b74c3a96f6d0bacd45cb373c10ed3223377aa5a565bb39f6c3664bbdf995a606b1cf3cd1dc13515bc6fd7afd57f6b152792fee27bb9e5433e619329df0d18adea0d983d3da72f79b05436ccda2c4fa54f495c5d62b3a5c67e96bf20f7fffadef83f3500081ba77182050281685cfb503c41402109ccbe790b0a6ca5a072e6036c384507045e2102cd65d68d2d32ee99ae5e8ff3133455654fa577f0eeff85f3bb53e5469a572d508aec0081d3ebc306014b375fa006c234a9a8651c13fe0dced35ded743fd77f6a0b80f64b0d1bcd0dd9d5b4b239da187f2c7fce58f6af47fa373ae28335b8d7ed275f45ce01c7c50463c3152c2c98b377b264707441cbc655e2d0d69099facca5c6df069a13e728d628101657b7a89f621d8a721dc9b55d235a2165d68de17f9701c54344c4bb8257e8b3031a986e410e74a8575cf1a9a4b1f928d4132035ede2e5047f92bc539e0ba01e1d904ef77c613f7ffb553bfc2fda2b3df4bc7564a6b50790b9afb69dea655ccf7497850bc14a0802982bf6d9dd8d35d78f74f9e7b0732adf19f283208af594961a87c4f06f9ea272f73758d1a0226e0ddabd0ce2d98784d59cbb322b7c6187cc7ea9becc324e97ab081fcf6be4862b5b9d2499bde9d0deb5074188989a4de27e30c2d8b6f7b425e6725916f143a16e0beea992118f1363fdc94dae7630e92ce74b323a396ee5350fb4fb736618623bc272d7935b11c910579cee0c63a10bea96baf0066ce21244db55560860e59df98b2a68ba2a8c05cd010f1988578aa279f0d60295627f1a51bad913665825213f178f6d6ea6221e5beb10cb3093a54a3b77e00cf52ac9868c3ae0cfdc4944870cfb60aa3093187fe2b0c52c3a2053932a9a89c827fb8d1b93876a59d7261ecffb0293f8b59ae58804989ce147263d9a1a2f7b95e20ed826fd674fd2cbcb2a6ccc93de97b24d22cee1accb74889d445834496a26f67b17d3fe9b8e38cd22584fa53287bc999834715dd2d4ee21fef602399cb152801ffc05fb42b44bffbe771ad20f9698176bb7c1bf0a44893d102523cb67a617112195f9ed24713bcd7e585b937907156d0a610a939c7727cafb4215f16907d8d230732e46a79bc31c6ec5e0b83f8ad0460e9c5d7c56eee3f98a7a671c515ef61e8392e65bf4bbaf4ac4d290e7dbb5c750a5aadf582114073ca39c16f1a92e8458ed5c34b5a26f7f1c1261881e7e2f881a53ca78fe9f41a05468fcab13a99f124dd2a28e92be9dea3bb2bd512d67e1805f0439e8c133580601b9b9b5ee2dc818390bf27ffd88bc601de2c5c8b920d6a117fb66cedb7521177106ad7a19cab651584bf7928c9f6badb812c93190e1f12c3f03e65dc82d86c62a55fdbc01ff2ec3f5fd4071891445baa5490abbf5f39a34653ddb310926c4c8931926bd53de75b3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8649999c321f499230184c28366f059e892fcc9675418bc5265b93e7ec1ad2507782450c55c314426f7e16333d9582fababf2bdbcaba7b2bc466e4c4f38f79c2ce2693824e1bcfef7ddcf29dc179521671e9c84a830235fa336520e96346291b6336a795fa7e94b56636648483372164a616b884d5ee3b40429fca34117aa67482beb2e47a8fef6865fe22e41cc59e9c5bcd1ea880cbdb0ac1e1389b31e105eff9292cf5177b6a0c721cb67aa41fb9661f6612e80c34b2a969ab0761f2665959f7abc2d6c661008cc8a0dd744dddff5407c0167a3bd010fc1e24ed925f8d1973166c009f8ca318317b9ecf6241bece2555a1b3012812e02c9556b87e78add364335233d4993e97a652ebda41a04f6ddfadfd1cdd2106e90dc555b023b651cdc86d70e5698ef7c1496f3bc24772beb912e3fe8d96ca42124f50b52c2d048a24ad10a30ce67ac1db994f9025aff92b17852c1be45a93c7670f2b169227219df8d753d149bacb1ffed64070c31b67e1307d44ea1d20a8f3abe0250628ca3e19ed55850148f354db5e48c49b9dadce27b92ee287d54406d54391e518b551c653580706a7cafd66fad39bb343c9d7a54904f89631163bb09be289df875428e10bbd1944b23fbb5773e6bc741b1fa77b6fa02bf23ce3aabee9dfd4775fe0f759befe9599753492047759732fb5745806d701844a3e693dfe9bf480f4ffe53da8db3df40cce13bea09adfef59bc59ead9d480aad218ca34c1866acace975d592dd83a6766469238e6af4568bbe42b8e422738b096cf0f7f883d3c3ee188a0a6263e31de79e05b01e30f2bea06ef76e4ad92114159d93e16a4e95cda25d88b8bbd09af2461c3c8dc10792dec0f7cbb06139fe92b460085b86d1b3925d7539ce5d5c7e4bd010be8469bc34bf26fdf1d6f94126a402d77f9bfa0657df4f6629ccfce53238246de32c436bfb3fd41c2a90726b6acc59066ef424f4fb95075e5b88060796d71259921028e9539114757a7efdb92032571c94f0eafbf67254da9f020acb9d6832a5266ca4bf1dd496a0ea10299a26de404757e30392f843a0e5af60eb72a41615bb2ed43f41307158b5c4b7be467c8dfeb4bf0b7c14026cd83ce07add16164ba6a4216786c4fcbcadbacf89e2365cfe8aa6f93475ad582c4e33819345ccf7b5ed79e831a476747ccde8bb837d7f4cf4777741d9e93a2399b0ece48b357a79ac356288478875466d44492343140e1c8b7d4ed7224dd5ab05e4a85769923d38e5b50921c951cb45137008f1b1d7bfe53c399445c1772b3ced72ca0d88123c628cd2ea7f69a47e41ddb3abc13cd609683e6fc8d0506e8bd35200f9c66f47193555d4a541f394b63569768aaaafa586c478f74fddf3a1abb869b6be0e322ad2e12ff7c74833aa4fa983682b3c4d8e95ada18f7efcb49f5f003113abf168d6a52dc9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4a15ea116389516c9bbd9b17d86272627d423d81d9d2495f68b166f959a9e421733e77271d384aa752ce9e85b432762c94f64455f227dc54cfc16d047f557c9ff37c937c5eb0672e68337d95040e0e91be65251121f1c2e5dbef64f6975e094a5f24164516993828c33467da20590518ff4a92d0412e5f361299e87f5f85f4077d2553fe97b46016b5e8ad5f949655213f377c64ccd945ac3cd30890342a990fd1da3e4188adbd5a05988e79070bcc5a92e361e8feb4ecd51ca4c805abe1a64e952912cbc6b1c11c781bd1a13f1543d7a31736f4e0566db5b5bff949b37c1c1fc81dbd87c7db716f7babbc35a5b870e424742beaecb7a5a386ede9731f7a1bde9addc991c091b64d5dee8f5255e0d5139f1fc01bb27ad1c5659aeb515a881e5cff3eb9713ea742d83e0375a3ffbcdb1c4ed612eb4f78f422b52617f35f9d82073803e14507d5fe6b86933a76ddc292f66c87ae7756d38c23864ee45a468880e3c0a93bcde8f6e70ff218c0ba8ff068a7a52ae741b039f31f18686935eec99bac5a3897c38906130e901011da497c6e2ed71cd04e1eede3c306c1b945eb7115793a7888e9dd0ed3da24f4413462a9f2a06ff648d20805f6cd410caa0e002f83ba355c725c8102c1e4f031e66368eadfab5dbc99a0fbd3c5d569f9712958999db3fac7a62ed5f6802434bf74a854d3cde956a53374965c7fe157c0a71120e6488cf3b3af2d8b7456b95e84f6c83a6ccefaab88579cca2dd643c4d0f9005aae6b7b88cef9b5c0039cebe7187c8c4f237bc54d54d7a6be931d0dc20114547a7f1b0b7273c7223baa387d9ebb10e168e84012bee924069692dc700e510381661b9f2a1edb5da584d867714b24b9ef1d1478a9777326b765a95831203926b2f3a4c135da840d20e589ff76c34b8dd892975e5f9a306334f349f8e5e6c7a702c2f6e8ecbe849346cf999d22e3b5208e29f3822aff57a2cedc261b60cc101ac0e51c2e4896e00936387e663a93dd0050f3afd4de0d23536751a5febddd219d3bb276e00bf2ba1b36051bff262643a0f72989ac6cd9cdc19dfb8cd90577d3436ae42e2c7930eec5e13d1b14e079df0df5552b4425d72ec03ca24544e33c58ef466f2f857e9528064a72217d4ce79abd3af21eff37788e3ac6df90b366f4fb92f3e0279049b7e3c4c9435a579e1ed3e833c0ac5c1bc6b4b3690d3d4d477b17e93f93c20df74b7927e6468ca7210d2b1666f89b605274ec699d90dd687a145e975b7888ac33ff12713ecad47a90455dbaad281cc94d28faa2147853c0c89b4ba56a88dc741f3377fae62b0740259694d13c95a47a7fcc25c870bdd7edbecc7e25d1df16e31af555fa5b993ed4e332ac3eb88755f72ca035b40e14ae99d3b857fdc8cfb012c0d5834c3209dfcb9cb31c5383408ae172347dbaefebcc112c70f01ca6b270fa76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h444d6effba1f709f40a836a83b96c9602c7297d0881b052639a9007843ae45362ca080f87d5e8488594af1a9bedfc5de8e5495763fa717496b13ab258a22a2ebca47f87845263147d48e446947f267b14f72c168db1784f8ac9771c836248255bd9945c7e5bdd7810a33004b3effecbff23a21e49f166b2f02856aa331e0c58ac72e975da9f461facf0cacbe0567d68afc0857a5f5db44477013dabf9a00ce765737c861754a9b18aa77387c9df42ce4f91e676504e672b8e3313e6a74fe41246c146d80413b4e1d7bbd0ea04c3b83108fe0c4d41959dceea64f6d2858f8a2641c83a4bea7116bc1286eddbd9397629b441b49b64c4a585d04be84c7a70f28f1c68d0cf0a89cd73db67bb9bd0b84e4fa072890e003665c0a89b23a9920017e75ff720099a1d7116545aa23b9d2ab1e6264099867a6f61452814318edc00a9e91a4bcc3872f93312c336c919bbcf7443b21e4865ae261bc6e17215f2a9b5d022b0110bc15d08401d1bb1db3f1dfb5c9dcf142e9878a067c4da2c8ff5b15fd5407185eac7880dfab0b028aa171268a3391f0d23becd544caa084a517367de7868f0756574c711e3890b4065cfd98cafb60a89ace43232b94c3a04d0365697c15a745caac432b2354c77b398e0d99acc17bb082d9ef82873708ef0ed011467cbb754a2a13ec2499a5ebebf9385b4c55cc42bb8c71e1901f66091d8e61c0dd92f9a215a0b31f5616b67b3724637100d27a515c60e5739a1be242a19ef941601459ad1b719fccea2509b41083a89c5f4bb50e8478d636b2d34e3dcf37073ff5f9bc5e26075cffabaae360836dd72dbb56aa272b6aa7d8e84bab7379abceee6cdfce10f204d2894e9e6a4a6a92b462f39a5daa0a28fbf405449f057282cb41c66253b685624c60215702fcbb1a575f8fdc56e15ac68d3e7099266f9f53ec75d30cfcaa1475e4aed6e154b08e85cd1e9c060bceca3c1191aaa5eabfeeabac04c91ed275097dee3ef569f6963e72f85bd505a5cfd6193e17f8c316a83c223ee6fb9d83f4103dec2b5c7e30158e1b1e2de3eb7dfcdc09953f760d6244e1ab570c2a9d3873f64d40b9703bba1ca3f99727bd298231b32ffa8275cd94552745f9ddb8a93bec32543ef62119fd62b2bc61ce3d6b7d48eb89ca14fdbfd354abe17a3bfc4ed3884aa3bb0c3837088c8e5910a529869153f02fa334861de3a0111dc61ef9d16619bcd7cc50dbb84c6bc9d90bb1d0ed0c2f0d3e5b976d8c4be9d7e97487ec11b88be981ed04d7092d54fe1af465fe1288d2cfa5e89316718380b27df65c6c0401affbfccd407181e0971d74c6138cd8ba033485c38150e6f4b71b2fd1e598184aa2868e710bf40f60e6cdfc9f696658e38ee76e1379370f5e48d6915ae4dc3bc28e06c57cc027723b2071716a8cc028f445725e26670c1373ace5aee2fce95509c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h32146fa581309470e89b5def157d54738894b93676213dd2e89cb798a9f31290d75a8cfc339eb05ca08607306fa8f26cbb59722fb842ec87dbee993cf8c1143a6b764bc6fd00ef4b2f1f2e12a470a3236320e591a4ed2c418d4dcbdd9b29fe2c941ada74a90817ace485d10d1c86467a991c41515625b8a8e574541805797a64dbe6de561cc5dc56b9cdf0efc0638083a785d064bf7b0161f900904fd7260fe2486c920176f0e7b130935ae64a57aa7409d0d3adbc9561a8e1246e94b2a74ffa62595b4208f5dbd707f5cb0d296fba49f5e022a3e0e5ab42de1553b5bfed13551d9e9a659ce8d711949f9bb63f65b58ed56764e924ce5c97a2b7cefe63e4f7fa429ad2e047ee3debdd887ec934a123b82b9a4011f9e8d9a7247521453866abe9aa95a4999d758311055cb902c88700bcc150dd34fa8aebf3eef495a5595907f43d02f0326b09729a4edaed8d47462b09d747c1f684f725b162d160a140fff16de883661ef547bee50c9f884b925d60eab800aaebb607f1d6b8bf1b35dc4a29cab7bfdbca61171adea047640c1313515cbc5a2ba2e7957c469adf10a31b6cb9a259b89bef7b93080be826cf59f4b3284cd0becf5d7bed93a7deb42613dfa87cebc87b46d10ff936ba17e976b727990ed95324ef03f70b104f61826c1065a15a3c28ed3693644873f0a9edb2db17130be4b90caa696086a4811dd56eff8e8acf90c1d6604304db0553553696835afca5dec65825154fa9cd39de716f6c609c4c237cfedef6dec1edc1f8d2289b7d5d2003feec6a35c66b2a5a61f939eed01d51cf3ed31652cafa3b901d55fa753767395bf762f272c230fe0139487e5ae8b827e5f56f063a154b297f8ef478d2752a86fdadaa2f7a8508d3f0730cf6a9e9b217f12e2feda4969ec838f29badeb6e2ea6f842a074a54edee2b3072ce324755c8e2c66c79e6c15546cf92a47e055479d6dfd03992f123ea76ef60d725d7dc4f128873f3749659fb1a9ebe102ea9ac4832ed9758aacd8927868632ee2eeef3987b8a32259da68953b8b99f22e2501258c6f97687c440080b29a216c56d1e71253c750c72ae87453795ccdb06af37b520e729777eff77fab47ee23fe71f56d6ee7e4387c65a66299b65faa8a35ecf738e9c3d95b4f553b0e08f96f2ff69d2ac16ea6e89d97a6c542347f02f24bf089b446561872192daf7de22c5c847abf89cf4c587362efaec86f85766e35216c2f56a7aff9394de2b21f659be8213f6e30a3785ed14e9a5a9a0e8d096a13251790630a844ba0fa2bd0cd05a337328887eea07fd7fc2c59a8ca51ffd8b8d97a5a1ceb8f2cbda4f9ff9b83e11477cd14854862f97568d660f4d38826bd3dc61301767fc6befa460b6d7597577a3fcc04c14d1add7d31efa6132682ade53fe301ac350be334ac8478aaf938d94297f46c7b81781ef101;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hedbc12085c9ed6b8e229daa5c97d212976dd54d45c33b6f7ac84f588791917d4c7b955c778d227b858141911395195b3d6af6f6318c68407b77ec3a83a8f1c20f76fb45029cab70d3cb564f9f89b72c32a2eb5856b79ebd971ce29062fdb486d7a58c9e7f73cfc6f184c9451272ce3c2c0658696cca2f936eeb2e4f63d8441ae57941fe45f995282d370e5c1c26effd21d47571bce5d5b6bad6fd86d90bc1936a095739afaffbc01f3967be8bda81da6554a6fa35ede20508613f9f4095340a3370f0e44c270c02c8ee8cc418c183be82240ebe8908cd66bf0cc563bceefeaf88d1bdea29b3f7633baa72967fbc0724c4749963daf68ca458ed20c7a3ba6044287ec348bf46f10409a4e296ffa40ad3cb2b9857b9d617911104d9c5686e4169f95056be67d7e3de168c9e9f4f74e5f5a9166bead6abd5e0437f8d7ee4ae002ce500ccca6a8fe5aebffc2f251c9a376777c1897aa7b2c0b0aeeebe85fc1d27cefa269ab44e7df7dfb2875acb8cedfcd21cf149b4b938aca8ced973c8062ee5e89a467997e8c226620bed496d8061bfe9dc368032a9618365d0399046dd6af7683602ba6c402cd73f0c640833e1f1c848724c86c7409e1aa92721cc2019245f981c59f2a89d597edff74759778e61cdc9a49b53590c6ecd977061895c2afff3f109c32c5f66e3bcadedf606da3cdc1f3260033e60f8367267fd9e3c14773a8bf0e505f3ee5c9d4660acdccd0391f7f85c4e19683bde2629cdb88757ee23907474bf25d0660249488e7ccd8cfbfd8b0ca85a868e0db71590d5aa2511d66329895c3d9df785692a1a9e241ab1c506b383b3ed7924f0d6f55e29b81cc09d3a447a96a2b06b9eec274ce38288bc3d1da89c5448c72247c31c14cfa7242ffe55281b1766c5d649cfbd92ab92c5b08152da5abce2df3c7294f98f375ce7bdb6ea8924edd475b7810b90c0081d2b2c063354700eb5931551c558cd02a76ac26dbeee145cb00a65e547c6c22c412e26bebda900941e3235ca326caa7c81efb4932976d11b9306952fc5edba84885f0ca350103b77905d4f87f8825a449d3e84d7b67c8a4d3f926bb7bf8e0d0c6bd5f3c1558fc826c25f00127e7a8fe7da3541744a62cc2fb787f6d5dc4e811f15ea2ab86f254049e7b65b412d634992f3dd509cc4be786cf5466e44b68fc928a7c1f4f1a5d4e741a5833721e42a523bcc0bb75467f3a01f7885de6cab66accc5aecaf9f52bbca8bd29a6c1baf0fbf91de8fe40b3660f21bb4eff87878aaa633349af18072d65b190ff2e4e427af7b95286264c117bb7496536ce64aea68acc1db7c929057c0879e45e8f0817d4d9ce885c8aefd84f7691adb0bd9f0085e29556e661618edfbec834a0dd94445a99d2a2653aa579f0da384ac3ac24c2ab883e67b200b0d3ec45c280bdbdabfe7913a7041d5408b1dabc8411;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4fa493cc5d13574daba90f2dfa972d3233e39274921742694d204c860243cde0e07e823faa7b1c9af0f6ad09cf8add23b24f50ac0c40175c69cb8f05ebb3e8ead56772634e73ddc12ba22a7f275103e2e0555c26990fe69e056c9696dccec187f3a9894a0620e36d697a1a0e9641954cd83a1b7cedcdd5cf093d7be3a0f654b49573e79e87144b1f0d019612e1c5ddebdece70731151fb8824abe3e7fa6597d2d7cd26f1ee346240a740b4138be8d50bc6e8ab08efa88e49f8fc2977481b739ef62f9d89bd00e681ed2c863330bf5f39706909192f101cfdcb811e9411391a598d330521ab6b99fb9edd9a7ddf36aecafde9e92b0e674733185fa8e96d8b5e2daeec9cb08475172c2c8f3a16a08b0672c334304049da7a92c6ca4f0c3a9045a4ad84a2cae8268d8cfe537d05fa60ad4ed8675e52d915742d5f74cc00fe94ad9ffb0869aec5cae6009a20665cad6385762b32079717d702eaea4f0da59ebd4493edfef1dc1b5730cfb0cb57c6d7b2d18df95e53ba4aa35a2f258b66c59f4dde92f0746dbd33dd37b513469453edaa5f8c0fb8ea9736d0ef91867ef7c6f5f4e0d03988bd7541b7454bac132de35e5eda905cab9b1326575fc2157a62e9ec6b8883b3fd66784fd9af14eade8c9df98440b1109127d8eb6da26d5aea62aac8e973099e176eaf26f8fe6981c03edcecdc2d385ccfac79fce0707149f7399f8440f342a67c0e31835e98ac6a2ec9a49169e472ba737de15235d0ca9a79bb0a4c5298d87d80cbbfbd22a6fbc1a5844d586ab21127d957ce3a143c149d2bca166a2c5439ee44c464326ecfb665b7004c604e7c46e00ad5d6a4426ae18fcf22ad780bfb8dbf545ce73195489eb9a5163c6db26df5c8acd1014d36377d6e8a42989143656c885e7361ab14191caeaa9651824011569d0a37f0ea70ee1ad077c9401c4c3b47c96ec43eca15c5588b12e88b7786d91e2335cb4f5067ea0b8a3144f2dcb93b403070762d6e1084a47bb4f6af05bf093c77ec49ccf8d1ff75da709ab4d116c324afc58ac98bdb4b8fb8895f85178870bdb8875c90d94d1a8ac46b0039de70e7e3eb38d0288c4bf0fa1554f72e9f98d755c7720dc66f3d3e0a26306c7bc8c015320024afeb7f49a7152b27f7817b96b932e21ed8bfebf5145baef07b80cd363330cff598767f5663e2df03410b85cd4d01a14f167c2c142d6fc448d6a89fb52b5be15d3eecb675694304e0781eb58285d8fd125992c7cc9abdd3280ddb800652f13acd3341218a579009a4593ee97c1d9970b4d5ccbd21b15d6963ef8e5862caf63ce060c5309e976afd95d9ade920e78a21d4781a14d13dd8851599e8efd72c3efb57347d5aa2ae0a6ea0a1b79ca9fa1a7a5a5ce59d55bce1e166aa83e0d0c2ee7652e0893f06478285dba1e672ec2f2dc9b79b28022faa040f58b9469c73b435;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h933878b246e6c8e3aec3d28dba5363672203d58820d6cab6b2155c1a0d67894fd2cb4232d637b1893420d9657f8b4186077a3a1cb9bae7d4b242c361e08eb0cdbe91eaa3ddb4492b33d335ce6a2e7d0be9231b5d2076e22cef343874a30a5f44b3e025189e3d1e5b5bda27576cc59cba80401ed923f72c02136e7d4bd97c2a9880a44dd1cd0120f3b5302a919a588e29dba569b339b4939496f35baebde8fbef0127f57395c3a1bcf5c86fd0490064279dbaba044c46d2f21b54439c2d3610fa9ffe9f5f100fa5b95c14410ad535b4e3d9f3e83eb427895e8470d29fa18002aac4199574b27c6944f3973f54a492c37b126bbefa2f7d15baf6b5d367f6d13da2236b2c7179cb3af2f32cc5611528e86ccff880bcf755d0d3319433ce10adc25b4519fb3b2cd5db9748aaff36a2a6564f874bade4c7c41bfd139ac6ef630d2d33f16723a82394ec14e4cda401ead18459f8ab7b68b363d2438d6652c65bcdbd937169da8ec53ac8a9cbf67478682f22b61e57206076078b6d622b1063004d1e59458589eec167f594777eb303d49135342dc480c316f4dc38a8e80c97e841b27ef73376f50efb3023932f847975999ba0a02728fb96570bdba2d029db4a2741fd6c9f79c973801d14952b860b17f7377233f6a22abecd1d31692cb99c76a59c0b04071c291bec432e9f3cb47f59d0e283f255a3fce03847c82db96b249c4b8852c1e40610e3a9df38f708f599626f2f155ee8dbea9e97ddd74f2c8c4485b3c0bc2df997eb8740900e5e5aa9dd1402567acd6befd46cb26e98b45cecd1da16f826956ec083bf7868574c96a4914c1f6226c4ef74824bfb6c851a44055825c532d3684cd8b06bdce8e78f041fc790477b1028880eb7e75a036fce38813d43543367b9585108cbbd979ad9303da946e480f9b98608f6474d626fba7a0591c531a435867bfd518813d374fcdbf6fdf0c3bd3029e5db2e3b41a42199c1aed1268b5c87c0635d06cb6c38c881769f7f492347dd5175eca89c8f91115fedf38a13afd29be01389013b9902bb1e9cf7cfb2b72c96ab5174cb14741dda952fc7065206f899588b6d87c2a8df1c2d8a4cf9128391859becd37523583d98ee9861538959f6549581c46eea987107b2919720afc9264a1f2c1bdf803311f39b4ad05ad5d0cba7ce285527a27a371b55cdaab2ee0b801fe5bbde111db83aa46596c1f7e0738b3595efc2bf175867b1b2493184f2a5b3fd7ed95c3a5a06d837c16e83a84be6e7ca861286dcba774a28d69a3d9f5731edd58d96e21d4cbc6252618564d99d8c74f2dc8c056e3290e69e90473e139e31a1a4b5623e16dce834d13b8c62422674e0492573a156d712bc35d138edb5b6e7a8ee7c8af7a024c3b8c6635e709d5f78554ff8faa48bc1781cba58181d4ae8fc804c417c73f2d2b8c48daa7053ecc7c96555;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7ac822830721fd3d9f32735ea5b073a88e4dc88694ce9e3d58ab2260d553e4c5ecb7c7800a1fc004b171b7921e42fff7d2bd8139f65bc974c929c9247448cab6fcc42fa10c9ac9503e1857d9ca3c0815477bcb464628eeb7e9debba2fe8b594845bc5f427ffa4166fb584844001e450909ff2e9f5a0c4b890bb7a0aa8195741d2084538a9a3d9459e101e6469bececa40c94579fb7edde8ae09cf50bbdcc0fdf92ba2c2da2f3ee8c99b1c1b719fc8f7d6336df233834122b9dddc521eb818f8b78d2da0c9ea8a1618cfcb17a2cd23deac62a8c6a8ef9d71457496c8e6ef1c0acd14520da65565d4e484a5d476da4e0bf68783974d61a91286dc7d6bfd34c02aa561bf976a253f54366a1dc7c0002aba9f2868633b258b0847bb82cbb6105fd2b8708fcb653909cc8a8560a08b9a0205ab1ace9adba5cadc0a23630eb882c76cc4becc6ba9b2405ebb02bd57e6add0b16a73eb9d0e99b9c6b4f7c62bb45727b323aa592c5435030db3ecd151e4aa0360e5e31e8fa411b8b4a1f5a5dbdf0c05a7352b1bc33ceac9e842367bea697b0bf093c036c0d9cd491f5505edc4e2163f04e73484b659672cd4d7d229981d02e620c0538f6c676997abef46d4520c751748f5c67d8adcf367021364830d7a6cff6e4e2a46e228bb701822dec81f2f40955a82ccf12ec557cb1f3c5c2bfe7f0ee15fe51373d40d341e784271dd57fe70f15b08aae12baf7cc8d9c4809d0418468268dc59d06fafacad220bd308781204f6719d4b2b1e7aeeeee2a9d2623056f920b9a9a4dda215ace68611b7e4d8abca1bed2367499dfc69f561969a2d69bffa1147561821143209da1939e53ac88d5b9ef737bdd92ea94647c7cb7453a6725ad326f05636e902f25108a1818a1642e2e170c415e622c8bfeb9252ce5241594a5219312252b0032193cb94dc8d3b00bdccc79c4d0b5027d623e1b4314ee9bafe0fb90832c77acd3279d049276d1110c0227110f918446fdbbcd7166f2a1e4953ebccc3c5989032d44f7c2df2491c6b3239c22ff0fcfb735598add455f3b7a22a3c1b0466b5599097b50132f6e2a751b5b4949f6076a9e4284c992589d56c8517603e66e4f6cd1a8ba94eef48df9c4925156fde7528f800f5cd01f8b376bcffda09fc3b71ba4f3ffb1c85a842a01ec0dd4989adf789e8329debf8cc7c10dd2e83df5be191d041ef6906b0430235846d8e4ca15e6278fa51611e3a94f4af0c118e3270803dbde6c9c84c86b0751ff683e3ed572ca2bed3fefbb97903c33043d8d2fb0e452d4f3f3c54c529b6b1407aa61ed411b0eca789f8f80922042537acbc8e82717de70235c63980727195620185d581c31da4f12ad6a210e05fedcb4f3390f3df654d361529b8287afc19f8575a655cb702c8a464e3cb64f6ca99872179876013f20ffb2766c7fb0b6b23f50ae2a2110e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3e8837ba7f97329f2785ca527cf61d0e05dfd0cbcc5b9e0f21bc20d62ca2ee6f645bba3d89a9214bdbec265b997d4a40074d2b4a1d68b59d65afdcaee3b8d2f15ea568e9e9296f06e01537c8b106487ade487da3f3a027bdc3158786aafae9662135ee68e7a039a47b7b685fa6afbfcb1ab2d4b5f7bbd156499e566b253a19901bbbcbe2e63f8874d92eaf035abe5ebd38017de9635e99823778525b745591725e7753ba03e3ea3fcc469c58b44d62e0a55eca3e45624d2e26c11804da4fac71edd7e47b8144ec75040701ec7891855e051c291771f656708dc7e80dd1b2ffc60b269c3e3417789aa035255626992a4942165094b43d4b987b17ae85a5ed2993700c9c2e60dbcda7114ba01b0dc89228676a62bc1850f9a27c86115241852df510c65542843123869351bd8c3fd206d21333db99c71dce3a94f4fc5f4743099be97c962587976131e52fd278d46f57605778ba45395aa5ad04787f8708d9fd98be03eb9b381043b811c7dd2fd110721c72f9e6f56ef4afc325bb76f653ded9e9f00721b268345fd69b951e927c9885f761a053b4f392d71fa32cd9287be55df5cde3823f8f5f6231b2a61f077d96539b906f00cd6f24d5e2f1311b73971f29cf63f3459e243427b9eb831964970c83333d195c17ec51a12b3250ca627a7d6c68b14c910d86260ca9a2018fcb3c98915a7d9aee7e0e5e3419da671e13716357d93441ba1ff1766975f728295940789d90b2421d5702c50f625d9d65a52c1c8b5ed541bddfffd6f0dbac61f45c01737117425404114de4e81c3a9f4f6c1f90ce18eecee320ddd52501535ddee1b36390b164b7516fcc043656c51701cb8eacc9be2d6a0ee122fe8389aca383ffa459d1d546fcb7c99ed21ada0e965cc675c813a5b1cef8d1fadb87f230a6ae292d618a715f9060c576aed76d88544b5f5e8563acefabde27958fb2c5d2797674fc4d631e2360d90a15b6c85cae4df09818beeb3ae4ad904ad96cf0597c371ca916de2355ed4bc895fd7379e20920b915b6665b09ad4de59c0ab17ae22f8f75c631a6f82cef5b03f4d6829ec5d10a030b23a78cafdb43d5cc9972f1e12e2035a43625f68c1b6a4659786a578574af2e7178408df129fbe58c596383a6e3ee71e86056209ed3e1c1d7ec1f9331de01f032c0cacb6d1f0a309606889aba387e3ad25a2722f26cc852c918be928d01d9e5887ab1b325a1269ac1eab09bb03a656e26cf540813c8f2be84d5b1ae780e8e94726bd5a5b9b00289679377280eb7f0b6156b11b55fe22a1427dcd53a484cfd1d912736cfc409f8e74e4e6abf9d91f01b97d46cfcce7c08d4dbe48d0c53edfa268ecca11924d725b404bb40b30ca0934712312e4e3405513707038016c2ebba0c4da64f31aa06fd7f2f2a55f34ba96c1889ed5436cd8f79fb1616c037ca9457c29b43c6d1b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h48791f5f9421641076d04c867f15e7603f77ab4854945125f4606bcc2dbaaaadf02ab27bcda19d68825f1b4ca1aab1463ad63465f113b78c5b186055651fbb8b06e51d4b55b381ef441f2d97dd9190781b951b74520d9fb2d16cb542b5f56916e06c5f4ea0412d5eee89010a95d41242ef66dd7bfbbf1c542320c7bee5ebe38ea77e31307e9e0d85ee3bee61a4ad21891537b88a45cc5d1d2a8c7a9b0224a701959fefbffdb30a98271fa0d29d70c083fb91d305465db0be39ff8c06c91e26e90ee892ce3dccbdd73a69dde8a5a34ce1b334c157b1e4e4970dddc862f92b944d3f0213393d86f8930bb6fe5cf1e5af31a1f4fd864a57f83adb01d0b85fd8a616f43a2a5be4c65d0385dbb073bf37c2a04ecf71666ec6f5c64b4719dc6fca14be588b9fa29323b6d946326992f01af0e6d70190db09e83b50714f90593bc8339af4ef0d72dc49889a6b9e58eb1fd4842c4b33ca479917c311ed48b4e9e846d9a29270b07620ff494bbf62c0d139d84cc916a07eee8e42dcf9a2769376e21b4b808eaf8184e9ae516b6e609a71ab5b566dca46c2c530a2fc8614d443ff8d5b10755e3c904e748476e95ff24b3810c347533a78e047e228d39390685599005de7b6b8dd6e06c7bf76e377277291cba0a4a003926634d2fe21f5cdc1e551bc15b98c1347629f7de9ff350597dedb6af45cb3b81e8cdc4210375cce00299b528b89eb6875c635f3d375f3f3ae49da2305a5d10e1cf73a5168523e0bac5a9fc693ed7610f2cf07a2fe0e4ca22d0486f5109fb7db7412efdcfc9251e7c70c187adc2e8f012025e30227cb9de0ed8112471bc994b331da139ceb2dedec0deb747f2a427576bffdf18565cb5a85bc22ca2db7faf255565c098c1e4e3f6b129e19570b7c67ba95b62cf2c759cd39d67d9bbac2830fa90fb234dab6f502582d491d99b2cd918d2a2da6de3b1355245ae9c41eed02ac1d4fca23fa59d34dcd84c035fbe125890c2392342b9a6b86733637ede76772f8015d17d5cf4544e7659a2026bed3d6bd91cbd61973cf8d00bd41d3965de1d36c591d31123782d0a704dfeae82aa8e12011506b603c2b834ca7b709add7c1b6362ead384d7548188c76ea44ee87f099a43ac6c736a9dbca5910375ed979bedaf6297aa634f059b5232a959284e8abc4b7615be7bcca5ac0702aa463edb6c2e8e27f63c2b55ba1a026840cdbeae8ab78f675cf74b7ebee60c060e656c3f86bc5436892e0b7459dda35dd6791f0177fb3bf77a412d41bab51eaeb0a2fed6ba97e0aa46bb083c34e334eb84f70f471d4e2c06b1e72893a072ac69e4e257d309124ee6ffa89e2d074e442151f23377e12becb9b9060b2ea14088647212a5364652f14e78806b11b075cff25e5b3b4e14e18fbfb3a2055b6836ded3f13f241a47695f2c90a553bf79215a8a3d33c055ee873b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4aba0719ba5a5e9fb9f5d97a02fceb9067549c786fe405658b852b8ccae5e8f8951cd872e4d4471f324e5f4e69fb2cd172972d0ca62a39be526f00269cfdd0159b5189612fcb141f29d7bf6356f6480665fdc2172bf258152dce27ea8d0d5a3c3b1f3c8e82e49e6fa8ddd03881d25d19b02373602a3cd214a6e14e2f31c85b2edb20e58e74f2bba088f5dac9bd863bbf37e69951921c6de272186262c539ed241b2d6e2335a8a5c121a17999d3336c4c6384ad394f088614d1e78debeef60d0bf03dd0eecaf5d2efb1da786acdef744747ec2c1a3b9e052248445535d452b0b1736397f47281a2e9bdda71d8403253bb83240b5a008c0446740529d7d21dfa141f058fe33e5486800c679618fb8bb267e2bed05b5ca85d53d1e2a957cebed53d3e924928b09badd15f7b321f3ea4359501b9801ea80f24d65ea61a5fd48ba2b62d3d6151cbdc44c095366ec1b16b458d84ee93462a38cd17182c0b076bae3eb03cca202c5c08d980a87c3393cd24c759e3cea06dd4fa295876e6af00c35c39a2196294c13203ac64564e94c6425ddec861d2cfc3a7ff76f12b01732ca6267fbdb992582047504703db1fca4077b6be6d8988d42934fa18ab37f79d762d47e1a611e1748e3440f8f97c9dc7ccbb5cac12e5611b7717c3e7a25fb3391d9893e8d0f84378a45acd1dda15c2f306538b5acca0d2bfcd68bc2dcebfa44aa5fbe844ce6310c6558d6c0d5e5ffe7a7f9fc670ffe8ef03bdb018a6d318b5386bda7a64dc61a236330e1902558d8fa5fa741ce47bba4bd63658f8fd095420829a2b6b3db2087297ab77771dfabbba40c7911abd413b8c799f36d98f0d7c1123780ace8618da4d69d69baaedf8b40d6c4f59b36e4618d4b86b8ae174f931fa61bcdc25889730d073a06b48f5153f943691408839a0c6dcab32c952ae7eefc9c1ca5ecb5ac8fb71cb8db73bd2d8896de5374430d13e25d38a3571989e90a5022301419ec6cef8acc93ac097890e2058d97651c7b05fbcee9a2caa4ddcb7037e2721d855d1e0986b32077ed7938825869f7b8db4407f857ab643c3ca2fcc218466e6801f82bd6703e2dc289361600e51975ae677d8f097aa219db45ff11964951c3eac26560ed2479faeabdcaeea15909995503db7d688482211abdf0b7fac3cb332dffa1290c10d332f1343fd1194246da12a632b96c57226b592ddfcecfe0c26da68767ba4bfbd09eff80c073b1e8c93871d00b109e0a10385feed8199779da91203bf57e7337aa3223e00b053300ef01c7603e24151f4a901b84941a3b6890d8f9ce6ab2af48db22394bae37478447b7f29b5e98ba62c3a38ae27ca507eccce3bccebfb88edabaac6b8e3a7e770459befe0986f512dce07904366b3475c05847b9b46adfe39a7c98540fe9e0d8f1962d648479980181aa8d6f80fdf66f732a4a2d35fa0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h76558c4e849a7bba516c9708c2a15af25d9de8f52f0554d7f11dba2fb511cb5143d55c5d2de0d768d9eb74c7ca0e0fd2772bec2d496d0ba63c995a73b8fd82d04b982468a8a35cb30170aa2fd5517cb10c5e98d9ee005eea6dd586285446aa87b506236d5812ebda9134e50487f85e0009c01966520e8ac0b7b15aae94fded44f796e145361986da2f3023f9999b5a9accec8cc961c1e51bcaa073d16c5e1407ee3d39bc6d38224b581eac80f13f93ada6eec42d7c9b3ea7f10d24857bb111e62cbf0fb8665279bc650bd997e736371332ffb4559332cf905cf64bc7687d1e99e422919542ae851fb7809a917932706d1486d18b52b45e7a987b148d4a6a293cb2fecf225e58406c30767809986fc55e1aa75e0c692ffb61b5fbd8396c475f4a12ef34228fef45d5b457eed7cfe5568ecac051189a582c66a19de6dd6a8093e109152f8bb5aaeacf801b236cc256b9236d6a120ee24980c37cbb96c6dbf9f7c314bb1a629f10325cd57a69a47c2b8468cb120ccfc17976ade505d8e033c4839c2aec4b93fa3c68003275cd79aaa3623f9a8965723c02ff897f53480693d7f3fa2e717adac6b6f3611695f5b67b6b9cc6bafda0229e85decff15e94289a4e87a3321975eed1037ef4b28b560c9a094ec3113d9772dadf46046bf3903b7bf8da3982cf646be828a48c3ec45b48288a929a1cd4b92332ba2e9a8db4246450081926e06ef9a70d00a4624b4bdc18647deaac749623cb3f4fb2323a454365a408aee5f6575196b10f1530a73df2616bb9319570050d1196cf21ef6e5d32eb672990663304ad9be2d82bafda9708f3692b415afdb1fd75551d68213a08d56a4dac0b88afea365b8d221771ed029f9c669ab955fe651360b5553fc264ded2ddbde25c6a608b8843964744ecfa6f70bd40b53f00c5ab6c784ea59a1dc0b9fc84cb490e2f7d64e340f6f6f5a7a1f711e00604ba82885d7144aa9161a7595d2cacb56e11248d11a5da5ee377800b7f884b15e22f9f8e6c01135dfbad82d34b60311a0b19e137a632273106f9c16d605055549001b91af4121e0460afc8a13362b987095f97d1acec789f9cd284ae9a6fd0c71f985f96e4328d4bbab1ccb13858835cf57dfcc80350d3c3d09cb5f0b6cf9ca38f05f575fb96e7d1ee8e060775b00e4c4751177859fd831cb6c88b32529f28511521b67e26929e2b3a4fdd346f385305cf506cdfa47293e9b375b742bbefc943c67b89b86e567ee44b135cd00f10fbfe1a43804755da956de858262aed81723e1d3873cdfee1ae3cb30ac0b2dd3eab0404907f3581fa436c930ba60a28752c9919a75977a3615290425bf127cd60ac736e897b174e1e8262c20d40fa14a81b79b5a8257d6e648f46c633c86f9551a139618d073b74ff2491379e082dcdecf0a560bab317872ab8647c6681e4466f2cb12b6f4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha5e43078992dfe22abf3574dc04e0569f0107c6585cb09508285388a9e0cbe84fce6b6783950c64686723ca9811cd58e0953ec1b79394e4c342bef6a055fd1a33c049161ef069788ed6eab05be64c76d456d81f92a7ee2be560ce18c8216f671d3dfcc821447876377a9429afeecc8189c0f43b3f2759aeb8e0955d4b032fe20af836cc3d2998f8763c53dde2f18664db0d5e2a5fca258b96934c67bb87c76a26fe01a065b7b42ecb5400a5e5ee9d588bcb68da93a7c95c391cc62dfceedd80c156a23877fed2c2c7239fc942dd1c936ff29a63e7f4c9ab58299717118a97c16e9c2792e68ee6ef2a8493637569985755dba857ae8d3452a9b1f5f4c296b02dcb8bcd18e4ec5fc3e598bc83dd6541ff7e5ac77179b7906fff13f8894761606fa426575a5dfe79b4fb61fd9bba3df403c0f3b1f881b781178fe560a134859ad0ca1b86c3d378e010f271b648f0fe0cfe512b86fbf9821bdf01280400d25b12b195c4c4ebf6cef44b4c9ce79a91a2bddaad122f3003962e8cf0158c9f64cf9d71c8fd2504d445667afdd3a1bfdca9fc37f2773241d41cf12406a479c57032f4e9d2ca5e540b15fef92433eb2ae7a8ee62de17356be337b5c7d77b16bf59bae2e3387ee112add00eeb1cd51fe775c9c7ba7692d68f3ae964a568813e76f73e654d13da17bdc94ae1b226efd213a1f076e1152fe40f4c3457978747ae600547e0bcf612ce7f5756c8dcc1bec60eb7ea0f79709ed5b129dc33be73ebf7782d81826113dbac277d8c471d3ee51af013baa8136bd436907eaed394268d6171b3b433fa44590e0c73db177dcee732f0a8ebd91e9129ddd782f0db8b908a7e6d6d1b1ea1fd8be57e0cf898c947bbfc4be47a7fffd3f82517e64af8a8887a13ed5685938718e79028f1e48d757594840eb6f036c097b218001b4ba8b7a77ddf619ce871ecbd93eec19d89ef0a8e4f51cd7813d4f3c5f86fa07ebf1098131ef4cc7c6a1878083f34e5acdb4df7e7eb564ac1631e3bc069f30df6f2f9adedbffec6df565e7e4a87017e61f7585979e12868ff6c0ba85f09705e476c8fe42a44a2f0a44d0595e051bcf8359c502b381a417dac4237dbce4207fb6cebd8d41aea529a45bf4ece0d51f24b42c5c0df0f5a3f92361cd956c688ccac31eb09937bf582673d992d8c84065d44197f8df02590446f42db537dc5a59627df1d560ed0fa2ec33f7bd4f114d0c777c48da9efd63a525628f3554dc74e56767a880af93257744a7ecf4098fc399cb6e1641bdcebe6669ea2542602f48ea76e523e7bc99d5c731f6d93efe74566da96e5c8b8b69c838da9e32e2e429c1622ce99b409d0f18df6592281c8a8bc2f083cbb0f0ae0057529fabebd4b88ff75b27125efe1d3abcdeca1ded85b0d22b8ee06ea3f1bca36da6eb6a2efa757b4fdd9f3619ec4338f79289cf245e8dde;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4f409b0bde88603d9292184d8500c9899a97d8e18e09ed98680d99f1946a8331fb6f387a8765e62cf2f8aafa1f5323c35b58a917a31ecdd5eb48d143de0687cf78fdf20d7d477be97e41cd63f9c9a432dc716a4704dd16e6f21f3cfeb433125df687745f4450154d2f17dcdbc07365b75bea434328277854118b64efd889da0e6ae3ff956e27b4bbf8eb0f6fafff0eeeb00f02c3fd8e96cc9bf96880b37794de52f4a823de2599d7a1afc018d141c4415bf0da551fb9ed951691342704502eaac922e8782f1f5007bff37fa47140d5e37c8fa7fd822f205761d27e0f33ccce813ec3f579dc6a775e4cc18ebddcbfeb2eeb0ebe54697e74fcf36ff9225cf3cba4184dbaf780e1666ffc70f232b7347c2601bccb46beec1dc17ca1efca23ce928ea8edcec1a4b91fe903aeff5b55953d5eefcc165ccd4dbb24bc156096e9f69939daa5586fac25df1bfe4831f14610289ba86fec0ef8a5c54731d4e60afd6df9f30ed64e64a88ef0c1c7a3cc9d14c95e7c2eb98846ee4dfa36828226fd7291410983949a9ddb5cc71e5ce51f5ef41c272e0e33c196087a7308d077973092e23cd71bc989c28a7a6be3f1c1032339afefc31b96ed1dce3845a24f0a6f2cbba1522a26aa880fcb4e7b58f5e5de4ca3328668c76f038264df25f0863616a9bf01986a084cd61704be0871f0ac4bdca1290ed066ae875a1a3ae8c8f45975a74028a4ef7e27bd03fb53885b713308d4011a699f655a5a832649c92e63935f071d8b3fd49c4b6da6547f58a64d089a49447840ad230deafc957c5fb527d52b62f17a618a354ed0deab9cffe838a3a8f1fb2d14c04c586e39fead0d5bda430b0dd91d4696447576d930ec890440036ae948552d9ba702edb57157a1fbb9662d43be1b8b64eba642bb20e37db251a7572fc1b0fc478480f1b7a870380e6886c2cc32ddd9fe0508913e7c79ac5046fad5ef3b67b781e34eb8f921624b19133e9d7728cc6157d115c3fc846eae2de9af79e282fae7d99dd71da52b278bf1e462fbd905b9103e04dc25de35f98bc5f228f43369d1598e8cc72003571ccc343d1d2b25afa78ed344f05e6c673e21b4ed45c1ccd8d552825b949e9450069bf2fe9b164728393f0006ed3a481ab162e7997323973a3f7b7327bd876995eb123aa29c1a3985aeedb579928ef227290f4135afea29eb7aefd784778742d3b850b676e407f842713e0090c36e3c92c699b0b075bf8b1f79fa0b78b1d9aa6785fe301f8d44cc1a1edbb63da7d9827eeaf667c12a8aa8686d154b04d77b1396c21cb563d3583f97333ca7f696e37f1b480226f3713ec63163f231b50b2813342c82d8482dc073563fc4b08f81145df52528c4a32d9b8a943b79e1b169dff0a904b3cc3972dab3eadbfa1306e585fc2669d9aaf7dcc5868af04fa2abf46dd654e3de5572e218625f7af3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8a035b90a450c3c3ccc9b4bcf772cd2f3ac5726f55b8779e03440125ca0b4b7d1b8b422a9b360e7fe48fe45416eb4f4f3847d8d556d55eef5e5f33dad114615b80229669f01608ecd52c82aef0b77013cce6aac4e4a5ce9e64b6d1448b0afe98735004bb356720119fa3266e5cefa59d8d46722b851af989c11261d649cf3aaf07a408bdcb900d7996269e46ebad8f3ff1ed63b34f89f47cf9ca1e913261cb6ea6506ac0316fff80218db3be5aa37184622a6816a2580875248ad8d03cf9bb50603c55f02d2a800146e231c3cd8a1c9b62788e513f192f4cf568a558b4b1ee56be02c8909313d9274a09de576400e1ec934cbb07dff7155db0a0dbe53cc7a1f0a69b71b74e72868af10de6e34be5a1339b0c445fb8838de19d005c7a08027179eaf8051d1dd88260b163fd7a6721a20a3c44c3a582b3067c344dcc39b742d6a6373178d1cb757f98b2d66e8ff81977d4bb07a0d4830a262746a32caaf7b1c2de071fbcaacd0cb60231da388526116153253299d2505c4dc56b2c4e55357479632256026d54ee7ac025192140c22ab7eca2bf83c49522b409668ded686d6f0c21ec2871333ed8350261c7a980bb280a821466fcf700b4826b897ce45e988896d1cb851b172ef45966cc7436925d79fc9be23ed7a831c8ffaf71025bbbae81ce30a2849dbad264e59bb2dd0bdf338854c238362a52d4971db5920d1a8cc82453c50b53c0e56a0188239bc6558ef2044eeb5c86e36fe266aeecf501243bc80617613911556b70ef3a2753164d4be176abde11cc69f997e483fb13c04b30bde649981d5eacdc7d79b37e3f80900c7bf64a9aa43cc519bead1de4bbaf238452f882318664bad701da2f26ba54cc5e2a46bc588b779a1e6951f3a160abc621027a42dc423d4b31011173dd5159d924f76878958a4bb0ce7cd530390cc692a0c16d7b134d8389bf5292588020663ed1e56eb8fd590aa172ad1db7991f107255a6b95e89c47527601992fbd90330d84a5b0709bf079dafb1b284002804b58d5e5272f23ed8274bd4172feed5b81e24b3aee2ec300f171371a722f9d3c897159b4c0c5bad40647122aa60f361c5209d6e4a8aad386ff4442d601c169a728fa0f51ded5b75a20a18bd285ce1b66ca18144836e0ec288af964e5d526a37f325cafa84c64306918f14bb03dba44aa4914abbcdd7399c4e8659d274ef30ccb3b3e3fd9bec8a256bb75d57009fbd081f6738f455bb452ec2d0c4bd7d87b5d37fbfb56a3b64b3450e125c39be2d4f11bd891130ae24689e30e43ada7255ad8c3900a1536705f77840385f9ca5fe2ee883f48bbff582576a56b516f23278b484262f10d783b17254b28c571bc0b849cb46f7ac974bac8517e95fd2805200854506ae9844d21c8ec6d65658f7f4c82dbe9d747085915777af18236bb1cd7b7e3ae9fb3e6c99536314;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4680dd2d60d5d66373ad2784d69ce2b0a2f43c15b3d6e579d69a0bbd60e89dfe2606069c33a94d63a950d31a720808fc17227a0fd812220aad93f18d462a47dd7a4e6083f03777fdb47f62c27d842bd0e11d1cbdde6a7b41ac2ac867a3e4f88a6d14fc2d1af921c149492d31952ecc9078cadb166102cab25d56268557ea7b6a3c98105e615d612c7f31d250327fa3711fabf6be97d41a2e75a95082eeca08c008c7bf16ada5c48c77261b27d94e7adb99060a589e13acf03a60a4075d96d0242aa1db17419d83dfaaf728655a694749dad702a5c730aa4cd089a72da7257d26cc4943241ef58e1b4ea6f769c3beb3d4be9918a000a99c4847c52d7b9e6d4ba4a987fbb75daa1dfe13aeacad3d7af4a9328438a770dbce2e3c48c74476b6ce5fabc67af7274d024e74cf204601c1c4979e24e61bffc712a17f316880175333a104021e97cd60957b4fcd5aa8f2f95aea8c1c767cef37f49bd9e9ea61c116924c39cefeadca74cdf3ba66995f059bfb0771f64e336683848a781e4ed7420ce4287d10936f6eb3f6964c915fa56a7cc8507bda6d47481a220d7a532ab4b5864ea20c220765f97a71d237eb825b949d1291d5996e116d226e0ce7ddd1ea74cc4d64d2418d263452b5ef94252ec67bc005c9d9fec64720a30aa88aa18b89a0b92bbc3a226b71e27cd820b0f77f87b86695f664205234795f5c14e614c01a594b196a4ee05c8fbd527eb6acf8542574705f830c6ac9a338e397490b19c6313cdac5c4b9fe7a5de59938d1d3c9c1504cbe46b44e8d161f27aa9f7f96a0b4911836d3da03301e0bf70fd69839e097d49a108f9e6a90dff5cb825a0c90b799711b8a163ca3145aaba73410d049aa78cc5e3480520598d6115f85108fa419fb8c89ffda6388ba7ebbbba1d2f552e4c7c2cb287fa894d2e4820d80fc654e97428619ffdec23914f484821b021cc0d9c0fc56f61abedfbda0becd4474514fcf2416c5ba29e0069ad1068a47563c940050354dbe0b62e74741d0041c4ab3c00b1c4e9d1e0cf04002ba7a3d092956cdfe0d3757a859a893da36dee4672209c6da8bb6c1df3e27b82bcde0b4fb8150d2d4f1c977c2ca54cc1439b1505add3d5b35fd518a828f667869727d7d12b65057e9e15fc740a7b0193e506bb362121fc82fd43ac0b6b7a90dd4cdddba0581bb02392f1b4808b33160b65b8c8b4154ca36bdc1ccce615156da4da8505986aacf62843d507af1ef915965a902aa0f57fb0d4700214830893249b761d6870a3a24d06f8a448bb3bec2a74ba4c46fad643dc3290ea6d765c9954b1a4d040b3d9876291491d23368fa2022d436016e83a16ff5a1c21223f78a720be3080bd9da1dc66273bc6d8eb3edf4306af92dced3e8c63c89f6cb4455f47e714c14f70170c2841f5ebc03079a90f44a27c58b4ac267637de532f522af8ec8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h99c6ef7d213e16e0ac109c95da3cc457ad16faf0a5ece7270a6d830db0bdca68bda372e97e0352e5a7c8f733f75b207e8d630561540a745f62e0be34448a69f9c8705367f1a96314ad6a73e806eb778232101a0adc0f39dfc9f751e7b4bd92c660da1a2ea26e977c126335c5a4ad4bf60a19509ec1f8366aaa41794b20cf61e8d95affec7b0bea97cf4884661351103b1f9a4b887535a0e6898e55c8fff49465a616da901d5b99b50d713894245abfdbf353403fa0d38465a4a2bb94e18480e502f8326b1cee7a05192b6445faa8c2b945292eeffb3171b10f549ccaad0f7ee9e111d4220645415899fd8c28281d0df72ced562368e408342ed4ef804b5e5607754a307a560a5838cf6f36c94a702c2026af0e1507eed20b261809e295dd682f8f8e9aabf8a77d8b2ff6da50c9357cb5dd670d661e6972b25c8c1d4648a3c8ebe6c88fbcdc686ff34b29ef10ec9dc36c6308411b54c253900157fe11479bba5587155c1fdfecb09439f42be073eca23bfaa57425390813c06e2a8a49efd0ede2e51225485be64643995c209d48566fe5e6ca0e471924b0445b4897eeb62cf35e84923eef68ab88bb77f50a75cf107ae51fcecb0f950f2a05c8450047790a4baa0be7406769fe217f7b74966e333afe2eae69f3f6d820985d6382ccce19b38f92c715618505e7cb931c8b75b1a8206096987f37d78836dad0b92299f096953b3667fcf9a4164e978c60115220fdec07fc33f3b01a8feb40ae9bd62a7568325e96dbdb558fa2c4935e4c0fbbb610ae4b9247169691f88d0d2394c614d890731d91a163360dccd1de5985ceada6dc0014c348a996ca25c66a483b1fc97935865c2e826d2d876a01795e48b724eb023a76bb9ee6990b4c2624e88040fc5c6990f3bc6b5abfaff0448fa331dc65a8603cee71f52f4f851079ccd8a4617f88b28a53c3de35d39155b9f6eea3747115424629e009c473f6330f1fb0068f2b6ed2a92f226b08221a2ad10b4010625849504d08d847f5284278fa8127e55b92569f68646476e97db12a22de5103020a4ffaf0a7a967bb6a879d03a73895e4240be9693cd152c30fcce0fba8a4d0cc34b5fe0ad679ef69c48fe598d4be0bb1d4d06ce7a75686335ea86c9571aab063f7c8ea68c0a7ee7a3bf3d77e5e295016e2c638443fca8d2eb9dd6dfdba229c0e75a41af58a2984c885367455ece07a8e7189feabb0db36c2f2ffff69f238599ba01aa97da1fadcccda2201c1dc62fef5a90f34310c03226e53f41eb8a22b0cd574ddac04c211433ff1d4fda490049f49b361287873634cd505dade6cbbc92f3256a009535ac3ac1b6ac1b3974cc8ef42268850edcfe3fbeaa9e9a4d7052629d2935361318c80d4b7157b97e02c0bf915e04c5472b38152299c0e644705952e735e621eeb78b62d550179e0fc461264473b5b99963fa7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffd20a7f56b850db5ec376cfcfb33dc0dd189d90e189e16bc8f611d3b4d61e2880a196dac39da48266b216d6a9f68d46fb01ff7c0b60fc2650aef682d7b5e102e39370e05d32450787910eb5d63eb40965c06c31b9700e4197f6b68876d6ade788e910a75927f7615236e67742f87a5e446b2195614610756e549c97809b34a0239651289ee4b0853a3249e0738f0bdacd691df3c3cda276b2b6910a175201666176766ffbe7901fbc036b97c9ad01287932d21aa25b6a19d311b9bb3360514dda99a3748fcf8e9c0ed48441813235865b1af5d4b47630d7504495bfae7409d38e26cf7018843657088b1de8e5e50266232eeb431eddaa22046a4d30cdcb9c75c614ff2bebf36e25dd6ada6511733ae8dd0f527c30d84dd3a5e6646becada97b5598257cd8dee25d20b49b30dd88c3af83aa21925a6a5b18da39488851f26a75fe750c21685b63f94143fe48a44d5339352248e577d58e8a88c4f0da26b521cbc1b38186b71a75a5513815af91fea69ab9ca340ede56e5c071e19812432c2aa90e73ff07a1b46b7ea852a2842526488947996a5b9313d3bd98a263399a91444d0a0c83c984a1bbd166c0a6fe15e469f73480972555747a002f2b2cdffcb859bcbcd66931805dd48f801444a3d6a40bca1b24fbff4232bbeb7d0689cb896cf461419e44ea5e734cfb8bc196b1d4b8105bc705c8395899db7184638322f7a8f8643027b023a7b63aac450413d45c7872cc8d431488f0c1e61848838766e3972d4749a0f08990ad41e6b2b7d25872c26d89bc9672f6d3e7c54b36c139196c8c678f9e0268108691c6f54f10e592d946ad34657cc414c7b3c723b2c02731485024a947669627e790ab88e1b68636ebe7024fdd760e6284c8761f74922f278e2e3fb05f9a8eb7befb0b8d42401d407e411196105306b24cc64f03d8ea6225e83714c9c3e90dc760ceddc30ed2b931b43bd1bcaa7c4fbc453c6f313d170eae8bb207e7ee12338bcccc1f4cbc42851a3c9f065f959053095a5ac021f8d0da92c987933de791966dff2261ee59d7f4f4ed36463f7d57a8595c2f876f579b61a56a00509d98ee530932008ca2a47353ea3c9ca5ad26ded293c097e8214736f30cdbf7acab58c38ea2194d914615f5e4e7caa3f656349ad9b0df77e610978e6fade33fe47fd17eac1b379f7725dce145a6383565c772deb59c36fd7125e6ba48659ccc97b918408b40d2b5f56ddc7fe021d4687afa9a8c133cacdf2cf0971ab5b1b0d989b2ea127e204bf80fdc9b2480bbe1010ea15d400bc7f779db1c58a59cca116df30d1875978d6974ad8aadd1ed5fef8eef7be3a5cf1b52b4a2a855640a429cafee2b8fd9608186d9c3d0733a30c51c88f341c4a081f6622a691b25accc00bc12368ae0fc6179256387aed463b7f0d51e36396ae9089bdb5c17a94899b53a304238a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2b910cf5e347677be5c11534226dd6b3b824746dfb6b3522498e9c1a4965c036adb4d9ba08b221c4e3eac50fc3cc75427cc5e4c54b4d0b17ca1f5bf4b0dbef3eb62e6f30656cc367c6c196732abd72887fb07816c943cb40bd7a356b6e607c0fc6d8478916b7bfa811e1de91b87a0b2fe73e141a1e290ccbdce65915aa874580c8efb7a1aa27062ed939a19194cd645ae9a5487084ffdc48abf60ee1e57376c8acaa6ae5db504da380c3408d83cce0f0f926a9516a95679b110bf34abdb9de5fea78f68797705e1836a3c8e6f6cc0d10790650f58e65b8bd48704760e3b3f0b84d572a37bac802c6388c6ea484981edd19299553e51e90e823f6991a35c7a44ef796316d8a07abd32846a59373544c6a1bd1d548aaa2bef9e124f32f8c52c5fb147c536f5faeb46c575f43e9eb6835ccf94ef734661e4ef268ff326f7350e7b18465404c8101a460be91df5242ddef1f07dc18661280853cae2e4837dd7d944322dddbf033f0a349218c41a22dc0658f930952fb8b3d78d34aca3906444660dfeb46eae44c0bd5f8dd82438fe59b3e3f1a0c51a98219e1da2091796a7f29f1b5148ee8c51dd469346f17d1d666b152f6e1ffd1002f2f99807435c38c867223a29a8b991c054100f55d5f428b1d86741190c3958e63fe8ed6fa384e57a6bbda188b85511a263d798a29951dbb7fa1ac073f483e70bffc99608ffb4fab63b9e4900cef2695375505faf9e14c329eb9fb5653d54c87dcbe293ffdab10a6c62e055a9137687c7e8bf408c60d38725a5b6fd2185d7384aaa9cfcd6ff9b4aaaa8faad6c602a8dea05f0b871d6658bfed1faf005056a719f08739c5ef9a70e30ff6c0bfbadfbf6ccf796485a366746aed39e1b3439f8914f72a27b63ed9ccbcc03610d11a21bb41b967db2c712259d6eeed1c7709f7db46198334b474642a68a4db2eae825121efc572f20b2281803ec42c924469bffe831f787d4162a6bad754fa564199087d1853205cee73b7e9c262220e6ad234e218d9ef1ae588d793119dcef3e1083756a8d2a04f42b34166faeab3890420a3f3a88b49e958858f809fd7c08eaceb1b91a3c70908e5af089873e21719f5252c84370f975e3e2a22723b42fc8f86e9f2832235a42b25e63ea3aacbcc5b91e07b030fee377bebc80c0fae9d6921944d2a53ccdef416830bdf2bc0e651f94bbaf7948f406cfb1acf758f14aab2939d86eaf82d93454c5b225aa6a8ffd75d3d8b698f740b2c54cec11bb1abdbbc2db16f800480a62fa4dcc083d7769183d48c53ac79e4eff9959c1f1915393a61556874d85149b26ae334f282061439eb93e7f162bc7b70b8fae9193e1cccf0e4fcd2e498cffed5c330fb7903af4a7ff7d8a5a827818de3d38ca3de9e89123aaf58da71285887285ceaf83a92e3ec8349887611261e5216086d0eb7d082949f7a762c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0c5de3ca622b3f2f798d4169e303e9f6d231aa8e28b6c494487201599a5f4390f9f5f7b63c187fd5511a7419c3a183a4dfbcfa8dbc8585e18e54dd0aef065d3b8e309864e10bb48dfa89e8a03d88fe71579e982e61238a8fc41ba3ca64702b69e968d2d4243afaad9b727266b4d05efb05342a8fd78bd2239745c902b6dfa11f7f685e0cab2abd9c1497d6017cc4dc3867dfd47be909360033313a069f1f2b883ea37a87b8e1ed2a95712f6442b36b1f4f60478c5f69998b7bd0bc6ce974d8fe7acdcfe64bb8d81fd717a7b8930e3b478d3bad8dee9f78c2cb3fb901c6715cf7154e42557ca3f0c07968a52795d33819305541566652abadf3c608cd2514262506f743234a69475fb33ebd9372dd57b2050d2be67b003fda3f464c77e0eb3cb43a4c386e5e5a2a9bb403c669bc81901c1d634a7f255e9ed54aa6e43ede50f72171511b9f75652de5e01597a51592c229318392b18f29bda08434eb70b1c0a21f0eb64f6a293767fec3570bff63ea9a05c65283445712c2e61951e5ba81039d443fbd39319dfb726eec82a569abeefdcba0168077b4f64f32d049854e5ac73f0edd022cebdc54842fb788f7cd118719b123a6977430598f2ede4d0957222c7a7b980d9fc7f3a40d435a9a7399fbf7868fc901a89d18bd8c7c67561ea1c37a3334878983ea1474e56425d1dcca613df50a5a2d9bed1c68e6aa49a6216e402adca8176fbb9c4e08865587e30fcefb826c999136af0cc6eeba1723566d31446d3f634bebbb4769099c2c90db67bf30ad3aa51cce54027dbf2bc9ac9c533a22d887ef82bf3a010e7e1c78356a7378e030a52aad1c60f00ec7b9bafd42968df4956f75997744e58f348179dcfa95a3f7b10569fccc12c8d84df53ca8d22333253d70a17a3caf7226ebd45d6035f4a6d09a7c9e4a4fd9a3333f196ed5e04d75049a6dcadac25160a927eb2b007027734e94f6fd4d9d8e39de360fdc9983c98bdefcbbde912453f3c470c57e1d438b992f9ea0fa5685a52750c2ee73c6719440153ed1ddb0c76cdfd6d5aca7e39db5fc15a89015a5df18691f0818e3b90d1a2ccef1e3bf36ec664002f15c38e64c541707024a75a8a34989c6c38d9db64f52b748d76b2d79ed4134462421dd5cb88677a8c1062739e39df3693a47970460a016cff642eebeef6f2cbad6c5f48f740b8e950b1f9c9fc7ea56f038bd850d1380525fa1f04a02a4293954d37f79173517cba7b766141e019c4f1255dc4dfd9a80f24f5a1087a77d7bec573a3fca679213c57e7645323b5b114bf3f04bfff5dd18fb701f26c137f9eae6b8f0c2690d71037c97d42b0f1051dc06b441a00384c1a21359ed08b8818a6caae3bdad46e74d50eedc88fa72b52aaccbda25006a8b6a6e097ad659e53bd11c92619cac3815ae49da2c4672d88eb0623e31b1e950d8d756f9a3cab95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h65d3d83c48de233319d929073ecccf651e07c0e274c6df7aa4461d661386bcbb6bfc829e8c1c7e77ea06871fa87196bb89bafdcc57fef5efe617adbad8a1a0fe1169f460b04e2e28f4596f2b8c583adc92c3d4579bd74f78d14c5a9222a4d8eacd7592a3815162d1a9321eaaa6cb643852fab6b43e0ad6526a49d3cac55c728caaf4c668b7a216e89ecd49f132345ba44d85cf1ce20b96e239583e396fd5c067aaa357eb7a0a6055a93950ecdf1255b0ace0a4fa78ede2d99b48333761a5b33ac0ca07d93ae86cb98fcafe155d430d9fc65edab885f1f21a4208e49af83cbaa1d57a038667b76bb4c76291c3721cc17824eb3b7eb2270711492e71cb20ac28a6f1863f60325060a3ff95f5f6bc565920d0933117ab354ba0924491a65b50aae705ee77dd869258e2a31fb674e85cd6a3b2994cac40a0651ac14b03f2509ce9649da639a7d98ddc34308e9748eebafadb02dbdd29514e085f8b2655e495a740ecdffb9f5356e70a1cd72f20f25a4b5d6c5232bfd0369aa23d4df929da2c4cb1646e77117c3f92d87c61b7e811ae051a45d89803dd55a4fc9513f7cd4659a3830b02640da6f6a0b3d584ec21f28aa74f9e1d8621cbdbd689a5a34312bf9fe7a777e0d1c155fd87bb435464a1644459ad2f86cf9516c9fada9696403def73d1785339a25795c1c099f3562292783580da61c8277502bbaa105299e0b6227d87785f5273bc5bb824808b0d899dbc7ae6a05480ca9deb3642940e5cfcb4cf9030d3fd1427ae55335e30e1c120bb543e249484f6e00c895fcf72757b0fab1be8f177aaed1d81d276b1b431ef029a86f98b7cca386ca8db6606008626969bedf2ad8dc24cd2ed3e36de8997b4736ebcfd48386f1fc994e4aa71dbfc7faa9bcdd7a3af70fcbde217d57bd834c2ef92aba0b8ca507031aa0f7cf10ac8dfcd697efff5b760309d68d6fa30d29d5c72997052a39f4b3e027cb2ce73b70f5844d91662d97f319b5d4148dbdd7f43d263e705cb2ee1aef59392427c35c973bd881f9cefa9cc833b22a7b12e669786c21ec479e18c4d75d109eedfd0dd674c8c0f095ada63212b792ceac053ffff9e76b2257326c2d88313bfce4df2c6a87b94ac5b842ebcc18799416f27c50a821046c2d8ff30593a681ef02da58251f3cd3bf53498422a4fc6fb3387c2125a049a2a3665b730a8fd530ee868710df06d7f82caaa9534a75d96871d0a9c3d25837389762c771aad86f4fe03ec9da02d8efa7e36017a33e5429b36da8ace2e6e33b40732864e7e6f4c99fac2d47116c898403ac85adc7d79785c17858f2f3bc2d0c86cd02d88cdb838605b6ba45a87befdbfd147bf7e5c6d6cf144285c9dd0fc28e2e1e1883e78ee9f447d6b7499cb186c3b237bd977161a64355fe77709abb6c027bfc25c96c4565c24b41627ef22175c925c6c90bc2e18694b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h93d88ec7614c823c3da47ce4bb93765be346edd800fb8eb1aeaa4f3d78ddc8ef6ae048899f90d954c165dc1c5c54659b960cd357158e3e2fd5b2f82be5f5b2c2835083251ba1c2710e488139fea69bb2d999e7d75eec8e5974039a3a184777886cf7b88cfb8d391f21c9f14b2db57052668e9425de74b4be4e82bc1ff21af3e2c0464e85ae54f31dd4f1533391d9d0860a4a3e91fafc7723558a780121045953327a19cb78b524c2d50b23d5ec3d431fbc6a406a4b0b6a5b136fa4604700515a7e6c3f45594743183f00ed64c05d15c452f3c3db948fa8e61f28dee7fa4d797d9dd1744ac3de260b078caf6cf77f48e461d65ed1b5798627103eb6e157d090d97861c6b6217932c354a7c36578f2bba8576226bacd4913673ee42dae0b139dbafc7ff7df3e1164f41380b599041859ad9a8684a1398b92e6f3010c3c4a13454c1e072764c8625e1eb130f8c4731a7e59baff9ed82dbd6b0b1cff7b2f5bb5ed99d0b8e67b7971d8b210af52869bc963c9ca37562f61303cebf742a608c55e36f9443c75b34a8700bf3f0148032bfbc29c04d2ea07fcce7b56c24d372cfe92749cbb11c024d07e8fb944eabdb6e53349fbaff96f9734fd4c59f3b6dfdd95c0dfb554529a559d64d316db661c68c734c98b783a554168a6df477e54afee76ebe36bbc6cd9a74672e67624207a93faadc682329e512fc42f3051779e1f4ad3f66e94e700f8b182b4d8e36f11d8ca1e12bcde827ecfe9c379a05f05b54a5f5a3f07dfc07dbf0dcfaad00decb4b4befc86fc1ff7cbd3461a801874c9cb2addebd1a6b855dffb80a708170db66a331879dd03125991dc7bb401731a436e3a8e61d83e8b65feb452c7ac12a2f8744b319360c6f8bedc5d4efb5802e2ab6c1e560586ee575f2ba9b585fa1c7d45585c4d603d0dacf6c32c3ecd3ce4a8623d72ac4fd40ebbac436a4824c833a64d53cd7a51bab39cdb4a7d322c32c340b187403e5e0e6603c537f0f33be7a02b02660201ad7010d90908236225e07e859d4564105e1b65bd4285577ddbf61dae3bc2ef56da9411735dcbf1e7eea77dcfc1f82d87b7400cf5de32692ac23cbe1ae352b3dcc2f8a5ab85665408a70b3b05906b88e89b1bdf0bcb0d6638df73d98450d5fcfbf08c6ef188d312c4af297c24e3cac4d10eeb18dd36666820404e30ea4e44675ed4da8537996efe1ea8f2fba7fe97a5e788b9559e361bae1c2158b966b9fcb06cd8de61084dcf7c0c2473c0f390c75e0a523ff8d39b6dbb6f58be972f971725e9e3f64ff9128571307e469a2a4d327c4b7aa5ac1ca2b7208e5e42ebd7941076e8c2b37425b0ffa9bb07ad7a53f554795f063895c9c6d34bd1aa0a242114dd1393308fced36d85dd21184bef437dfb19b25f606a93a2eb3206c46c0ad6ff7163cd074445576310c20b45cdcb34d7b6de64d9e95ab0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd3a4bef48b383c7b32cf9988fe0676aaa7b24a87870dad3d45d862bb3c71ec5244d3743801c1fe35ad5f748acb5f69996dd85ac12889dff02d24c0705e67b2c8614786c376b455be77d9e785279309b2b33464300b750e0f8104c86722c8fe7f10bddabe8d4677d2a197bc38f24cc24293eef06aaaee7c41422a4218c6b7bdfce643457775efcb5692f3eaceb01300b577dcdc4a71321ac5a4f2f56e9f45cf1c4d01a42075975c8db938058bfd8579d8b89bcf7508d0ccaabbc8194daeec5071744b0cdeba4f2daf976ac26188cdcbc4b8617353cc015024e2cdd2cb2a6c3d51ef5f96787666ee8394841e1da8e9512a31f763c49235e7bef971f4fa2c577fa12703b04fa1bacd93cdadba9707cb422add2c07c0077a55cff27af89789db4040e9195f8944969e43883866aaec88e179b0513b48aed3401053840dae1831f061764f49792b428ff69d96e01541170d1d188f47940af913aca2b63d5617a08b0072d9ab83221da3caae851d1b1f9d6afe71ab9c8ec5c3689c79bf8938b30f97bb6871d826c9cb2cd28780b089c5b2405e94b99d27814de9cee2c71289bb398d151cf2b8695ca2fe091e49f4208e929d313453f96bd753c4ff9fe62c5b086a50fa428ad34d4c87288127039ba58c88a22e0bfde10257a3044a41cecdf9a6eadc75d1ce3a2dbe4a9df37dc5fbe3b3a041f8702d85c57a750819c66fc363f08bb8167a5ec8891db644b7732c3ec069f278a0dc88cc3957e763dd4886f418279f5861c22e62cbb886d8619aa2a1a4262fc3098f2efa37574ce86d5ce180f1aed24df389bcbdaf11e67d4f1953bdaa345c317486cd0f7ea521a2b05a54d5a8ad6c2d46ef1a7f440c7f7dbb4828449932adf230552ecff6d1a970ccc3e7748b44daab526aaef0fc2f3fad8941299fb043bb7d954c83a10fbf6398d9cb33ce2e5705f2cfaca75d9665d39ca52cfe4449ee2919f82313496c38eb5e8f713f2b52b93902e5209f3b530b216bfcbabc619670fed7b6bb288ed8a66eea68c90c5aea7a208ff9662c5d539f4da241ea9ad6961872e1d8e0d875e9c9eada64c0b56451a91ce4ef064b8e0fb618b4b52a6da5f90f8f97e692801ac0b214ae97575c6101cb99c7584c4dd14714a7c48e57805c8e9fd4a6061dae55048d9e657daf1ed1461c0a02a403d68b3e3e5dc05a1aa6336b3da1d2b2e55352ff220177edcceb7f0f75969d582786b737a05fa48504359660e0417569cc246e847dc413f65532ebf2ec2c7c58bf7e28ba17b75fe53da8c1beda1c90e08f5f00faab34d3d45702be42af610354e218ad60caaef98c3ea7b880ce716da7ec9fa19f05b4b598cd6c3e4bbf216d0a17edad248b503db9a68ac237af9c6158d9da7673ad37110356a0dc4f5f82e7f34d8cbfb65074205f4100ccb64f96d03d01556886a30460346214655d14eaf998;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4f1885f3c40352c9ff1ff42ce9bf2db3ce113c71d939cd668e56ce209010acca5c59cd683a93e57c65b60a2d6e178200cf5a46a0c7b872a6215e0e7cc9a3388921a1513ad18c429535a9a2c5b1bc7aa1a8e19413a908d14ea801b2bac2835fd4a01b5d1afdb37fc47db3a883f3ee1fead2064f543d2d3d42eeded1a1b469f3f6d0a11a960dcd82eec2a93f0aa083c106a0d05eca2904e7c728ef1483b7043ac4cb0d7b2c0a685ecd3fe8bf732ac2fc225f07b3fc345e0030b4032bdc3c6379911d2207e8d4b072503b8b5d940eb08840998854fc346dc3bd36174ca7b15be35a1f3af6e2b58e1a92fc3bad2fb67c7d1ff0096b566315de50fbfd1fb0cdd498174ead9b602653aed54e62f97d711c5a3f2f1020bffb85de013c3b28ee13c831be85ed767aff0747148c326922328a130eda2ca11842e8a6298ae1cb5d9a438aa9c8a0619d383d1b3e4683d4de7a7f6e43c157e018a0c8da57a81a1263a1a5212d0c3e58ff3916586aa50206683251575bd3b5a3dbe860c20274ecf9c34c04410880d24dffb9ca18f3f1b9f02f64da656423eab8e3c89dfb082164769e9b614443e29dd0cfd528e4e0f9bbd4035eb3485839cc8d2fb508a2addd625596bd3b88c89fd2b381938da112aa7f6246c3d39ea65a8e399765a51e13b546d0a4c3259494f8619de204231ba411a88cd7ca1c73b3a45e1c8ebb6a7eacfa5fa9798049db6e0ff1915e0c6643c7900641b7a9a4af08377ffbb3b001937b13f896bc231949943fb168b94d4b155236008af20b00909bf95d4f1a074aa7a3a1f2a51ff70ddb29a8f3969b8deb8c97fa8fa8f657acf093698b6bf9b7a8799b25257f91dbe3f04feaced4e53516a6d26b8db4a6d817ffed351bfae6f445ea7de450fd21edfd606201b8b946bc29d4390bbaee96c05ace2d17bd3b272d53bcdebad5e029b7b67829d67216081d942cdfd4c363d1194cd2283981d17897be681f0be1d8adf873977518c79a8ce81e2f3567dcf86c5f0877c158471a2fd3dbabe6c823e44d909f9cfb2e48b689c0635a040e299746f47715b2a44712895774fe4792ce406ff9a0f56f3882ea62921724bbb56f96a0a1104ec1b478f413512629a347b1ea485a0680306966c75ce07a58871aa442d7bda4a5ab26150fced4632fcd428da019dc52887d1df64216a6e39e845f7102703ab7e688dfe84fcda0b3215396ce9b4d4da1a1300f7c7b97e0cb62aca0ff512b1c13a86cde9762f0f995cc3c52286aa208f96ad12a8ef4c1c2d94bf146a25fffc22abc35cff6ce19627bdaa329425709a4d7dc1dd90e9ede581b3ec7594ffe346ce428d0e7f84a5c7ff3c0ad89380b9314fd04af0aca78e81350c29d4cfb9430e45f2c2d1a4780b3d41839b4107649eafc584f35112d5f3657af43e0b1f86aa58c8493730fb03222145fa35ead0f8e292bd3e567;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc08f1edbe7d8d7376778ab9d02187207228b18fe36b4d9df3bdbec8639b7df3ccfe1e2411821b01a1dc4e25007f18e09b97e330c011316430bbcf3d92ab2eaadc8cd62d4a2d9db74e9662add51493fbfa5e8e9bdff60ff789b94dca72f987fa3560a5c606fe4f9a0d4b9d327795372b2e53e4b5811a2ff251fcec0a7a601cc79ddd438e572133e5723b7932bed5e409e78207905c0b728d1c5ee6448eab633af820f3c5d97a2240e411731b6895950ab661a17c314c68ed993b6a2806e78d9adfe9d2f3eae9f0bfb5478c440d3b075ebb2503fb9a66862509df155331c7ae7aae5c17e11734b75dda7ccc0a546ab3f1562e2167ddb77e626e6eacafc86fbd1939cbc23369a3a64e45638e0b335136b8d69c25533f5b8e6f2f77501d02aa5ac0480e9fd69521669dc63013c007e729ba7124ed0492e05ea7a43e7c9fedfdce01ac97b366bc34e1a7821f9f4ea5e82d73845089c60151b7744921bb98052acf6abdef037aec6cf592006e06b07e3f83028d8063c3e209ce90696cebac9a608fb02d8ac8fccca58d3c2d4e1f54ce0d4c47e23554e6472f09fb8636519b1920dea33fbd7694c1cdcc657ff35795c33be3b9ea7c4a1f03b737df40a606d999b774aa43dfb48d28a26706d0d5c85648b3c6175ab12536fced91a3d03014e9124aa5de3f3699ebc66207b0db5a31c0f84ab416378aa5f1e47c7a702dffb7bb8260526e917a860396396f07e0baa5789addde1264317ed250161d0e3c91e056cc524329022e9b69bc5bbb3a24c2da4a82f499c896967a1304f96bd83d9e4fcae0be4611a6b0e93114b339329fd4c3b99cbd6c53cf23ec6e264e9754edc4d867384d462c13283ecd20576e6db2c18204ece523c3656efbc9126c5373d9ae0a4d8a69f104e4eabd456888bf04f7384a93c1dbb9d99025cb27bde8fbb763fb741ee5f187f2b6276f4b5a94ed8e4adc7c92052d5665c90b455f713f1c7cc671d2af9f4ea4a50d3d07a3678e12b4bcba3c66716ac7f3e900a0f6474b76f31f841bac5d456b8908f1f707c386f58a281024bc5a14b5b2ffb1c676c0ef20fe318e0c7960f1e1faed855c8a617c09e5afd727745a946943d30d7561f6a664602fb5c2c47b14e6e89c1d7ec0f1cf457b5740e9f8390835836db9889fdd7a4fdc7d368172e0a4ef689bddb1fe6b60d59d40c3bc4265661050e2339278ce15076540e909b31ab45cd9666c32ff7559e02856813ed340cb89a07a323438cae312201d31c3d2a5eec88b9749762026f751535984721fbc9a04d9a7f558a5d746a0526738c125c3d587b82a9e73b34bc638ce3665635991501b0ee4d2d12b5d64d4ec72c08334c279c0273bbfc7a6dfe7c1cf02440958486444e3c4b970948e9f29456621fdf5ea0b4164ed73e03770eb8ddac74825bd911b85a2064d7c97a3113ba3967b6b943f76f20c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h77c7886641e2e79fa000e74b036facba138e454c1a5dca45851ded64ba1900c13307d55a010e0c1510f6c0f3a47fbf69bec5803d80b754e286c8178ea03682f230583782ae6cb1792e106562879138b3c9c57620ce3a86da0d5992a0597e0da9a261db32eab0baa21f6f76fcea8044ab86ceab4f77c2d37b86b25ee81fb29c2254f3103b4f32e62ecf33c5c6f211857bad74b5b5e56679d80fc6a377a2995db620a0b95c27eb0293d264792e6b87d824424793c1d62aae29bce1f6eb2f5e47943a911092dad8a5b8327eb0667444b64902fae6655e6f208cd1f8540d12833ee65bb1b0b54a13c13b09a51d65fa476b00fc489b19b7443fd683929b3424479acab0f37eb2f510d5c21a07168ed92ca94841b42ff317ad67741764b020eeaecde3a704cf21617754778ee776454506e93aa220ab516d37ef2a3c9a8e124a0643105de0b4451ac7b6f47ce79a2a92a8bbb982ff5b1abbd2aa9eb39bf4da19e4fb13bae9f65f24471ba7d4b2e77f2f6c36a969de2c25b8f0c78d833315511c991c73682a44d555885a28edd812d03fb289f970554248590b8ca2cc16bb270310f9a06d7d8e4f28dad0c919010f22934ed4fdef078d6a375b9708452b1cdcb8b1a42a8965b441237125148620e55afa4a9bb53812f97a80c96cb4f4f9ee3e0e4ebceb4a60c39cccc701eaab52fa2f6b062f782a0654866e708160111483ec0ce1d2330fa5528c6699d41f64022e5291d855265d22972e7a76ad2e546b8e7ea6cf9ffca470f3c82ebc8cf6fac61916c1864ef8c85a68059423100f109971aaad0a2afb471e4c18916dfebc97c279f5bb11f8dd67814b2d33aa91eb34e1376f885b6d91499fdecd92e0ac1381bdcb3efd12fa72c17ccbdb40bae149688ae90a549e131ce17dfb5b2f5e9bfb5cdfc475af878286cc469f0a45bcd765800f6eb7b4c1a1e654f603eb9bee3864b2c99a48de2c7c1c7643ff1252ca0fc440e787398373d3c03700265d89c8f5d284710f8b73ba31087fd2752af261eafda38fded38b841703206191cec0bf6838b641e1d992d2840ec367cae744f8c3f3d1d0c35d843e89028da5ad6563419dda11b93d807a123bc16e4815027d42f1eb91431134c4ca12ffc8e58c6dbbdd965ac806642b78e6a212eb9f260e66ab317931f3079e06620669816108a58c164b725a8f8d8605acbd7792c8c35e71c5f8e4139e54040b870dc6c2a5fad934d34465e7b9bbf93f413260998302bb1989c42cdfb95fd20ccb7f19609c507d54c733b1ecd270bfb878092501bc9fc31558382c32a3beb7d68dcb3f16704b61129220a51709e1c3098d5889d04a9432b2d30fdb1710ef75b1970300dea721af889ba3778e0760de6a5bad608e9e0586fda48376cfceb744bd5113140ff1edef3f6dcac09221f07aba8315cd3f92f465a4758e492f5d577be4b545f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb21fa2fc19c85e98945307e8d2097bad6e901566e242259c4611e77ea6e92259256c12fa81ef73abccb9c290d73a3b37208f7a78102ccffc760e3de491f5af82e0253d2a418f65a7109468e216b17c1e4c5f55d495d1da85713b4512b56f502cf3a482d4273d501f142fa81ffb667b4f395b5f4ec5e437011f1f2d3d7e7c98c57fb74b5cb5caf1b85f93ea33170cf9785e0542100ecf1f115ae331ceafba63ce659d769347eed2740582f216cd0aab3479b23a132aa730bb4a1c930bbcf929c90cd606dcae5ebeb957bf40433c75f1feac22bfc194b931760be4f4a1ed87db19963852ca2599f0ac17e6777a894392cf315fd2c1cef56d1b133e75b5d9935aa2d860b8c3e9da57960e4e2b076b7b98f785ea6785c899bcb1df5e6be0f4b2af3ff4aacc93a335e86b88efa6e9f55143ea4af5b93bfcfbd2b64fb9c926beb30dfe954f7f0ccb7d90d0ceefe314a813ee8ac4d5a15a102beb499ab9c6c1d7aa43c0ed600ed940d568ec7c0baee4d859d6ac9fc8946673473b03dbf20ab0b2a2ff63dc399fdf92add75234f0996687f4ff2a61b8f735990b7b9e88496939ad36750f7f5d6d2bedde5f4f52e3150248874ca5973202c004bbe7277d8e988a405291baa54bbc8e389219c899e352dc395a5c6f318cbe623f3f09d03d5f94cb79fda60dbe08fccf7b52fc702157316dd29a24f186594c7f723110dfa164109877f47a81e0e9f936176a5b2157a42b7e139990cf8771c189aeb06ccb9164cfdf022dcbab771a4b314edd54357b078f9b3ae77672a99a9d38cb4c87e9277d74291bfbf2d1e783ce05add722cc4aacda50fe4431eb7aa326856f99bf8f18ce4ac091999ec4bb6692f3e9f10a4bad551dbbd46974b3c0448b2858a55f698ebf064105ce038f4ee112a2a03a05a8c68ee286379302bfbdecb43ba0da8dad4c767d1ab2723f459fd5298a87ad934ab5c0f9edb77d7290f075574f6539b5def290e8c318ead1d8ef508c5258e689270f346587443ed8b59564b9cacf43bd800ba7449988a66d69d5d9cbd0e730a7278126831895bed541aeabc3a1e28554687d85a36bfe61cc5c7e11850ca174c61e71c1d82103d9242316ded5a93d70abf41979fefe26f3fe0027628e5dd1c06da557d3b96990b9497f1c12f77da39fc3419b70ed83b7eb059f9ee3943b404a731ad90664567ad7f363c68295e7b59771fb43b29f733746f3357b8230868d6ebc7568c51a95192a3fac9b839191eb4607e93c1f97edfa6a12effbeed5904415a30760105d0c78a1b48ecf6de9b8e6f944773d5d8aae18b5cdd437907f315b7c78316505b3feac62e4bc9b69e662975cee4d4078031d5fae55b2d0b3cbe15d4c62199b35c0a8be95387621a9ca0dde0341ba391111df88ddc130d0534cdd956c78267466e69e5ad7995c97f5da310891fa9c4bbf7560be805b97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4dbf7825d8ec519971b4f4ae589ca1db297e812cb9cca7b0397de8969a3b96b80af2543197c262840ca09fad75bb02fc763180d08271b674543a00e48af5fb95c3713fdf27f8661c3db8f0e65fa3fa82e3e7f8efa56a68fce30e8888afc16376ea045ec7d2d0502688211df5888c3fbbeea067ee6db6c3c6d128edc2b32d587ae62d13f3f34ec2cc5f63f01bc6384560a726cb8b7b23513b356a220495b5d8fa42c126fc7dddb0b43b4581c6337fb2c4f01447d317e0f178d9d619f8a2e99f962a8cab78e1f944861873ed4947cdfa244fbdc4b9b2fc73d2a26256068c5a56992511b956a7577fe2c826c6c6ca2809e016c7969671857b6fa3998528e54ba9542d9cb9f18d8bbb7e408fe0a269abe3b1406260c5df61acf51fdf94aec6d9d0f98fda23066fcdccf4f7d4503bd2e599e14d0bf0198c7b94c80241aec953060730fd0a5e028d7a25bb46e4c0d30bd3955cb9c141fcee7c38a128c18b1c2eb024f30a6907832a30613e3d58719dd70e3a661a47a48a54a85faedff3cb239a9dc0220d6653893644704eaab861d6b0ce025833032c0c4be9662964f30e916479145df52ad12ab84e7fd3d6d0df60a7a415ea1f177be90bac8ac1fc0284bbfa9af96225daf1e32289287987258ce325399cfc6b8d5511841694cb22c7f406cd665912b3b8b1f16932124cd3e956c61539fb0e85ebab92e1b0a2576207e2aab9b9a695bc77b7523d5bab5543f7ca8268ae768928c4a044923790d0019adfc1c2d76202af314b3efc68f6308198504de2e9ea0ade8b5e2049c87e21e0d519694a5ac6242177bc246117e8c582625b85136c0a1242453765c71a09292aca1135f5f83670403958c18e3c545ada4ce5b730d501ad7aa562204a6ce0fc2c146e0fb849031dbfba9ed68f4ac183dc091b23d6d8fbd31f85f57b4e28f2361688ebbc892827be5eea823321b2de12c79628e5cf1dcc58ad38393c4f8e53911e05e15c0e04f0e31b2133fd09f3295724576ff39a981b7319a734319f83fe1ee8bf71f8b92183828f89f6cbaaf5117a55c91fdf1944b58f16856f8289dc1aced051f23ced1551088d1815972c14e69af556e2e92810b8fdbadd3a62c7ba1399eccb2c525ae2c369e84eebcc86b9c272405d85d26e15da316b4169fdfb2b428e51c76b54f6f51bd36745d88130ae8be0fb0705178a8bbd4e95bdf436862b04e206792460721b7d84e7150c4dd69891287c2b7bb9fda6180797f6b262c4292737b5eb533b5986ea621eb0bfc4b4293a0c4cd719d46b498f29f9ebfb007dd78cbcbf2ef037612847015bc0d9603242e8002f5a2e574dbf0285ff16531728f9a59c6a08d7f7d35d3a7791f007d163f315a36a7fa48b429c7ec15d09675e811a5da84eb5a70b43e30ad3535e928c4ec399a5edc86274ddd24147072ab5848529a764f52c49f7aa07d459;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5f94b689b1b00ce48e6b812713d1eb0ea8a7e7c7833e8018d0d5138c1ffacfe75f60f9d2d7a154db56801b2c11b81404c2546572604ae1aca45eeaa986ce7086736c5109105ceaf425d641290995d5540cc845d31cf713bb87db936d820b43f56147f20f58c9c389de5b295aff0aad79edf6b40b17dae52aa710fb230563760aee78442574a9f358eb126b242037973ede93deb6e9bd27ff280ec16678425297714dfc3d82a0565104a5a0842ed335f196a71c77f49e2e91f665c875e3f7df4a7f5daee812b56bb6e6ef1efcb2ad6927eb35c8d4eec9c1aa043432d5b93a7fc75d502efdf213ef26738d22f3aab7bea15a14bc150e3aeabbfca0ec049fd35f84340b9dbbbcda78468395b9d1e62de6714eab023501bb46f1619f71b1be69f135488c8a5ef27a79e1ab07c7b80fd44e26bc248f94903b4b8572590eaad2af3857d5de653adaf88beaa1d70c3f1f99565cedb54ac799759e08ffb77b6a78f4b45ec5b8bf217b75a4ee98290b458e7731051222fcde900c5fcf63c457eed2c6eb3f17939af877dd19a3bda98c30a1394500457ab0b6aaba65d54e095ef73b691abab9f87099862d02fa3cd6496caaa8db0222859ef040a16cd1578d7a1c4ceff0ad8abefa6bf66549a8fd2199f7523aa33090f9965a66db868527526657eb887f985feb3db00ac2c9b4dc790c7c2a2fb0c8e7c304a891ca587c2a04f77f32e0eec0b2a9ba43b94ce48082da186112768264e7d5275caa4df948ba3a846a71c1393c5932c757718159b52cbd65bcce3eeee9b3661aed189c06d96a31bb72d85ddf729973c1970a27dd4f7bbcac9dec7e6d172b7393d579b4b1487a52697780ede931a26c6396dceed187e6a8dd18486ce175d599eff05d10fb2c81b4fdb62b9754f5873b704dc300c82c7df0544e04ae6fd0cc973091459e8043b5118d714386bd644c0766c5b80c3d87bdd52d947e7486b2e9d740708ec56322370d4241af1bed64569efc0935b7c90c3e2d9f771f87adc37f3d6157f20cbc8081bce75efdaf88da8701248c5b27596cd2e74090e3ada6cc4f99a499ea15abc92ebc7ddd946762bec65199be21e4f0a64cf49fe676f8c5a8be613993a0ba94f3a930b1b3cd79c80e88b4642e96e172150cc08913bc1c8e23c3ebdb9e6f81ec495cd94ce6abdaf1b78f13849b1f66fedb9ebf3185e833ac0a1f53b98f8b08bd24d4cfa8134b045c271b45365247ac4e9b47ef2e804cb74d136e647ea7529677c6468128c5bd2e0d56b785b4278a29e92781fc76ce61b720ddcbe0d62423386dd85aa38058288f43601559eedd8c827789045a12765125046d9c15b5ad4b66ccf9ae1b10a3cdd0b7dab834bee4c16fc98cf63e448705c22d7f3cb5341b9dd362dcf6c2c22f089db6074c7c022fbb6e8291fcc1e174d676e5e4454837b396524a8a9269ef91f3b89f8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5858926c0b2006ce3a534b035edde2f9ca8c52ebfd471540ed50d15daf44f6fb9e62c422e7a736fafc06b3327883ac15d6ca0a6534f5f785fd13afe0f1f1ed3818600cd12076fbf94093c63f3b0d3fbda33ca35dda6158e9377786cb40466f0b5e9078f7a8fbfc576f9b014763994bf84440512808470e3110f669dd07d6f8b83461c4d22f75ecc8e2e6216c4bd33f84c7371c25d1f88c89642c6244c43230af0e20918444da5a8978a7c26bd8a12f0aa4f28f768bf88299f78479800226b75feeffc813269b82e92ffc79922f1d9e6698e76ada718ccbc46fb8824ba3845df51bd24d474796ae495acdc7c0cabb6bae804f8d0fbb06f365aff0bbcf0dc918a29879fbf0e79e03a6751f8e3419ac60e08f95f3d49c7aaf865384f779e78f9860de8dce8695ac1b82bca06d52005ab40d788f8d42bfb8d99808d51bdb016242f7903c3b43762596f2648281035d49160c69e7b2260879a14891b6e03a02899adb5aa1e8975abb231e5195be54c0acc2da5710e20a1280c9c1a8f8f34027c4a398b81abff6765e4845de20b877f786c3279d5770f306f44517e3d0511de6311792fe124ea5fe843eac8611ab7a0b1282e07f50ce3b380900ee94374fddc38be8674916b2c1b27f2c20471151179ee55d40c2e106f41e9ebc0b59fa623f6916c442d80c20279c6b61e8d4bb20858934482f66e2453ab4d1d89dbab219f3fcb8672a55cf38c160db5b753ee5cb0ad83775e2a88d3f071d7b0c8adf030463078dd8430bd4445a98220b2577fc00c507017f5d54096dd06402938eb9d9e7f395c60561e58a93de12354c2e2e933456eecd1966a4828e60d32b44ab3cee330f27e99badbd9ce5bcd1441fd89e93f0818323d3a82bffac01ca71954d94edf13c35520fe9aca74f0a767694bc41f89bbda372208165edfe3b2520ecdc426e21a5ad2416165be86879dfbb9dda6da8368f2346f8e9438aa9bb1f13d7e123077e7a4b1c1af03e3b01ff6dde9c4f16d8c6a00f47d0e0b346a502db5af56169243207d4b962f20074fb9bdeb0605d6c6a7be175709f7eeb2931587224a257191ef1658f44f8e275d07711a527023980e29e46f74d5379d15d50f58ea5942542c5b0b77e5d27be2edb9dda48c60f385eef29caa76dd1f33267d22121fea64de4e4030512d179cbf23fe27150dcc5fe8b1cf66c5aa67e09296d41f3eee7d0a1e8e7079341032a8d85b96b317a1814c9bee9c575f29e9cf8ba19f9da87ae3a5e5a5a92fcf69c234be38340546db531df6de3a4147d7325314901c26ded2057ffb8cc9f3c99bc321b44260db157a0a64034764d84ec0f9dab091523d40128d31b067ec29069072257a0c789e3dfa7bfeb8f332d8cb91782cad3fb29d76f6606e9bf5e9d7b570fc9eb0c21606f3884da7ad79b9c4df4ad219bdced8537803ff6751442f0de8c568f48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8448561a3b2731018a0e09283ef5f04c97e1a339930e460eb3503a070b580d7c2922f7955193416830cd59f247884336aeba8b7cc1d840076b64445b0790465092f3e16ae8062d777a6e5d589b4cda436f30ea59a304437c8059a27422efe192f778645f0466d1a7b4b55d3e69a9b068572a95c8c201a832a2df5746747b9da0819cd04807e1b48c0a9bf555cf1f6804f61bd87ee45fc5d58e755c47d28c2920363e4d1895be170b45135e0132789f377ae529e79978b834b4c8aa7f623caa6d60fe10ce2cbdee6905e8d84895bcdcfc3a50e80d83aa6fe7383044d1ce71df49123ba96c3c2a7e9a4649c58e46d1eb85df457b45bbc926a6ec98439119d8e19f835128bf0f25c88515a8ad7a56608227a5bd89187402306a6075ec51e06d9a01c1635450d05f70f2854277e38173e34e17292fe32d63a64b757618ae73853c80ed66989986403be9a0373546caf1d01b159f6f3b14290c47408fc06b80da707b90a0a46b47518e46263f3e44fa7df6f625f1975edbe56bade89addf477209366288a6ff17f766fed6c6e3e8527e0bc918c839576f300768ad78c40f563871a82dc781717075582314403596f31aaf1ae2d871616e11166eb8a60ebd207054039f9d514887c3e7b2b8e448d8a9ab5d6ecf5e1da909f5c5fde5305c25ae56c9f29f4dabceabc608875cb202812db8cf9d0ae3ec6ab3b2f56ba27111f2416cf7108a67df8f05e495d63eb3fb6aeca9c9da22c607d8093b3e3e09be36389981f9ef9953248d6e5e538f7cda3f34acdec5a893faf9174d1e3850967168d7503eed04cecfada226c9c2eaedd7cf3c05f7e1d71dc8a6bf48bdc10e72ac035ff38a2a23eac5ddaba3be9f3ed7c9f53bde700cd68a93be4213d432b609ed28771330a0c0d00dadc8cf346c31c2cab6f4ec480c0b67ef531fef589d462c9a666986b14e32dc0f23324623b2f754d25fe50b7311e07e1b8d63616e9911f7cc6559a38d226d5adc7c2bff7a9436b35cde1fe07dd61d0e1f638b58401ccb77110022a8d93d5beaf85d43c9473285e9b8c61bb9ea4ab47c5a9eec5cbe6a15bf2648bc18a6cb6cd4e66a785136a0c84dcb66972bfd861ed6bfc35a558db1cc9a0173d9ac2fecda0f30c111ad0f6b7006cc580adcf67ffa65a8d434e66c947188005cc2ec7403b4d141f7b6b345e7b6ab34d36a40a1903bdc3fe0d67391da853937f0d14d04cd4f1b1e512613dd1b0b31ffbc4f11b5cca78e8622e0be80c0315b8b011ddef07ccd4aa6598969468817e616d537c12957877138fdc136c5415f3799ccdea478e8281913cf568a7db901d0f5ab5f183e3b4385d2d417240a1742a162c4a5fbacfbc3e568a7c8e0867c040c15f20112b405e20978b2ec253196d5510341c93f4794ce9b67a3a4a4a007f43ffc19d404eb8fb6483ca8e182c62113002cfd12add191b8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h578fba4b28f663ab4eb44dd9b42faad8502d1350c52c2cfb1138008312c80a852855ca50e43d7a88e8612151259c05bcbcb3f165b4a5f48ab53c8906684f6f23b4268b2eb0c50a3a53a51a5b466a52902fa8655760fc603d21b664c6878e69360f1f20df781ec2a525836260aff6dde5f01e41815ba8cab13fc9e60f04c8c03a27e57953d57c61ded924622e7c48e6cf74e77b0cc8b44545c9f81d07200631b347f017d2bedc6d1f56403e05afabc05757d2cdf93217dffd2eb8995014f81d1e104c815a609a40c8a3276726242a78f5548f92d741d069e49417d0ffa1085387b10649328513da4cb9fad9e5072c5a163591d216cff11611002c8642cf7fdfc98bfb732512cd33b5196c65607250a0692d87cd96668fb809bfe0b6d33d3b7ee472fb2ed5e28b2fc9d37e257d8aa54d619421974fcafebc9a57c47b246a4b5e9fca803b33a381d620178bf4fbac505d5b53b3b8e5dca38b90978a41f64a7c7be60665724b52697ca64c35afa97f2c926b38d273906d78fb41bfefc2a5d3172b2d4e538d2b2fb593805526b048600987bccc93f0151dbd4090783b910d09e8eeb890a8ced9f3c3afb5c8ca8a36f896ee3f8b1a38cc004b845a7150c01ec22ed4c045ddafbcd53f3588840b3cad17a453442ee272bda38edab84cb12256c50c1fc04728d7f9954502fc09d9d07d19c643b36afa62f46653b61ed4d03cddbb10fb700c0507c1e3eb9585a9e52e978afa4aee2c0da6378cad33b9d603c4c7f2b5c47aa3f976f82a9d1e9476f71cdb4b2aa8e654a6b527d78d6c6c0cc6cf4cbf03f827735145ea632bf918281a30fa6b0a12a009ca78fac9beba61720cf7d86fe294b893748de1b0e2373100d0837673e84504ce7f650cd5dd7286d6b4b24b0e5d97aa42daa009fb5cd4e192a5746c7b5d3236a7b51e0e431fa04c4e0403f2d9577ef88eed2cd83d7e12fb1d85c584e3604b710fbbc8222f2bb1d54c571aea25cc1e5a0741a94a248c0c384ea178bd46736913048fe14d62e0614455ebb42a82c44a77ccd0bd06ebe8608131e624f34bd6a482a934969ae36f051630fe140e1e91a0850f943ab76ed30912e6fdeff557a23408e8e91f22b9b3b067e8711ecaf72b8c1c7f8691ed418f55a06e4f91921701a702b75cdfc63553391a57d11ae44cc13c0bf3b726f7adf095a2692af90e66b0565c199dfdf506b5a785923d62ee1c52fd75b9c261c931d7a2e631f927e3dc7b1850a93b6dc78933040a98293fefdc9ed837d9bb93d54a25b5fa9536df339de3fb0e81bc7ddc1b8d512249e21d95f3ab00a327e7b2cd31dd1593df30b20f146e0c53cdeb9f70f32cbd72766424acd5bac1d14943f21eee9c94b7fd7ca0b4b5371b1205e2414a3ea162ce3f3dddb2dfbae06bddd9b104eec361d90c9a54bf77779c43996b2400385b84e98b8986b7229d9466;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h36f168246c211b447e605899ac26ee6592aa8edef7abe419cc4558b7ed97149176a3473d3d510052d518e0fbbadea20dff206c75c294c1b5fa63f5466bbcc33ab3035643942e51241b9e638b87d857167ee580c931ed644e9b87369285cbcb5613e2ee830d37aa4f9dd041a34596e4db376b8702ab6d69026f4685ba8bf7d39c4fcde0d557618a50370393a70a98da450ae1b2667cd7bd6cd035510d1fc79520cb1b719f21dad1c5bf734b8e377414835d8c7e95d052c0c704228f86ec21b6359056195df1f0915e693aaa9aed2bdbad699bc4f8a2185a0c6ea8a5112f10a71f2a236920f53bb5788b800619c64002d2735e3d0928ee5e2dd25ed69c7095d1490f79691d0d477708a8493c2221781f8b18534bddd186ac19f7a32640180e42252fb6e590b699a6847500d0e97de36b68855e7b129983b914edd9833dc2638cb304f5b5fcf0e5102b2ccbda1b6c4ee4afc3a28df5830e2e4e4753b10ae3ea6b9b274353d6708639d297f1f599f8cee3400882e6f72e8411b71199d07ed9062ffe7346dbb9b909b89500914a8e8a7d0f0abf426ab1bc204c5bbd143ddebc380f46a9a0647bd6809f2056c5dfb10c45b63833e5a25651150f51a249a45f22a157f7716c1a6ecfb103cbc16dca2379b171486a08c0bf960e89a03ec395ffc460ca3eed3080edb0ff91dbfd59f14a1ac77cb76f8a793a9511b2c5f10c7fa4bddcda0ff5c97125802ef2365aa13007d321284c7c1beff78686a53d1eca0c97402cb4bf0b124060e92d8b92fdc8dfe52459fa0ad47738a59014d19f110382664f6b6223fc3afa1431617a022f1c38de7dd11da4191a99f16f2ddaac855a6f39fc21bb1df0b6e84fd2f8515a81a992c0fd122ad29a41d19e2440372253c43fd83095687950f3a172ae1a47aeb1425becd1dfbf76a5bf4f436973b4b05ba9ec84c3a2abda697226b0cd0824b9f275906b55c705638648816fabf5b8c58ad83208e60ad898016f7a269d5ccfeca813b334f45658c4523c7b4a24a8d49932e502bc4108232362c6c046af9a69b006bc49183666d1200856a078430b84cdd9d05029fbf70016e10d73e0a9835134c6e034bd5bce12c0f4d5357ef878d590ad670423a761d93ca52649e9d43e0060230b2669df046ef4f4989aa86bea845219c794ac365d0c9d4db32e7a0290e901412b14f6618b9f63708ed4cf46fa1a9735b5061e990aaf6f5eda078ead82066b61a89ad271aa2163a74056ac1598cc3ca15ee3d532096e6461737342c07276fc0121ae20b9fecd4d7f5a1ae0d08261c30047707880314815cf80cc86f7066ae50ba308dd7cbf3207e96690e1b0a87d111448d42de7738e3faab80e7be75d8d8db38b0550eb76f222a28c08ebd2e22f8863002036571f99a0b755c8e3c33eff6d3da837e84dbf5991a90503e0f42d6ae9e5790112f773954d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h99e9cca4aa47f0faae5fc77859793c4a0f2a83a1300bd99d88975a3820ff47d42a3908da2577ce585b1819600d7d697cf0bbb9f63dac740668120437cb1e937523fe24456147e1923f3804469f82a872a49c75bf98fb007b79f77b6973a14707c25aaaf89c4d3eaebe1835937f52fff2cc89b73bb5dc6a2ffc1219e7287ce8fb2ee0b77c41cbece026cb0f59e95b02b84e01ddf28f265f3f1ac5657cff15f23715326909bb7814621e29bca61f98407aa5855e56d024e26ad5507c9fedf5ba7019f4c5ca12bde50ae5bef7f615dff38f904533ea7fbe85fbb05bde7944de779f7afe5f4a2e7f97dff70f6a547a889305b8b89dd40d696c23cbfa147123cbdbde98bb2e3ce84d27206d7a15d5568a4f1fa183c39052b18676bfbbd97c07043ffd3ceebc7685ffbafa161cc26d42977ca3871febd925ccfb4eb87e039effd6ce59331d4a670837ec801047eb4c69c3712ef1af65c3bcec26ca5aac86208ef8561c3493ebe409aba0b62e64e61b2d80cf2a0b8be3278dcf62c1f3ec1b89faded865a3e749eeb14fa2e9cb49f19a761151dda6153f803ed345a7aa59acfa667e0c561b6a061b55d053472b316d2007c1bc14dc5b1ae092e5af6c69691bec6aea6df27a514bf7e7f1061e3ac24d62b4e75f01b744e8b0bef9be309c37046103f20e0744383ac368ba5d03837fa0b983b32ef3242435f05d83962b76f45ebe7e2c67c3eb75c814bc45eef2327dfee99b53457aea9594c4b22ac6b8901e4b05002c3a06eab5b149972bf0d9d880a2117ef8194959566be2c46ec24c85abea1ff5d1cbea00255ded32a8111c899d288173179f9034101b6dbeb2390db0d5e083114f10bf8b104a531578ed0a0e66e41cea72ce901bf044525071b44d3bbe607404f84fdc5cb9fab4a7780f3b7eda7cc18ee03714a204b2ae2e08eb1739f555de4f1b13945bd57d8f672e34aec68b168e72bfc81fc7014736de9a01b4864b239c230fff814d379d5a5f9f9e8573f1d162a3dc2db2c00265dda9147f2087c8d64e812e6ea76081a3f37472e27e7b35112c89705758334241aebd043c222af60aba3b0c35e810d4060ca65b7d2c24ef71999cc8f13dccc9207ea96e69774304640c78cd16ac6c10286f4b10fe47062b3664158b3086ca29c27d24c93d3da1f6f157997aa8e55e4306f9277565958c9ab5d2462677ee749bf6a9638c7bc43dc637c3e7188dc704eca618b3507dacd2c652f8e0a6080eb949b8b5d571450bd83865e04609fcb07ae2bbc4ce37cfb7ae4de68febfbcde3316001150748375272d218fa9a3cc27e558321c335c35eb601dc0fc2adc457f45a7af83594531ea1fc7095e6b4c0da53473f88aceba2985807e8706ddb7691e7f4b0bcdc7b7de6a212b6cd9d0ab1cf236ecaa7608354ea83cd388c996d1b332f982c862d7b8caee546e52c84ca133a31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he2c2b25bca9e0cb9d6c178a4d2e39b0b30a4fc17d91bb7c1b83cf1a5784f5ffc57e5868d6ba5f6de73c51de22e21da78cb2c8911449249e216d40f1f05c92329de7475ea9eae490218865822759e990a124d03622c33134aebb8a93e0ab9b220ac963da889ac709f9bdec32d4a756315ad6f6f73990a0bd6f24272f5b3d72ce69108114d8890050d1462f89bac297e3657a877fdf83419059e7e8dccb0e6d12c1700076b3d8947c5910da8c4d0a316469bccdbe1d49e935828b55d7cc05511351e742eb2e028d6c8d0f19d36662943801cb6f4478fdd6dcaf54243741542b56754b996bd688d02d1608a76df67dbbdb7b5aad5590c63acd9ca07ab0d5a1e6cf86f65faf570d0c0f9fdcebaa99cd4cebd93f9d6d4b628bfb43752d50a34c1bba0e60fb1594fc6add8841059455bc7aba59f3d2d124e3d0f078bdbe67349e54d3688489ad6bbf652458738a5c024ff927d5c8f90eefc8f2060bb4424f442576387df64eea37ec8aa1a53ffa3f5069acdb3642bcd0e397d70893cf2e62a04ffd8da57e072a2c97fdccae7e04ed4fb38bf89164bd31959108ccdd13e017d8e0bfd5b8d567d5804fd354e328ba0f9527428f5d2328fac30716a18f47ed9cb1f3c95c01b4f31670064d0acbf619e4ba027696e33eea26c38b5e4ed4256e231b3fb7f814b62c32571044dd9699325bf3b01c46c6a2f03f0becc0e54da37d0dadabad21a928c1b707617d5dce65105a08682adc7ed88f61504dbba1be81b762c51be43aeb6d046466a7bc17b6ad6a98add544d70be7561ec5b4fd19eef2b9fd3b69ff70f5da52ae69a0e38650da35eab831a2570f86bcbbab8ebb1e71b086ecfc4104d9ff31221d12b2761a602fa355d9ff74c4c728522e155cfab38e0e4ed6ed86b486d6ed08d5c43254fefd7fcdeb8177c030e7cf218f62a65f60a93e3c4aa86e7f7dadddc30fe529e5e43e5d62572cf383c8b36235a49e13f8f99a62f878d4431ceac242927c9240aaab264deade2dee1a1e942d5b959e67a57ffd96aa83e61f151d00e4309fa02ad11cbcaf28292ac8983129d284974a1c3468b7f4b81a885855eabf67317900c8aac6e70c6e0d978275542025415928c813d63c342e3895562d18e3489e0c150440c2d528ce48165cbb88442651e0aa4eac2aa5ddb975d74680810eeab935b8ee1dc3fe7cd3deb54f22aa6130e56de8701e1401e36ee0fb474599c4ba6ebac9082d4517829b6a024d231c46c8a515b7bb57d9e32d1f5506ea12453d45c849ec531a0b014c82fd2ea325a3c78e9759e9af1bcaad9dd85c83a27259d4b4d1ef3fd30d9e72a5d1f8f7fb47a12318479c890dde4b5199ac67dc96399200a06f3deafb49048af632e5bc277c7ec1442d35fa5d143de06ce2b451e41856267ef25427665bd9ef7a7a6838865526a5ba646cef453a566d5ba7512302542e7;
        #1
        $finish();
    end
endmodule
