module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [24:0] src26;
    reg [23:0] src27;
    reg [22:0] src28;
    reg [21:0] src29;
    reg [20:0] src30;
    reg [19:0] src31;
    reg [18:0] src32;
    reg [17:0] src33;
    reg [16:0] src34;
    reg [15:0] src35;
    reg [14:0] src36;
    reg [13:0] src37;
    reg [12:0] src38;
    reg [11:0] src39;
    reg [10:0] src40;
    reg [9:0] src41;
    reg [8:0] src42;
    reg [7:0] src43;
    reg [6:0] src44;
    reg [5:0] src45;
    reg [4:0] src46;
    reg [3:0] src47;
    reg [2:0] src48;
    reg [1:0] src49;
    reg [0:0] src50;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [51:0] srcsum;
    wire [51:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3])<<47) + ((src48[0] + src48[1] + src48[2])<<48) + ((src49[0] + src49[1])<<49) + ((src50[0])<<50);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf653ab405d27894592e8e539a4f5471db063803c4810186c48a5310a82a02ce662435288805f0c450b999db994e3b50ebae9e00750f20e149dea5f54b5ed20665a28e57b4715dd3b9d17041f89060cf52b8093744;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h351321d07758c213b10cf321c26d7041bfb61c6cab3da1079bbb4a4e0081036d6ec6595bb5a49ec812f1a4c78b0794f3086eedca4000355a427802bc98a896bd95ade59269cb33037781c5421599ed71ab7c3289a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2cd9ec208fbc025e2678800a3bacf182534b2dd93161937599337df3cc868bd2f98e9bf3cf7d63b0bcfa318a59d03bad0bc4b2696ecb4e49e1fbb7ad99506177aa63a51cd803f826bd0a0bc9442df1474b4bd7ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53bff27a737cb02af546f96dda6bdcae3e2973b2f93683eb9216809bbd4313adb025fd20abf36e23c1650002fbcbb7f308213c63fc1c99d9cea145116a74f9765ce674f1c75861e431b03dd1bf482a7f82d1172d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb6be7e05d1128dca60087505bb388af8088b6e20c63d5d053a3a7ad8fc94343e4180a249677fb947a31be13e5c7051451cd26e332543149aa308b082cf76b15587857e28e20367103eceeed796144c68a711fd26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7242db549528c053976dfba9eeb09b16c58d7fcc106016a2bbec4fe9f1434f801487e3002f2281ae349c0fcb81e211b55df97634a24306773ebf220988204613a76fc737f3543193581a8cbc35b5179457ae1b5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3bbe42169dacd96b52336daff79e87bf4cce9a99fdeee0d0f0e3815536dc2a51acffa2fa58daea4ec08be2f742d9b8c6e779cf2b3346b7b3f34131b7e8003520d0fe987b757b647a7006e7dc808679ea382c52ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19d5cd85fa7759f04522008f30a61007cf24e9c0842403bd103e2035a7f05590de088ae45db8d6b14a56752d2e03efbcbc5345c464c84e8888a57a5aad9249b033467f6f85d4cca83e4e3ea22c5dbfce3d99a2a1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d20df5d77bc268d421f991e53fbe30a90dc21a12cb3e4b8f9c78f2019aa8cd134f0af30d60124d56dbfd1abc841235ffc90f44649ed90e8f9a0a994cd8e4486286c10bb147f02d0cc8d64d4f59cf0193425e0013;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34b9e3b6c7b7da7cc23dd7901ba50bf1f6c4013a43850a839823f6da87337d46484c8ed187f0d9273bac964a9a0f5454a06596c2643c7e3d600f10f010f1cde63ee03b9f6d5c9b2753535146445f0398cbd624fc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he95bbd152ff4b6303bda1c574f0a920f78852f4e898980b5065f02af6c309f094fd856e4529ff289ed800a7750a95f426b819520e03a2809dbb7589df793664378b8249640bbbd7f712ccb1e1530d9a20103b323c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4224171fcf665d6914ee6ef8c248e62db08c3f9c6327ad5549ac6b7c430aea345b8550afc42f4625ddb5304c500e90a650942a5cd53032c88799ce7d9ddcfb32b1a76995eb6674db1628fea85da5ab8eb685d0fd1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf78a280a6731285eee482dec0f59ac91b1e5027fa1ec9dc4a04736cd7e90f38a18db305c9722faa17799427913707bcaf5e57c84af8beecafe3f2a37840daba6ba975b2246bd15af95e9addd33e661309ff183b7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h351eea917e27f8460c35061a36b98fa7bafc4c56b533bb7c352bbf99ce818512422267dbea9beb206cc56d4c1f62117482d2e0e69872432ce8f7b1e0bcad3049e9bea4d3faac18badbe44b20e508ca7810bdf5320;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e894360742d7a4a7f8dc64797508b85342275e6ce90d7f609324a8f2182f2734528be22b9702da97accd2bc08b44bff9137468108f6bc0cfa201d30c591f9d2ae42250b4c0969e89c06e08e1028858b053462017;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf02f412e9a83ca2b8facaff2feba449a11926030f2c3efb9631e8416e25c46f5342d9e551712af85e894baaad32a0626aae1a5e295bc60bbd18ea3e125dd45e88c429103f86e5327e10734aae705b3734c82c066e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22c5411cb06879e73737f120b9a41ed73471ab1e9424e00003366f87b57948624d29a6ed2cb2727c066c0e4154fb3bbb46f380da6802f67b76e740b78842765bfd0ca6f871ce340060a9bbb05dba7821e9e501826;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc537440b822f117912716bf1a0663ce01984a49603ed2d35ac99a69f356bcdf9707d1903248f326f68665c8486ab99c49c2cfc4b2e2a2c6c6b0b47808b0f87d148dd8bb97f6ad8f88085e26ceafdee12a021bcfaa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79e1d0d372eacd67af2fd168d404248277814f81350dd350238e3959d2d0651805e81feb05886d79e06dff0652b658e5dad5eaeac4f550ec951cc30b368380b38eaa971e1c2046178b1bd4c62b7f19eb3f4a6f4a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf504372eb541fc7ad6955980f75542fd57152869b013a92c05e83951e94a8eeeedf86c100d8d424b7a66744cfa0d5fe7c6223ad5ae887dcd9d906adb059d9c9376af9c2c66e3df3ce8c1140e62d68691e9aae10f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h433290a884b580453aafc5dc9d37e491294410f503c3048661eb71527ba0e78d24c78908d71fc0537b7f3977bb29b2ef5ae49051e6fc2b5577387390b96ce0cc3b425acb1881f2433fc61801e0ecc8ee13b4f3b1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bd32aa57a2d7ece19f98056a39b5c3384e287c2f72c7b17728704dc208e1a317449ce367af578aa97cbc3a7f3708f89257d8b11e697e6a986572cccc73189b87fd6372287add06316c5bbbcf0f1624c439f0767;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41cf6cf1a9ce4f53c45d1f0a81fbfde467eb8cd37a5d961ed3578cbb6ca12b8681e43717051ccf27c3fb778d2eb12a732daccca4f516aecea2727e3662a02f7a1c44f13edae193e4a695af57b600ce459251bdeca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h933bcda085dd78d08ff3f559c74f7fd2740d5088b7f861fd47cb5f59590ff2f12c1ea77263c7daee88d74e50898e92d7b9f93e92cb2b6d934e072ca5fa774f3b46cb96688855a95c81e7080029457588a9dc2bcf2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf6a4bdbb0c7f5a63b3c5ee51c6d33bfeb4eea93525542ffb92d1d98185824ce80094f6e8053d26801b44c273160c9180ad81e527906baca23b11fb98e196d77d98ed20cff1b2f3533bed231ec623e5f1ba071022;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb49af2cf18d90ed102e2b697053abf2dd12d0465487cb737c58c7c5cbced018c939a820a234c6f62d07b9e530ee3fb048104d4ac9e52a83d80100d34f0ddff1aea5e442797b38405e86194ec5cee58949509e0c82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bd5644427bf7b7bfc7dd8b30ea909c1c019a877ff73214dcdbcf71c553596f89265195a75749a68ec6afe9e4b17364f04476dcc73487fb2e01a794519dc59ddbf1647ae6ef227d14d5aa1b3e402296128f57d220;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h234d3bb20badda600105bbb8083e4a28336889f9ba887e84040b020a56c1211a37f9bd0748e4408d35855b0ddb6002eb0f4a67d961030e4cf807c87036e8f5830793c5197ace949ee1df6c4fd11e69f17015d8255;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd597ff1e6bf9a1d5055352f23eb693c3cbd62678c5bf4fffe916c5364581a5d17d2e3783893bc58fa8b4b88df965040f93ba25a60034680c8fb53ac88e34475d64a4b2f77daf21c7d82c8317a0735a1ead0696cdd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeca8e4dc980a89d1e7d9cc4971984aa60b513ec40577005cd5f98d12101171856f3f6c3266a1a9dc3a6e8824f2a9718b82fd14abb1ac6770fb2c6eca5c2ef9deab8ba2c25d930b7dd32cacb656104d7428a16833;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b04f0ea2df460347b0220d21ffc0d0c8868024046c277c90ff284bc3bf7f14056fb3e489638a0ee41339184c46a8279e396b68f46b07b320f9f650bc260265214b0f783ecc38dcb29249f724b3a12d75cf897f7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c8d0608598ae8fd8ee20781045308cd309b87266473656715b638d563bd758d2da25211c57994899cfc1226742d04024792379d44aa0ec7f55526c17c9e06eb48afcae8f9ed8b506ad5f7f5522e1f3624f2a08ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe32ba207ec032a4bfde5d898df9094c5197b89177ca03ba38c0cc50b6ef5a4b4eb0e589d43a1ab54a85caa210266c1e43f13a3194cdcf14c3712f7b232984f5cc919c09950a8ed156e24cc4f93979bd17bd97fb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d8851eed38c1553839f4c4f46afbc98663d0d41d602d0ae7fd4021792c35335120cc446de82ad61dba85ee8057c3f33c137bed10cbc117eaaaa968ca399068ca1fd547c704e16d1ea8e9a8682c264192d204c85a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3876bd021d75c1af2667e533dc30bf0c3e9a66cfd1ae303191725f2bbcc5262e91beb22e39f96348d0bba6348d7127871c8a9219e369eabdcf24524b25541faa0735777a83965562305b9285fc9e0286248881f7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46acd031ac8462dc9bdcdf5a666f778d3768aee18b40f005ecc8d25de403ba5067fc5e335fa1ebde4c9f078d4766f33c78444e28385ba9cbd9c33f414a39b99f6c45cdacafa9eacfca3cca86d9daaa7ee8d6f3ff7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76238d8b022111611d13aacaa36d7dd7b2097251d48ae7fef2f0b892ac16c35b732684fe46c99a92abb61620fe966e4cab8a9f4202ba2101ace71cca8fea4852771c334174024269f9e281a689c1322225c33f07a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf8ac5193a9da9e04507d1112865666688b2152f1ba609e60bf6fef80a7831942ade7f788d3cb6f9117a8e89501327201d13534985886f50c87e5e034dff0da0ae9db50aadfb823eef2e9bc1b33433d43c462a960;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadcdab90d8f5b07e3a32f64b137d2c0d2318a5a3d9a9d70ee9dadb90f01d9de80895fce8d03443774569442b7e0c64c54ababcd95bcd65d2e788a42de1e5f27955765991d8579e32f4b20ae93543a119007ffbe50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3871d237921e84d40307d8f2dd45aa78635258d5e10c4ee48a19fb3d57e6c38e35c746c82f7f9baa12a1af8f15e62073f8864a91cbba29ff3fc5179abb9e23a596f2d8eb63cac237ff9af34b5a429d005734c8a09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb87995a527c3c1893f53c993a9f8566506885f00037dd0500bff35cb3f953927b976117076fd976d3bde950c9c482d985cd05a57223b8f437a1d9b1bba4bd20cccd8318d3a51891224f0c6118dbd9bc40dc212d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45c91c97df6b5281c47702049564cde1d6941494f30a34ea5fc7ed7e953bd28dd155edfdf5ebc17c590178018c94664416183616e5ff5582cd094717e72759632c26c161dd5027c01b0a5bcfd2006349a78c16d96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h118ef421f742c0d7cfb4097969ae84b6245478434d84f331438b5709390e2d26bd1d21cf0734df3062cf7388b767c58996e673225ed7461883f437a37804d561d3d8ee9e938a8035f6c53ad48156f3988b294375a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc2e97a6c171acdef8c361eb22ef35ccafc56509ee9c14fef6134f29fc62b139cd117ed808ff5fd99327d240ccbbe3fa9871d874c840fcf177014f9488a84884a5bbee9e88474e807cb1a58fb9f1ecedc37a1a124;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c640fccdc6e688f52a80a9ec8428382da9b0a106e6a6c2231210ac8d40e5a28bc2132827b3286bb21179a00f1b7c97f79b74b0cc68b9700480fcddcc582625589364e1b22fa3df668cee69414070ce965b2bc175;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dc5ceaef0b5e9ff6c68c73c6cb775b7c563ccbf8ec80fa66963ad5d8ea58a120edf5983f85d5ad5112f382a4d9064de10007e97686cff7ed19d695741ffc1015f45e3a8d770d67ddd82e7d810823c6843ba02fdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95add1a47998e4e2d5a39f9355cc7462377ee0bcf66a3bdb6e4675d9eba6c5fbdbf7a2bdadfe85026b05df3a6934e9f85fb5b59c86fa32f04d640952be29bdb4c74220a449ee392412d49bb0f5f86389058903ca0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha562c57ebbb5bc530cc659da483f6f3fbdda4c059312e49d021b387a7a7a34dd72754c9bc75ebabef0b521fb8a6eb73e96f37df4f29b0573751e8c8b317e5b240d872a150c290506a989f62e50523ce76ca1b0773;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ccc047b049edf475a0ce149995e50e8d8338698043c43acab7ecc8cc0cbfefe00009bc232adea625b3d044d9c5bbf8fa0ac66246329273896f305ef8fc86840e3ecba1d8ff166f58536306ff517c9941b8f191d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30db7058d42ddcabba4b5506e58a42081f8d09259e3cd23e42a689c3fde256b21358d07479ee99cdbf1a2aa942acf3dec5cae1c95a61d8dea0915e8ccd424817c3022c10f91e31dbb32a8bf345c8bba4365ee87eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37cdaed1339e5c80af34a9e8d7d24016ad2790238e651587843cba5f2f740352c946a844f8c9b867e79ba172ea6506bd81490673a9e2c352d69b81cf0e18f627f54fda38f44bda101aeb4091b07d34f832e36572;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8be96f05b0d2d1abd0f9aed986f4443a75e3e89c7300a81fb7b7cccb292badeb7b0a5659e5effc8d3ad8af03e2471e9a0d1c9efeb162acf257ce57eeb0e8d8b4105970921022314a36ae7710b7a62ecad41309bdd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d17215e6e821117d80666d457cee602c8201b479cdf81bc4fa7a9d7a8700db0f3a79a93480146062e983560b2ee17db397a979634189d2e449febd240ee18fbbc8022790fbf03d6d1560483181254194bf3fd378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bd3a318c47472d6be1d1ff59a0b3377ec58ab056f274f5c3354adb809ee4166bee3df08e013602560a2d79faaf43772efe404e547dc117d047d6405c4e818e1d4ea3038eb89c123b4af38e1a1f00fb9198986beb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h699e66987ae9a590c00e79fc37f8bdf0a87319bdb1b7a240ffca8eef9e7118b64d6be5df577c7352ba8f14814d008e3c1b8d123304b527fb34e71540d7d540aa9d601ad2eb6c893c4a4fd2192bc95d81ae3054399;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd617f091612972f3ea6d6873eec582dea78a086d8d511353f4144583da07e5c9f2a2180268647bcd8ec0bae0397ca66364af340286f5b40a5f3cad103f5ca6ff44552fdb38d6794a2cb3176581fa696134717d89b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdbd2f2e69550a9714689a999904d058c119a6a635d68e52f600b80c4e702af1fc125a897cef73c187dec908f33febca3b3474759245a7ce6caa69e29dcd3b5696b0784c818bb3b2faccb98b9b37350c1433f2b12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha18732b1fe2ba7db8dd567c72171775bd99e913423918da34ea94be7d54359f4d0cfb139d3b5b6e40375ac1c29a62b47fe6b3b4927a973a42710e1f694a15659f2db668dbb9988084bb7e2ed356ee8578c3f37410;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fc13f725b5477caba332cf2b40f7b44969b3edadbda88b1160438c40ca73f25d5951ae000785dbc400c62eaeec08d6b8dcf455ef43456bd23e434a1085848f4652f040ffda6e11678d5034654badf03794f1bdba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he97664da23880e078960effdc83f478089ee4db6971379cba11b1df4c4f0422a80be5d1580b8c8c0d2956adc4d6cee5d716632940cc86922df036ada8693221b6783912b52564a7992cb4498943512443cbdbf6d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c4eea0716a79fbe83e669ae315e0ea8c15e94d93404debf7c3014222f9bba91940f6cceb3ff56930faafd90109e6b670988dd17b9b95f5a01ea652e70b28913c370e6958f3ee424b703afa00d9ecf893d3a69b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2493e029b91e3c944bab73533f527c11ea68f6b0dd1b84abdd365f559569590ab8865a016248091db8e221aeaa42bbcea54105fdbeccd26ca969e06a4a908779fd79949d0d2c15e91eedf086f9bc426ed5acd68f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4c78a60bd8d686dfe65b792dbf621564ed2e7552ba9bbdd18dc3d20a63e443ac8c3a2153564863f86fff35a2a29c2022828b444067d30ac04261e603d18205262d5bdea6dca28f98c27d66d53bb4df99f5817ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf38404482650af4dd9ba98d9b26e4b21fbf7f62524f33d06582bb06191060b2b3a8b839ff035694f6af8034c06c08d16dd526d62b896c4fe9e0ff9cb3ee34feb94cc8964879c55dfeb03fa35fbfe80d3e0149af33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c3ae614e15143f962421dfcb3a14081472947e69b9461b2cf7e1645161a7395d856c4f056b5edf950ce57c81ece87eacf0115afca317816d419d45a3680db2bfd7e0c37c635b635069ed2b8638ecd6eb6cb94920;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec30757778f1006f817e0e381b94abbb731caecbdb94263bc720b240bcc94e0b099ee235b6e0f28850ab4a901725aa1e4a819f0a46585fd137d05dae8652b4d750c94d6f4e59584ae48aabe2ca3fcb230888cffd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbd6f1e6af9cfbbdf1056791d07c317bb86298d1f21a9e15715c5e0dbf4550b700b0cf3a2f5f184cdd9bf3b646affcd003082274d0154f805ca384c28031d06b2a364952358a0d71254ce9a422afae314989856e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82a1af4f2eb5f2ba417c52cf7cd6f1a6ee99d7d9fb7559cdc8183048643bc407793df4e2ecfec8536044603a901d722ab517a29bc9206538a815746db4cc44bdc9be33a1c740c09841f118dd9a35def37d7273995;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha21da3c086e5e52730949481bff2248ad6a6260247ef118ac558ea98b5d511adac6ce83a82f2128bd1a914e61564aa8d33404e2fb59c913ea935d0df2fa062b0d0dd96a298c546153a66978c36b4f5181635a6823;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6229ab75a1cd287d416dfc635bfa445bdc183cba4a510ba04e2c0a5db94c955460ef30154eb0c6e81484b619e9697bb39b95afef1146c7a0e83b1d0eebe03304590f7ab70b6e7f189f622f12dbb57411f9125ba7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5522b288b122641337bc0cb78407f46aea3c7361de9eb95f9a95c0061a3540f578a64699c377f2096aba62b879b2381b44a87aea693658721414af78060784fddda75de44217da73e42941535aae03fef074702;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c67df0ee8473e64d24903ca9e27313e8c40b6d166819c3d9ecaabe40086117da8a6e2b53aed86ee72eb9fac464d13645580594ec3dfbf40b2095931cb2ec92bc5ffd56cfc1642b65cb1129b28cce776d922f1dd7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd714e7cdf0f226fd5795f4e8d1989517b385208aee55d119f82ead0a9530ed58248d6ff41ac0348ed9518e9b92888161b4058b4d4d4a22f46c8e376fa740d2d6a66626d25ff848e14a10d05d34dbd6cc8b350ac01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha808255d16a50b967dc05459ecfca23c59d951fe628643212a37157df6ed6bffb407d3621b8db28333b8e749aaba5c72c7c19c9c1e4930df243d536408cefefd4ef8a736ab16d97d4647a4fe5ec522ff00b243e9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33258bd535363fb8d3a75a3bbdcbaa291aa5c8ce5b405d7c005f2a5ad0be559b619c83ade3c43bffde2da9b4f9c9a6becc7ff6803f14ab450c50775893eebb3b351242448599212dc4ceabda4154c56981799f1f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he99aa31fb30809e3b87c217f356743147cea0b05486d8e47ddd02a84939bc5fbbfd4b6b1c292ccfa5e802072594305e10b3e002fc4d6e572519db3cf6874d3bc7744d7ff40608f38c8c20df00cce57f842626fadb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66ffd2ba59ff7029bb80276ff4b074923d8e0fc72392c9d6e7df9742b174403a8b189883db22151ff808dcde7c660edb1bc03b9a1412c3621fa596af8e98f2d4f7b734e02cfe0b1ebc6217c57b0106f8df3802f1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he327b61865e1229fd974d08cdf99042b119c60c555b79e77378311b1406bbbe9c037f5b76f558506fc3b47c73da52ba1ef3fe4360e0474ae2ffddd5f307d064310ef9f18e67f2f85bc84638ff167d40d464f098ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3388753643941474d813d7693c4573fde9bc90e17ba2921ace8abba0f0a5143767f62c4c1a7b1454c7bc836a4e3e558350bd8deae821aed8828b6982510381d053fa02d4d0b35a72beeb41a8ca10d28b35d57498;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b111aa986d26ec8dfbfcdc01f8c1146df6e8b4fc4fa62f73fca2e08b386183ec355ecae73e0de3f5f93ed0f54302f0a296c8ce47ca95100599911d0de9cbbd7886d3716348ba7e582e6b54f4f5937a865c2aed01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd713d8dc09d688260651f0db347c3614670ec5b9b38388c68cbd3eaff23e0eaae41e50c2f8bff30e99d2b161c938430c4ee1a42c9e8efab7cc1656fd9efb6822397149b3920c5385a49037f80662a3e72fe0e9278;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21bd660c25f26ed4cac30d95a012b61889c4c0f764626dd2ea913d6bb63976026fc816fd3f02cac00489df80385f9cbde3edbd10dba73e96b4f2dd2f1cadd1763ecd6031f7d59858a1594cd323da766d697dd80d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b872bbde7508774f28431de64576f7e9bdb80ca6ad573578f75c744cef51a5079f7935ea396ea866ee4e0d6ee03b8aba826d8d27c194d46935e3f378c856e87e5261de98a4e4d1245b27468f79b31efdfaeb77d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28ecf7526d4baeed23702143ebbfa3d83aee20b38971054e3ef19b66e67260c023fb4d036fcaee5c297e1cc7a1033d6dc10e18e41dac88321a214cc387d0b056641b37040929d9ddf387fecf8f9edc97e6f6a4b26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fe8ad18f3c65143c7ed02dfd44dcfa6fcaafaae04c8e373ba65094c15d7d9d365571cf3f99b11a0288ac24f080c20a9383377a0012108a49b834875813338405c0768669c354b8cc429c7a942d396333b333df87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3151d30e0d8d73f6eb539041db0904318ab078c10b9a62d6cc460ec97155f1107a18b621b8290c9a38b2ce345d9fd2e1a67637b65d47974693cae77c379231ec734dd2fc24a4f5c4af613799d32736d31b7d908dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a05fae5ac6e75e6b8fd5a3d6ffd69800a37b27078d16bab50aa45eae56cba57d96c4dc36af88962efc4c6770a90aacdcc57937246c80997dd980119d58af2a81c2eb26fa57324413b7127a444e15127ae1aff396;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbd538a9d717f02791ef1adc1b94a855807bec8eec93f5c5ba8f3c765c04a2ae5eee03929a4d2bf5374ddf277b01ece4c9a3b11757189d644389abcd9f28679b90d934229da16991b48c12d4ae4d4e13b706bc5ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7333afd18e9330d3bb42d23a7ee16e4cb99d5379c450c19c55209ad2aaadf47ee6420b65e9ae2b10c6cbc9b449d795908f48084a846084deb2da5b082bb1fabccb79e66e31943ed45ba06df2bbd7bbe803ec63993;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfabb2a251412fac5384ec299d5b2ffd9385390233b412b0b9754361adf1d8ba81172f1b7ea37586cd1546a3762542636e6fdd1abb9409045c9c24a2b90b95da6e821ca229f926ce73d27e52c69cd48497fab19f39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h754ffdb9073b9455cd974b3d6f6736345b14424f4adfd3959448bb4ce72748c11f5b1c624c0dc509fc34dcf2c9437fcb7abc7c60258ea00c7e90208f0d93fb45597bd4c340005c5e1367577f7f22eb9a8e6bc2af5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h548e031f934a735a5c704d3480369b295dd04b4abf113cfcce18d86bc578c4c16f4368edbf626d6f4bae938c4da09e64e5c9cf3baec3cf2b8f5639cc0cba45f3c659b2cd85849d83a778bb5e66424eca9df2b3868;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9d0a44082a7ff8e44098ffdf6ba788e7407380531f899cbc15d6dd937fd0c8d4ccdfe82eae44a9a27b104f0332d121e739a98571ae63a4f634622ae21f6b05edefdc0b44dadcad33a79bdcf0b52e32e9bdc9ddb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce709c25cb3c3cc849a9210e18b4acb940d25bf73b9010656dfb68efc31fff605d3b6a7870c834acb1e51e2727f93cdd997f262498c458fa91f92f804195da33dad6a9b23a466e5c5ef3ee91da36c32217733bef1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h723711c6d501c0fe81c132d3c6e56b2a57810684b7f3b45dbdd7b0045b84f39e57b447c301c3f589e136fc2e92aabaaeb30c0b1b836d675cd77ff244c5350d6ab14f15b1ba4029a6980809c62fd6d181211231096;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc39d862e7ee7db098a92d9fac4be69095728721e40aa5fa00778fff18946d7eae550da9f31f529e0c0d68e36211242949a99c3b6dff55fb7b886564a1d9538488e5a891347e38e153a0119d065242834089bdcccd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc3b9562dde2f9e678b7d6febd71eb5732e3cdb351e1325aff66e765e3ab10c05b207c31e4ebd155e2f5e65816adf76f22eddc1fee74451a06578df78078d4644139ce46b9c459e2f7196124b4643dbee5d15e03f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64d8f81e90ea0cff245decd9a5e5202abbd8860aec29c82ef53e3dff069f3819beb6e53100c073e360f4f5e4ffb2291d5fda51f4d6fdad895be8dcbfd2f03e543d9da568fbb6e68dec95929b7a859d0228ba4ff44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4aa23bf2f5176493ecb4dfca6f2b25d60896bd16aaeaa758ac5b40b01b49b5a2eea937ece3d046679838d5339d26465a974981285fcc84e73e0ea49bb163915d1c1b62e9d865ed91a5a8123e66a737efbd44df6c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca62f2b981dbc0e803ff3d1148416205c8dedff8b7148d15ecfd4baf2ef83f104d60b123ffdfe59031fe52cb256f3d636998af7952b1a97187efeae84e35c2f9c47e61a6fd56df004b118a20adad4f266fa045b7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479d8f344c2ec8e8c36358eea1ca568595c94627a27f6a734bae7f92e0a95a7d570f2f14d98fc2cf0bef05c63da21ebc7b62079b788b07a104fa3fac14944928cf111ccce7fe458c32f2a967256e499c33057a019;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he90c222d7cfde1f11449a78e3eb9f8ad2dbbc313c0630efd705016aa0c2dc9aa79d42c959c48eb4b556ab1ca26775dca1dff696f05d37eb05dc212362698c8821156710e4630759c9cfad1c0f0f348a3cdba8c069;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46bceb7dce11b1bd3021dff9816cc0dd0dba12b88a629639f7a28669e51621fc1571a99c07c77035a0df53b9d67dfd7a53cf34ea722fc780f2e6c026ffed9b1fbdf235d0a1abd36880693db23715a9053f8bee47f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7b13f833ed4628aaa9cd8df4eb951ce2d1f6658df7e7b254afb3f2b67fd6b504ba043ac972130502e0a6c531dc644782f5d6ab29521134fedf4330388319402a65a2c312d544016dfaa3f06404939d443a818c10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c241eacf9dc8d08e7366085683b9ac05268b5e84617b0e947c32bb087376e959688b6be5c6393eb7c3b9c7fe633655bc2fc5a2a54d6922b2a67c179b3f209479a056a8b22d1fe3ebcfaef80cdf49c8ebf38fe930;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h274af37f0b7b937bc9a3f32a3a070e1191dccccfdfbae61eaa9d096c406f1c3ca9cc62cbf6d64abf2fe1773400589942400cf9d8e72c20c7d232071d463914d1ab3c0a38c9e2bc45522591ccabc90f71437d7a7ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h504ebb3ef9f1a1dd5b31800d33e41d1f3d7c24214b2724467f1be7227d6a48cfc0ca4f4f8e6da78f7e2753a24a47e71bb278438f44c6b79ceefa34915304680bb21199678a7fa7c458f0f02e8cba18fb10a90a31b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b2f15da3f53c57f921b6dd6d38f8aa6d96550053f8cb7abcda82bd259f5fc4b8398e1430170ac0670c0d8ff4a95cb8894423d43b288bcf17c1d30983ab03b0705e78343d3c089e5d0d29c79a80aa1e4e50212c84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5a65fd3de85feeb24eb5ffa55fa292141e4b4aa8c01b1467c86c10148f0158a0ea7c1e006698336834f3fcced16027728f640aeb8c0dc6e777e6583b01d5b2ede438ed062fb85299bc3d6ad15c04f92d5cdaa248;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e6f441250c15f48136940365024d71df991c5604bf754966eb9bd4530fadc3687918ca40cd439fc0e4b7648214ca2facd1d7d748cad70d391c0abaa862d8660eca851929588a4e8e4dcb1056e69d6f839ab7edc2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5e53b3847b0151455f5b5b789b8cc5612f76f59441df80a2e68839b0dfea19fe2b461bb41a6f7abf81b8f0450da551b1f11e68b564abf725986c3d96fdf4636bdd16a2fe761f762807345c3e72893ad08f016b90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaef3069e14367fc6190a54d82490776117b82f638e70fe5d1f2af49b19b263006c4f205c83e306f72d1340782d4dba3ed4777d60a7a90fea90a74f14332b4fdd4ee60805426946a9393527618d8de947ca1c5754;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a2730197c5e66df20250bb1b3c34ceb91b4ceed1e10ceacd39d42205ccb1226a9ae2cb39453d72e4727b76416cd9d4f25abd075c13cab78888466839b63cbaa9f02d7bc8bd57125e97858bf33d3207182a0f7a0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4334babc0fed4c5b4606dc9a274ccdced8fd1b19beb7c26d6e357e65e34657c860c23caf59bab47e06d6bd542140dc3b2d4ad78e7fb231082f74fee68fe3909e3e0db8ad85cc1cf7932af1aac624ea2bd195179d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb28c040d830e490b2765caa81d1d11885dfeee873839bac6e4c4ecbeb8579616101e5ccb9fc1e99f7509ad996d8f0f20d0b948680cdeaa9aff5dd73ef631a6a8a57575867359f2e34da237313e2445829e842446;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72fcb45c9da583d210a5ebaa07425f9c0c7b18415a315196ee207f35a4179312076e0e36743da36f2bdbbcd96eec81a4a948129b91b371aa49ee79c898473daf6d5211a7ba0075cf9f4a020b486f77d76a332d083;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dfdac0d114c6e125082bdfe5c3cb6ff30c50ae6c1205344950efe73ec8fae42bf1f590d6a4f9cbf6d15b2abc69d66b858ebc75d89db7cdc39d0f3d2e126cb690cc09093252f593b6102a8f518be316ad37847c2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3103dbbc7af1d84e1f61eaa584235606b22088ae615c2b27a57773c7a38eff45944e5aff5d330cbc524e3f505c0fe7e56decf1e43c106734c0d28e193ddcd1cc33e0c4e74c3af7f96b9e9b4491600ab76b610d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cd73f53c38dd4573546455f180413cc801d1c2175acde77b8a1ec8c2d96d6fc35ebed876174273e4c18791b91e7dcdb038d699d7880d65a3a457a79f6bab10255269d275030f732dc05663fa9e54451a35580bf9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2765777c8189f26f9daa9bc7c368b7c32dd18ab0fb568e13cfea7f1177872d3a5ec30d9b00dae2d5f43cd15ec4334efb0df53cb6fcb42f379b64728e5260ee7ddb61ab34e3ada8a7e28da8e0d2333dc2b2869320d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70e1c0b13d5a6e41e1e3f716bf632872110cbf5d150c9b028923a6dc42a8315ae611d58313b553630fc91f888256039d88319d6e1db37d39d0a9615eea3aa54a0ad030e686cfb5b591699c3e21ac42e47b56cd653;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e9707ed52ad313c8999cd5c559e08bcb8fffdb206feb580a94c3355e5b566f8c90d581da5834019bf9e0087d9d063c208aa03e49d0732c45909a9facac94ca1e780227008d78912a9e726432d5af45579e958aeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20518eb0f61adee0d610793c1f742e08c9488ff4e3fd8f65b314529b9ee64054a7d50eba45bd506c9577fa57f404dde9c590b19fca32a5f714332da09c71e6ece655b0d1b317648fe533e5eebef1d593a1508b990;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbcf40205c0cdb90c9e062eb42efa3cffbb313437df1d57a23b05e4e7c6980287b5db053d6e6a7096543494938021b9e88364562cded993d6f28f86a5758b2fa4b3484d214e1422d9e86ea53610a0c2c4c533c2ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2badc8c82af6a638f7104ab76680d19e5b16084303fb68e9db1bb9dbba0cb62af5e60a0b10b11cc9a1a036de04dbcd971ce45da553c3124cceac80db506d79305a735f3c49e7536b0a0373eb529a41f24e0a4cf92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1316925f65da345d12036afdb625039b2fff23929afc7b0385d2f5985565f5307f5d594d4fd3d0352b59a18be4dd75b2800246e7c16d801c740b8d763a70681fe9cc06d064fce5521b78180785ed72576de0a367;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf305f1ea3d30be5000de73b3387fd0c4736c9d5f262b62e5798d2e488c91012edfba0bd6444ddd1c3d769668d36d358b274076bf7f26e285aaff9c38061fc1ab3f91d698b5295b233809364e748927789f0a1e913;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb934784ab60368b6212daea35542a83a06efe43751a9ace7e52eddc96532b825450ebf712af6ce1fa169e9cdf65415c3e3a2ebad43dadef28c74f352b8042e7a065a0a67c013e65cd2c60a663b1ad0a0bffe0d331;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd95aa182ceac61bc0f69711d13d511751645b585db9a025bfb9cb5e775314f12b81a1e809099c99c8c55b4febeff82290cbc20d7b24255453bcd36ff33e046a041fda300ff6f7d2185c68523a0c2b8f5465b3c712;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cbdc3670a4653274f41c5d53533f1fb336ead9287dc900ff325203b1bf278375130857d31e1bc558b08ddce8114cf6fbb2ac2138c0dec38ade7ac148d748467ece8ef287bd4982f594f0f059afe5b7be36f7bdcd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bbf4bd203196634fd9ec62c7a626bfad96933043105263cf5d463664cc88ca0d36242e7505ac1b0d534eb2f508f9feb3f6025515757dd9bee1c78abdb2006b46a30b748d519253437a5aa7970f3ce228f9a861f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf61bc5edf9ff10fbf2374471ad9b247e5f3a173ebe7123663f9c4c2455b567266fa53f8255280d4deb06c05afa2dded5a5ef40ebc4e9309abd85a79ee372b1d9771c76d9fb14b5be593ea02d6397793a9bf4bd53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8db585da222c80382bb996f8c494b8273cd82207cf7d2980c9cbcbc5f2c3470f4f9a1033afd74efa5d59ce259c9311a9ee2a519b0753d8c1c805efcaed70cd3ec7fd5b921e2e987ad7f019a10503279a51be686b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda588c435577c4c2bfcc318215c1811362719ba898de12366bc52e26dac0fcd7736a78b2aac437da9adf0641319cf55c985d97c1874d6dc24093d9caea4e34da89a78980a44fd819b6d908f5946bbede65903ac63;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9445551d42782e1f690be7a70f32c587d03c4705077851beed29e2cd5ee652e9e6f8d3dec1e3bc2ddb5b2391ca25c64853c2362d7f609f1caac9aec0e02769ecc6edf70192e765d713011f6df9439fd7bb91eca43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38f06106b87cece52f20077341329834a038421206e4b88c90abf17597d42a41f9af53383336de51002380eeb3b9060d58a337f418d1db84336a8996d410102e26c40a8db681e5b95766bafd7f6cc72ba3e4d66c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d3e3e644218d76d8b5a9d0252067d127e9b962a418c475574a94b792689caab0d3975a700df46fdec18a49cc32cb880d93153340d601fbb99385561f2addec5f7fb8d5c665f677b7552dc4507da9cc7b2852a607;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87712481c206da05ef6cce5929d481c2810eb96f85900e20e78700305aa73fee5e3e17ce61f6e2d90a0f75efd065480c7326a7e902b6e87a0ea4529e65d05ddd0ad88f655cfb461de99fde75e1ef3741830be94e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29f846bee1b9fec3aaf88386c8084f316f8a15424131c3fe4c4e8c7d695f169bf3455d37cf40a24ba4acc3cf1e5459b39910d792c355de67c118b702cf0014b3d578320ec399877046b3c64f4fef45c9790c9a14e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62f48d9938161bd2d60aaab1ae9e13d95a27192e7cd09c1b4a00472f678ebab56907522aebcb0f8d1f2904d77ec2f5ab1098b001d15bd528930630861d5d187e48ba347ff78927769e7748dfec1a021e99a81685e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9b21097a31a52c9f21ca9b7b011ec6b70244985dac6a90a4b62dcd4fd2bcb9fad1e7d9c81628cd42b6fb431d23914b8d893b5fea298ddb03a14b311d78590a82ebf0ceb172186bbb2156fdb0be0275cc69e753f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecc6438e6265a4098b4306aed7022352011c7beecb74862947423c1811a07a31d7f3b0d578029b228676af6815807af19bc34117b5a294047678660295dceae8a28b4f6a5815cc2edc59e22c6a51a7490a45459dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h767a0c383d85b0f10201ab41cdaafbef2af369c3a1563310af5422da3ced7d951389b872d83d77385ca9d6dadc20bc52fb902c83a183422e52b78b82b2ca22000a00345910a8518b28e78065f66e039ddf50506af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9540e9923c9af1ca05a6a1477f6f8cf8dd0cf028b93c4f65d8989998bfea821c9d43e9767649d955d84ffef0c50ed908ec789f4167ea512eb6f319eaa72842f6f88b1af26d18316ed70f9650f51bd0477554230d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f95165025eeed28903b2a54434bcf7c2142ca1ec213cfd07cc7260325468131add0c139bf71ff7d39dfdaf60281e0c33ccd019d87bfaa5d1ec837891f7fa5893a863f7da6e92bbeb9469174953a5bf697c4c8fe9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16db244dd65e700b570788b7c1bd7159fec330cd5317dedb552bd6ed7530e7f6d7207f607fa18b535280ac8c3e0bb2bf6c790768fcc6343c06d1d059408ebd310686f03dd605f5cef45e1198d2e13ccd1e62b9bba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf23be2a46e5241d54679045c468bc2fa594e0c46e36e962acf64e27b1346b44f5058690694d1c1758192855a9dfc3fc7ef830cb7ac752082ac5367285d90b79c4d8b76cdbe9abed588b42a05877c70ca82ffa86a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h592bcb74f4737b5375bb87f2ff50243332289445622e5a0d2defe1a8b6e403e46bcae9017422dec7b003ee939bbb5d1638bdebaaae515d5b1d76932c6d8cf1b33d95b69fcaf962129fb51a1a10ff6365cd2ece60d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f1c4b280feaa7415deb07648bc417ce7f2d5f6deb8d47161cdde2494ef74457b3dbd47c40bd95c0520187372a1abf9a99040152a167656c765605b8b39bf147fa82b846935e7f7e3ede0e47988e90d5d7cdf24e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he51fcf6a0f82f9c9087aeee9c72875570dcd388beda46943d6e322192189513455716081cf3a496ef941fe5e485606ab3f764175f9735afa71a49b2b5e4da23bec9daea714a4ae82d10de26905ecc7c65d2d18234;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4848cfc2c5b98fe5d30a3e7471b2ec3ab7aa6110cf45dad0b4138288ab4019874b171fee16c2fd94bb156d9d56d31006405ae6a626bf5f23af65c7b41633acf3d54326187a5c4c3a364703440e3a64b411b81ca5d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba9eac86c835dfe6f3a99eae22b7f5de0945b4764d910b1545a621090b7b46a8374a141b2a7ba6051a9df5c3d81167909ed05be20ec6eb1ce79fd7430ffd9815394c868f93f148732e3b2bb2d778456d7eedc37e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9564fabcefebe14bee2dc2d6f4febffde85619c65e810b40c6a6ecf80452412dc26d98cc932403d96c515431882eec16425d27763ffd83cec2a5b2e155c91cc1e3807772fcb47af2f56c2bea06f75c2158e40e43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68a25d110a0b39a54f4dbed911b1e900d5bde56fdf274c99427b0ca4c5d7fdaaceb258bd21f5217c519db99526d686363aabe7b7839034dad3d4022236e40cc017fba32e2064155ec59074a498b04dc1ee48a77c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2ffd73b560e885d2fd3634e50d6417a10af5083ffe485a0cadae869ebfbf6a8a33099abe3de7b941db9c1a57462954a89cf3e7b48eb8a731c992e3fc38924c30cc01f45e13b39f5d68ea6bd43ea16e94180eefaa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h340a0a33a26bbd3a81b476787b11584c1e86c5cfe1e74e7db3d73261d8106b12f5ea0ce89e2978ce519639a6f59c0e188f3cf3f9cf85667e0b5e183ce3ad684a5fe0538334a59640fd01f46a9880007e8ba6b699a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6626e327d5f6e03a6380797235c339cf610a8a7e0c0d5aeed8461612f8dc29476c9f6b94da6f72fcc25ae278165508d93b70fd3ad0497840abf4d945b63805cffae8c8c3b3664bb4470af0da585225218e8297729;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d913a7e01aed63636b8fd6a2874ecfd71c1e579b08a1ddc38e9eec262b37695e375aaf1bd9e1335e2cc2c130b2d8e984183fbb739933b5b2165eeda70fc0d3823c68e6313a428940def6919f9898b54285615370;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5fae0b2b73c112df6ff34854e097ae02798d7f60b640eba79335759a7278d8939a5f30b6bb88fdd0a9a0c2fd860eb49cddd0a114c3a3eac36a2fc0761d55d3d436c8a0c881834d994a2b79e1c6b88bc9e825adc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb03efacb2b36e58432224424311573887555dd8bc827eda1cb3dcdb27587b16f7253c51697a8b5f3d52f41c2049e7dee9fe5c56f3e2fd6465765fd8c6611d376d3492e2b19da94f18eb3f26829531d9ecd9d2078;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7e226acfa2350fd2b3b22063d3cd079e1485627857431fafb014df8d0ab17bd1ab58553ff13987d6490b475e3ab1fe8360e195e69be3b0d93b8992e6fbe9b0c2fb442f0d07d20df5171f7a6501d5a3b65b39b806;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc905128cd103fcc9b4ee9c66137f2a8eedaf1096e6f0909a10ef6e1e8755ba6eb0b8977948ba7d510ab5e9c4fdfae5234ac4d3595d4218fbddb10d36fbb9f08bfda16fd19a011451ea2f940b7f8af946b8f5f696;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc8f7bdcca62162f0d6b2d01a808e6eb13320ea52ba6bb43c2c5c3d17eac13723696b343a65418221fee097a09e9b20d1b2c2595d00ff1eaffc6cc7f08aabe0e256abbadb5876cafe5e16313c3d488879408d823b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67c6a1be703cf4923e6bd4b3d316279612d4b746fedc0782e4a939d9674043d4303976964b8f1a2ebf422d94091c5eb43f1208e8e6cf5bbb60611f17f62e3c1a57ad4a698f0a91da6090d3864c13969e32ba2e145;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf171ae1ef466082027446e9174fe1c3385ed5c25ae162d0e0bc925979f415c3ded289d3e95d89c4cc8479326edac9d33e3f7c1826b62961f51feb7f6e2f4108dd1fa5e8d83e4828cbc07109400c73e435ca422571;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3690143a4032d0aa97322acb1b53fa3171be0be0e7283f4cdc69b52ee230a4c30190c27f98c0d7208ecb221c54fb6a92e70f11d51e09683c42ccca161ae3eb56c43e0d8f40535417b7361c86ca979e1191a35c121;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bf4e3c5c985f055a68c27325737ce9710c03ebaceed69dc0031bebf100c54267e9dad472906291e392599f10cb87d05d48825033bc5c7efddea007d958db2a932aac9665915164818ae09de651cddd9ad4023597;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h627fc8ff98ca686181ddb783c168cd15a094f4fc5b8e43fdc357771e616e10764151d6b5d48e1792010b0f5f4a0d2477f643448d3ed8f47c11404c41dbbac3894f3601549b0d71486e2d06704c4ff8aa2908a3b74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb6b26203102577ecfc1736028c531ed7e319bab967699320ddcca813d4faa4f749ef0090ae47ce0e9203ab1a6e51e92fdab9e711d5afb17459ce314bd8c1c4a846fd84bf964c270ceefbb9dd1af1b0cec5e7eb4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haecc515c8d7368a7206398f0c83dafee6868104832ad17836bee4c8bd3dcb260c6837e71a27a107ea706169450a9179f4e77c9dec70a01e58f90a229303211bf2404051f4e532bd233fc66177925e3635b49b4812;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he094143dbc34953021df76328dde928c83300920fbe321ee37b4f3b0163a106e7859d6208dd0e22f15fd81bf5852ddd4464dd52ab2eb52b9e56a9ddb5aace82eb633eb2a22b9c15a1bdec6c3e16d40a006b890ef3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2335a101cffc15d678ecff8b54d33bd8bebe47b98407e8399711969f831cc2cc907f7ab4b8c780663e79af4db1fc23678a76e9685f2cfe2dcede0a6fecde9e82caeadb9cc31092b8d9d285a3fa6598078b3170716;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7b45c5bbb19cb32c4911015d131ae7fa1e663aad3a702001796409091716dc39c25c11461103705ce08465768453d69eb544278f46f88810f001a36ec040f9ee21f4255bfb8874bbc64fd3d4920c7647c94ca8f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43a831d4bcb675813be0a8eba3561ca123b3e6678e50a90ebaf1326dcb934c0c3f0696b6d4389036374584fe03aa114868d582776d5b01cf369026c9d0da3adc756c598cdd875801325e0bb7e1f7e3480754d2625;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7cb514dff9f7c40d8fe64ac7c5b947a585533b87037c5df59efb554f076626ab7b358ea3a4dfa6df7d2c22dedadbfb210259d8d1cce9d7dbedda4bffc015b2e5f2116d353d6a069216c44b80a93579894d97ed55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h141100bb1e76b973be202282d05da0c2d5b5cca6f270bb5e3baa6c906dd65cc82daad0e71ad1fad99cf690f3275e8e02139d877e7ab2e7d60e5124e77aa2fa3a8ec23b66ef9d6f6b2d4906c0b7fb003b35e817f29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h229a5030559d6cb23e901b8695db5089c4464a3add1fa0bb797dc39f995306bd63a75e3e3c46175245edbc1abd1bc0dd39d8b89654ca481d07c2fdb1f77b05d3ee00d8bbdf012e50f17b3e519b62592395e010887;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a6f6e590ffbea83b60f545d1aaf136515ea68c8e1c2107df8475de95898e90a98a2b34268efe911363df5df3fb8c09600890d92cde4e8238523c58cfc9249520ced8108520618ad5d0c31c8c0bcac8f44c6c10ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5599c77a30b79079af92e3749a55e1cd1329a93db35912951b58308f65d22f0bc0769a167484c1a01144ab595f0216131855fc460ca386eb32c871a09808d7d4c0ddb3ed56ae78e3e1bca2517a96c8e0c3b31e77b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76a7cfce9a921bf8be7683d99ea3f6032125b436a4046805f0984015b6cf2024f237fb11348b4c222c4bd43d32ef28727506c0f496078af077d469b498627ca54a9308085452c4444bc281df0867a4e0b9f362d90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17f7c5bab3125e73c3b83f9920aebc0e7a1878cf50e9481cf94b473d3a4389ea923d32ae769255d8ab810ababe8f5d4a48c0172e3c5b97c02c353c639765323380d4bc5c548245e2ef4b79c58c528310998338a7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9295af99c2367f467fbf95390093b7bf44f9f98ff79f65f6d2cf10873324d8f9dab9beb65103c950d4bb82e910ce465a19e69f4345f7d3198f9c8e78ca95ad5ce93dd38831f6dad779de9c769704bca5700fc8fc8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h111732726be21bebb7ded4271490a0d70b7321f2c382b211398ee6339a5c7ca6ceafe99a917e830a5dd27f515eaaf850fc91225976fc0eef43e00b232ecacf415b5c95d62bdb099fd452281e7a68cd9f8d3758951;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5836be9224a14b1e372ad85be1e3d9115e159550b76b65c7a139e6718ed63920afbeae427adead3476cf0b47e65bb177e11658db2a6b3d88b5970c1f1b1fd7cfa5b9961a388ec1a82fe341b40998d40700b1b0a76;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeaa973994771bc5feda88068d26b7795efd4b90bf881ce90eaa10f0557b4c50a84443c52fdf76ea82df51490ae3d58880621ef45b276be2bbc6815d915ba427f117554df30bbb60328aa7dcfcd2987759729bcdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2005b6b06a6d5466b568333831108c4fb48341f27f270ef5979da34e8aa94d14a5f290b6874693377c72d28f2aafb8360df744930dc4dd316d3aa0c9541bc1db5722be88b40fcb87fe7f270abcca12c2401a8b867;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2e8b60a28dd510b7a53b9c4e9b85569782bc38d8adeaa0c46d86ec1c21bd9b4cae9aecf0788e6557fec08db25fe4fd482175c361d59b27bf3eb4af32ad241131be151eb0ed78ac827c7d9422e3db599a9b5fed06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5c9efb414ed2b9c8d9f30eafbb1c0f17f1359087e8e57357da206e6deaaa5664325a0a0068c301b0d5f9250f2c87372f013ec375d7025c399111c2ea47e0351b41ae06a5940d4f78ff3e957e1b3defa1513b08a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48c16875ee5efe423ad65bdac0db1ee143c7ba525c20951e6ce93aa82b4288643e0442fb3e9b14fe53ade4823dd31e702a5182c7f1fb8dc11d027e6812daa221db1e2554dabe1ecf413b8a04969a182852d85d66e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25b49f062823c4d5c5cb72f10eb681038c397bd956b70ef30d4e354c5a48e751c264cf860a2f36519f286a003889ffe76af398ac0298f462177ad274fb02b77d095acd67b82d92f92be4632f35bc55bab0b3582d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a928348789cbe6e082d0e714ff7eb5cc6f73941f4676c58a378465ad8a371420930747aa6f3d76b292b0509519b58f6c4a2707e3a6d1d08c6a5c8fed6bcd790c0dc10b996c149218b1e65afe2f9367c9e1b5fc77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5403d625aec1a79bb69b31836041dbd2ab4feae8cd3e1ab5c54f4e52ecf10dba3189e75440a601e0ecce908a69fff8d581d66397bed14da9d04706f4b4aef7427e226743e7b2aede970b16b863d0ae87ccea66eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8cd36d1829714e667b19a0429dc7b0c463f337a1c549606d89d744c8fd0a32997d26278cfd4bff80b4802dd71f37621c8d968b97785c80fd39713f1dd1666be90e78212942bea5e8a78d58ee51098b00cd7d8cba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb1740e9b8c4badda0213f3526c0e48d38b1b8d87f5b88fee534313970265e7b086790e67ab3ef22a0d1e13707b9ddbcbaf1bf0d8f30be1b6e04df4c91575099e6e81fe89b78ab2e663b0e660b65e82e4a25a84cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c73588b7c50ac2b95eb30b7fafc280f3f61a801f309d1d72accfc30413a7f8d503f254d15c35590e14b275f6819104051413e3a7a1e9cc5b1c0ff8573b228cf8fa9fb5d3921716f0c9fae3dc588fb80dd1d77b1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe958e90d94021f9a3470325057bd7a58b8f5fee8dababb337442d6492adaeae15dfc0233860ea5dc15d9664f772346cec821210e240909fab9c49e06dadaf96f2b71149bd9048827f9239476cd4849b41174e87f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46fe024fc8cf47394392c2842c1483faed6e26ca7bd99e8e251b9569f3d29a988e69f956240e0ae02484d720f220e107f26ada555c4109989a23e47c596de87a167d3e67a4f082a663f0bd7219973702283c30ee5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3784f14441c88e662df3b0917608fda9140214f7731f9203195b4bfed07324a24cc63eec115229ea70eaed5dc124c566ebcdbe7e019ac2c569f3db99a44e91618351261986c06b64e8780dcd6364c24481aea926;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h912f4c10e8ca6553419ee78a01d1b623582ca8213c726995afd1ddac9e9c89608efd89d54a690b370f75ab4ff28befb829b0c5c5a34d56e50fc33fcc782057f7ca8f09beba8031be00a5be6a059e96d5f90bc11ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7845a81189c611540c553a37445693ead30ad8c660f9e9ccebfbc1a11e64d4ae20f091ed5716d8fe6a4d287ece882c4ce2528a32648478c9d6b0e65e5c48f74e1303e30918e8916d8b19d582e5182fa83d28cb38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e465b05b6002cc0bbba82a6909731ecd04b4e022752849369d736c1877be5562b4724287a5be5a7ee95bc32613797c08ac803bfd807f8bb8cda7d50d7969a5b00cb26b51586d2e04e495af4c3c49f89398bda6fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f432d1c65340fc5ef3eb68515a9506fdc7d7dd4903b3488b56f6e1ae2ecbe10e39176204bf25395392993e6154932cdec19c0f4eb6b993e8b9c191686a0c9f60683635c8700d49f97c7c8eacba1ef04543f87531;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ac90f9b22178b8154408f99cbdf20f913fd96a3b097d57b7369fad2c4d211615280b2b5a4d1813b6bea20b2ff058d726ef71c0632caf46f4f667113ac86a24efc9591c09cb14f0caef3481606dc8eff4b042ec99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27f2743b5f6829eb0b4503bfb794af4df30cd64490dd2cfde49965ac0e6a65d6ff8700754ff59ecdb9ec95a87f51fceffe4279b5d6617ba379efc777abce0dc9f91c5f5af3d19c36d7bc8611b3cae94e432c79df4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h837095cd80d542525361c9ad74337d1b8fc6651facacb877637513c1069de10110c27f900442f2c309650c33bc8026117d6010aeb52835f161f9aef38e186ae823be61ff1130664c1636a1284753d56abfcaa62d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84a08eceb673793abad5d8bad521da0d484664dc32294539a4d96fb5fcf7eed0a45c0a1c8e517701957a876a71309a0ba0f0724e95a9abb073f92495f24044649f2981950be1007e3482ab4d981ba7f81e42a4184;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h644a643bdf4047f1e31df51f84dbc4d7b400dd6a8b32ef4a06d00e266233ec52040e08926f9b875a97d87b2d3d77043afce91edc844c102a29f385567a9e6fb455053f270180863924d586c5a98dae5ea61c7983d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2adbc181aad1e4cf12316d580967acf477b79a5c997177015839f670a69a0628ec92b58592686348a1f11fe208660429d9bcf9ea30432f85bdc0b7742216c6bd0c24fb5c8bd3ca6dcc50cc8efdfc1d982651d4073;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef886b7e315e75ba912b558b39fe279c3466d3dc6579b1784370c3930d3ac3e760d8a3a569cd684ffb54ed6c1ebd5bb6985dbd1d364ba2f507e4fba859599cdf447d350c6e634429f97bbc8d9b63482467e3ed726;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ec6c6a79f96c164de5adcf419cc2069121e4ec78bda3f956d85564b12da274591c4ac373e109f77fe0b57a46f25c186f6aaa14d50bd164b6e2a61994353c3a8fbaf086f06684673ea715386afe65197bc24b6a94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1770cdc1212da6fa57e34569a76c9d53411a9332f8c261ae774b50e437de75f3fb33f65a3c6b92c23b1e84b100a903f4a82282e74610da7b046733ce406a0c3da9fb8e27417ed11ddda689075e4ad4b22e326d51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1413a279216166bfc5dc7a095b5cb23e7e8b3a031db0797b3a4446b61c0540114d92d5a532b9be72f439dcb2789872748add35b764a342af52c15114da3e48fad7460e52268aac5ee936544083bd571ecb0964ecb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b2edc427caff1f44d4394404e86479561da740a73063561c77bed1318104f783dce07fc9b4e0c4fb0c34011fc79844b7cd8ace639a78e5dd88537d2ee346aadd1e2630b17457c652b81ea875f5d8215fc15b1ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8290748f49080efc4c7ddcc4490d470fe8a77974bbac04ff69cf914cc5b61fa77e0de4387d7723e51dda3da687e43fb59aa1af0e650c8bddd65b7f65f132fd646f10877a5fbd2781e07660725e93ca1b6ad3a7dd0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ba9f1cec953b3f7b7d9b9a2ad3bbcc71af2efb06f38f2f6a59e96df62e2cdff0f1b64fd01db455593f2bfb10a3f7108510237121a8e206cdb3830e88455f8d35d74b5da1efdee86e3add9bfa3719b67469b86d51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d34f75a8bc3cddba52c4c8cafea763f967c258271cc3900f1c4be6288bbe0fb60f25296954c9f427750af3bc0e5aad2b55d81fb7097e5dba607b57b2cd27f4c8bb25ecff6bb968d7cfef2dc0149a1716caae3aee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3d7391a8b7207b2e94845c5ab031a6f7793b632f4261f54bfa958febcd80d46c97e60e84fd37ac3b8547f39cbe24e7d2505cc1f201ff2df7821d7f6632147c2d55f972fd4d35485425263c7c07f94c47fd0ade6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bc3493b595ef05aaf798edfffd39cbf0244d2669e08df6f9f972911ead9841d39013331055fdaa7f252682633312bb334215f0e4fdb2160a384c9af70e90d5c4957a682845328374d1ec63d78270d747d26c4451;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93dee5556c1811fc176524f9b0439a2cb7cc1340115447b44ff93d74a1b81763b97ebe1e193fb56c5ff8fe5ff9bac3a51d398c83622e4f8d1a7d229159c60b8caf69720282ba909831e1b0ebde9e01bf0b9e8f1aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h725b7eb7109f76b77dbc242bfedf1663d4a268fe7b42c4a980578bd54c9974a23f3a627cd6c026c86f8739dd6ef4d1796c5fb9a8a5ef95ff17c06f33572ddc83a9366bd29b0272c9e2f8af0f70925faaf9ce5bab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7cafc3f9473a05e198b3b948ea21da56376c52dac6610c23c2b64ce968106858130bf3f7d243115cf838c96b4332641c7bb6497a58ec8c41f2122bd507ff579a8ac0bf5d59b934c3b4a90660c46ca2adfe5b852f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3dc0a4ea5f58feb9d2506d56bb11a79cf5ab291b9a96c8f89f64d2a3b9e4f669c5882b68858699d872a06ac1db76ab4035b9b5d8d39ed4b5757a32b21365988f76f359bfacd9a1ea719e1af4bf74e4142edf358a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b99536f3d42435bcad3aeae3d40f3284ea8f128a3437b3366081b3085150c2432dcf404e1fca3881b4f79306e0267704d72f08f31276970fcaa287168935ee1bba5efe6e0d664a252bdd3df059156e276767aeb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h787d121470a299545da919c9062d0b0036be7303dbf9cc87d05a1eff90c5f630e541bd4f461a86faf3ecc75bd17a74e5502381966eb02840ccb90fcf0b555706f7a9bbcfeecf52d143ee4b05073d19400c26e0314;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h268c1d9a6a6ed13e0097c96cb029030e09c0213bc8efa140114fedae1f336f33e933fb6c971a15d6e5911924ef463c6c7395f3a426571c21f42c4845ce1c83c72f2014fc44c6399271117715124421e43f69f0e71;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b8f6e04d90fa0ce6e1c93d9a9080504c1a516e08056da4b6f7f279df492d0d366c1cbc78b6b4664d934dd6ee0b934c584be900c07475a54c4c6fc7596fc697d1dd51511a0b052c842500d420275a430694851475;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52b19e97e789139f6dbf07a4ae9952c1441fe2467d962ef740a8e1f3ff1544073594f937c3b6a18062487c225aa43be3d1099e047e6388132c3e7792f60d37aa2942ca7abd10e0350de3d416386324a46a438a5c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc33220654581486759b8370c135fc67fadff67cb059102c1b046f4e14518d4b5f5bb7936bfa86d3d1846f1d54d0b06e074a178fb61e6e609c4c523e774174be6893221f572ccd0222bbd2abc78748ff5ef6fee8f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e2bb112e1f99c84a90d85fc31d0bdab0b4005560630785809a51b8313e18d468443b355ed13e4dccaf6f795260d3114dee1a87114c887fc4040698cdc75a32015e47c91878c21533cfcf9db147d12ebbd9a7a4e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bdb2ccc1027db5f3b8677dc6180a67a851d2dff4cd3e2d3a3adcbb41d5d97256cd10b8cfe867c5f11719eb2a9fb323e3d5030ced7568adc3386e0773a8a39ea43367109eb28a5f16bc8ac7498e69a4d8b39126b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h282cc1bfc2d818ba34cf6c72956ca81254a9a90c8329780e544ac700246738fd1733e326f078be1c1b544e9b58cf3fed9c405bfc8af2883a1a507cb48bb9d3cea07f15d3e7d529d08c9d2297969dad288fcf93c8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8407fa8b7f44d6645af6d4b1c3452200f1810c62edd447a3386c9592bd8df0489d8a8c4c15f28fe4318506574514623cb8246949ccf7f4f95483cd26585af83b0f359f03ec38499671034ea07b1861ee5058dca5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f6b597de659c5c667ab37ec458f7208df4ff3f0bd9be12fbd6e51d5a6b5960ccb7d3ea48d20553fd13bf3247a25d822a04927c020ec70105926542f6621ddac77b29c52eb12b466803c0a8f92094d44a3bbfb9d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had7254a72c81c56fe4fa6d4edd9b752c76273b4a01a202bf6640cae9333179f0a66d4f68e0662bf540035ba14bec32c99010b25f5ee5733cbaedd629338be9fde37b1e9e1ee18f15c954c466ff0b23c913036c195;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fed25cc4e6dcd0da958f3a6b4fa540fe351e846ec75934765494a46ea9bef70cfdef9ac276d5b95726b8815c5de4b82c0ecc3a66db4cef4a19312b3a9df77e65f3ed9473cac24ede4661d6d0d3e0e22cd309bc07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f089a5e4c34d442a29706a8a4a024a7a5d1d4b89067886818fdba1963f9dc84f95ae568b759724a819cc5b226635d051cee56e49f4ba7870e281e0514a8fbe2dd4c925c48c15f5e89f121fa4ffd807c5d61dfd9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ea9c01901cbf46d090bc91506bd0e18cfd4a6462e5f270cc0c5d84425828bd39bc6c0df38d05859ad1160f825fd1f813b58e6f7a188347d5de69af94b7698fc550f5dcff28bc47d03385acd5892cfb4efb0f36b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32aac043dffbb59d9694fc21c62f6dd00a467e3c275b96f874ead1d3267875632f308c90a075eb532a27de83f59e2312283f0add9bc7a62fae1325c634235d7e3a697130859fabf138cc05effcbe70a0e6ff2a804;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d10cfedccc8482f6f3969deb850d15a42d6922d1dea7986105b965eafa0a4fe00e9ecbfda081a5bfa7605f99e6a37427dabbc45473000225e27c0b2b3e2fe381e8e97dd7b9ebe53f97a048846e512c810266dbd4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd22d8805259372ac7237532511634e77ba333082f4ab53f5f9e5c18020335494a8754ad85ee47979b30bac06e12e54f4994083d4cd4f84fa97a04a8c02b424ffe7362b41abacb79ad7ff8abf8cf949f0fea3ea791;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h203eea4a7be826bcc106284ba9c52ecc654fc004927f03372855c58578f566ed3523a11b4d6206d9c13d4642fc6e405ba9341610806bf4f5a0f381e6ce270e9d757c0a5d4a36fb24745ae04ed1967406a01967a0e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49139356cdde2a12c5ba497bb25a452dbdcae1115b788db96823e2d2095f0f225d56a246f8ab76ea3459472eefc2fa964a75d8ded8ebc70f7ec0845a4d73a02e0bcb779f40da61affdcfe31a4a6974edc12220c60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fb6ea23f1ef1535efa6f67b1fc6d7e7263cbf2c0327becde7c7d0ca9710d3f75357b00525f1c5243f05b44689e90a9c9a0146a0f5716f3daeccb4ce76108ae93282fe26671ca5f781454ba94170338a8ee7059f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5c2fa13bd1efdb191b62324933f0eff23fac0de5ca063a3968a410646e2163bb02fda7691991f2d4e1ca30cf68b218ca2117a4e992ed3a7b0adde10a4e49a7eacb50cc013648d03fbd20dae4ebfbdf6f64221203;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81bbfb1b4d3a4c63547b586828ecf6a707634b352bc620f201b2d2351b50486d0bda7b23bd187e0458816eebe86004313fbfb1fdc8520201d9fce132ee481deb05e95268c4e53fc05d80c76b402e77741d5f7d19b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4c437539b71f17ad379a586a127f3f3779069df092de6302d15916567b84074e4530bd08f1cdc7ff3cfc14c4ed4397598ddae9f35d9680575dd15e3d8e50d1f8c6ba29f39a71fb85336902cd48c84549dd62dda7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd61873a4b62ac04f141c9ed14f20a2a67f68b2be9e7b509ed4b3d6d31e86e2215f94bf83e481f656812d43ac7816e8a553b9d6ee39358de7a1d371a08b576604936fffcb8381edc1d55d671c0bbbe027e0fb222f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5ade6f438880981ec1ba040bf141f051f52d9d6a3555a8dd34967f2bf0fa9988a0ec17d5b80eab454546fa5e888a69953e829903cbd21b25cddf3b061fd2f4a01d742cafe5dd36c3d5189545d97d5429d133a312;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fad5798716d83d4b0232e3ef60838c7ab55e10b06e11d6b0da16d69819186a7eb0cc299824a3a48e94620a37c3f5ef9314edb7d063423263f199ed91c6f7f2654b496ca4f1560ff1b18dda098d986cb8cbf31786;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1c98f1d9927293424ef3a33e8137f050b4b3ba8176fedc2bda4693f70fc98a9fcb85db5c3ead9acecc85a7b61b828aea0ced4338bb9eae7ae6f370a8cd54e81f381a4719f5476d36799835331ae31aee649f78dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f8570c963cb41ce98bfb1bb378e92663536168dd00f59bce3b82bac1d21272492321798b05ba04dd83d90c66ca7f58e560e22b0a961f447424a4276cd22725eb550fb95f17657f4feb3ebe633020ac098b298963;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ba9de67bd89ad6104c86932b6947161f622183fe4f0219c1c5e1ad545f644a833ee23d71fb783cabfb246949c36b972a18ee4d8cdfd1d711e5dc93dde63ffb19f5472f892557cb8c792e14106f9ad8273fd79fd3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd802637623bb26d54c9510cbf47f08379ef1d5c00cb762ab30670f02d8b444da2bd49e9739a68a00d0e5d01299b812bb0f770c766e60869e6a3e14ae56d4cabaaada88a1b3045bc9a8220e7732358c2d3b040623;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e6254b6c3b0b87b49656f7aebb1af2053b259b14e5aa1016618f914a2ba9fc898ee1cfc330e02327f5fa5130ca76187fbf4681a8bec08c6928f5975f9523718c816a0575101e5090d3013c29caa85c9e97e4d104;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd2c2941c14a194cf7a7f12902e0b50199d0488e9a40d7befc21754f46cc95dfdb3844caa1c1afaf6383f64f1e364e260544fb3d7620bb61824e208fdbecd36074b1a1d9b479df12f6ffe0a84afe6e3d3040bfbf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18577b8c6f248413b0202e1e7046ee94f4a1780fce3447e3e8dcb63345209644f80e4a02e88821565fde84e2b96550255d845322c82e57b6caa37807e3e30ee1bace212156037db47ae72f82a4efd7b024cfacf0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19d2c09332a55aaf44784fec20c6a25dd461be2f3872355b5f244c7988b6765d49c5c61766fe3041cdd00d33ae8ecfb55e365c4cd2202e1f3685b521846e7fba776f205793603487d24339191c18a3a329510db2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf67309027d4bb6855c998a2873ca7e23f456a0c76479b5a889f1000326646e66f27c88fe3822f053d7e8a8023ff3e088b7118a78523931bc8da3820ace8edfd11012fbd6092f4da0a435b60ea411b459569d257ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0da67178ec98c9209943173836021a7c14b9beb361732da699cf97171654ffc906ef003bb612e7b84f59a873cf84613c424d0d3a2de7896cc1f8c41343278f5641c5f68bb43046ff2544aedad1da3420669a7088;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ba7bc0b3778818ab97a6c860a99532b22bee9ceebde5ea367cd60485d0606afeba8e1b8a7cada1d004cd582332975a0e3f429986a798f226baf82dc3ca1272587e148aea5e30cf26e0d979f806939a927e089198;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ee06d535c0e7a7daac0fcbb43ad7bccf7f1f20a71bf57306cabb48f656e7cf6830902778ba608247d34e243b0e1d745bb1f849783f102dcfa22f311539f5d778f2656502d5c45fde9ce94c646f6a9133d74e398c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7274939e52018484e4e2124c3572aa52ebdbc857e4d9488be9f3225b32c6271d3ef8c1e611812167a68d46db0126bd211b2748a890da8dbff7f3e0d98264765e5c18e9cf204611782f1dc9b1a85babd3452eff18;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h255fe9b6b21543bcc694ba4ec763fda5c2afd3d2319fce3e025460de89205f129d47dd6e1767a54f5203e8b1caeaacc7e3a55631932359b72045263d57908bd454a912f140bfe69fe586ce4d124b38032196237d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77738467625688c270bb7f427597ad90ef616a02d4a26a1eec303fb3121852395f3bc4f0f65f89272ba46537b1097bdabfd8aecd82a6da88767a8dd918965dd4f58e5cbc3e52f96eda5029820a6fb9fb9a5387873;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd25f2734b5328b6b36f9acf8177ad33702a3c4c961b7b8fa97359ba62e28051573799ae22da4184e45c5093eb6c17d6a5957654f21af3e28d11141bc78e86c6adf9e801e3098a21cea43c56f287f76725d7a0497;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha814569e599adb83cd8a22c2a1c532e64fb607448a4e0bd969cc0352e22fc519791b344c773eb684f90ccde8dbfb0bd84172de3e9dbca162e9fd60ce57490e4c6f63fdd84cc6e10ef460aef4888765291832478a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb99b029b92f5274da58e24db974e1094822b5a8dd64ffea7be9e29595065f3eac31c925900ed51ebd090ad44301dfcf428490d35286787cf3318b2410253b9cda1b37739bb43a34256ce7e84094583497ba80f61e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdc7428bf883390e61836d6550850e175e48723aee3912065dcc080b588c9253a22c1654b451a9e9b1f59e88de5048e83b7085ad426571461fdc85cc36b73bb4125b37a1b51276bd0b4fe78a4b2943ed1ce3b5a82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf35381e0e1285d8f86c6df3da7287b73bb9425ce759d65a8518bbdecc67899b01ff179c0b99443666151826489a392b5718d772ecbf8d63859dd87beb239e0bae06ff902af5ebe68692dfed304a53e1b0e0b249b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbda5c15cc75d77d8fb9b2f6934d17000b71fac40ab37c3bddf4b108f159fdc2fb22c4aa031d2b21ba64beedac31a290faff3c52ced452b0c7120057df7304ac1d9f8653231b8b4393843d31c471906c6449f16654;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62bbf7cad3c4563e848c89106a841953a93c46ae61ded1c3346ea3cfc259b7e94cb59ec7f9d7b459712300051e4f649419cb64b7e1355ce431d1b93a15f2c9955dffcb14b2570f0cc1322f2ef7a2120fc06f145de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2adb94bee500c48bf364e705a8db7b6d09ce5799339f7be0ebb949003cf17c9c6594c5ddc1515f08b38d82d1f337fc0302ad374e192172e31299232d29960820efc3d1a4acc9248e138cfc0bb849217480990239;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h328e93b3cf174bc3602c2c952d86b5836d44f9b55112924fcde8cf335f80356669a53803006992e500d9f9ce30277381b46c9a1dcf225ccb9b92f0bf4d153797cecec0597b568d17eaeae1d47dcdc147e7a91c54f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1714cfa34fa325632d99270eb653b60fa8ca0a163bc7065f83adf76c070099e3e3ec57abb14e00f9eae6f90eaf4a0f796a0d433c40d5cee62cbda1779a08da9963390ea309b14293a8670ab5bb5a42a3eb3a55e3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h471b2da7f7519a143d5a26bcf6e1dfdf25a6bc2084caa4716ee3f826e9763e4e5217dc540d373a98701a325d4c6c422e7ab67666c326f328382881c68955a8b09382948f111be903235219b4592fe13c76456f174;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80868eb6758b03b59b148f12819ef1c93eaa6b956419f160c0b8395e1d05366b4fa75d9e3532c4560609dfa6fc05962176a74b36bc4205f5150bef1fa23c7d009c761e6b4530b756c5f935fa0527b3c0e1eef84b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a5b5165c2f0d517f905e624c4f4fceed82dbd6886c698f15beb346f370292679113847d11f86222bb1b2937cc157f688bc5f14a3c5865feab7f534179980fb6d875a4657ddf9c6668e234f2e54c99617cc1fec5e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54d633063608bde458f920ef0e1523f0c7de967beeef8635cad9839aae1fb2f3c1cffcb7138c7ea105406d8d5497083a2ec8867c86c07da49be612873500fa6e2c34b1ce3773f8fb364a324609b6325b0c42f7411;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9c04bc5b45f5597c45867abba1db157884af5ca22333ef3deaad4f4780be8c10055bb918c6689cfa268db84ce5a5c131b3cdd956dd9f85efdc838c01fa6f4b003f78fa682714febe2a32c15680de29a2636ae855;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479c32ea5dd6d7996a1c86e983cb933067ec00aacfc88b1a3574ebbef888f74e43fdae5dabdec2ca737eb0782ce7f9c4a083b27b5a6959df70b923c0489bff47a653915f080b7643a6ae6770321b89588b46f6283;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd680a0df690edc3b14cec27cf823a678e0a62860bbcd1587d34fea39dc80e41a0ac745216454e8f5dc59cb3df62026993e163bbe87b8070620b541740738615dd368cdcbc1e61bbe93d7f4710219eaef4a53a6134;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6df8f7d9f53bdeee8a34b93e229858d5fe62af59f9d0b2eaaa2685b3c68bd8d7b3b16d91873f90f16fcbaad67b2d3a73a595b56558b11bd40ee013e4a74d6a7fa1b74b790489eef9aef2c4c181fcc6cf50f0f3e2e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf728060abf5cf1433479e5bd7eb4b524e24b45feb2ae9b3689cc1a08931d4a78b121a409b5710947a4ee3752f94b6d81974f20af0b50ce3366d61405ccafe2ec1049ec85c689ee587731192a9e307fa0d974f0689;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafdd7b5bbed887bdb29e7ae142a7a54cb30be89be7b0575f84b9a15ee732da7c29fd8e60a4fdf68c022155a9ccf90ce76d15662ae041e5b1538587700c3922a5d9c8513387d03c224c7c546dc4422b180c50dd599;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2cd3e0a54593733262b1f4788f1ac2fe4246d8ef85e175ded7ea70793c662e9097a163a58efc84452d896acb7051db2ba9de8c739e93e3da62c86a4803793f76662a2506da9ec37b5efdd85f29e0a6bdbdd11441;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfb9b97dfa86e0cf32c4d0449f028793d01e90d9fcdc36762a16467c9ac1c81a2795b66207066465aac2a3bef6822eabf00aaf7d172ba978c26e55456abfa33981fc0a24def0fd505e701897b51fe3383bc8008ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22115099ae564465b624ec45f48c08da8c20ebcdca8d7c6cc70305b00e876d5e45a36d4ee9b8abb36b65682c4705b223d5a0215865e5ceeb06973b0c37dd83e19229ce22201397df0c638f8ce0184527208f9b4a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69fde0ca420b8fb7f9b1f64fd31dc87c59db7490012c8415fd0546cfbf30eace589d3596183ca272ce7e3a7cd312c2fb407545bf94e14914ecd97cdc8511cb525b4655690cb81fcb3d02804e8f7f9512cba6db306;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h671ee86070373012f9ae78f6f6ee4ac8f29f9baa6d30155f5598d13f106bb46fef00f209be71806430f4e98ad6438424807ad329b791140270c6be4a2e16fff9301794fad582306513e2787cb4b3589a6b0024f4a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f102023ac9deb0580a9eabf7ff252afea00eedd8474190e19df18ce64883419720d15ee5602e856f4672213bdaaf07596f85bd363bc0271780b2fc0484cd097d0112ab70b24ba2e7275d8bfe2a7afa45d1cbf84a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h363de8cd14c781cda899cb10397510bb2e9283904066264455294c18fee8024ef408c1a08816ddd85da489918bdeff756614c0bca1e021dd3641665e220f65c59ba5d07c5fe9cb63e419ad7b450a141e69f42b27a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71fed49ec376cc3ffb1b3f72dd197d7f313361d249d01f6ba735144e11ce0517028d86ea9d9ff918e0e251e41ad1452050ccb3228071ed8ab25d1329e648055b222c87bf50e55d57758fef58b6f8f53142cf7d4d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf38f1ef0b4e3ce196748654786dae3d4b86768b62d779c22a7abe8ba5d387508f73cf214623d1ab7b6910e3263fcb7fbebefa14e588b152456b32d9744594a4912d81d44730ec49ae9a5e70d2beb43a8ac44354e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65dc8ce888119027071d4d204063436de2315228da9c099c18b82d241f884feb5dcc7bc5e3efa69ab6b6cec556acdfdd86a80f5c87ab16f194c6c7a09b666a1cbafc0c549155406d4b7795adbfe6c6b1a7f84931f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee68ca32168c25734a04ffab0e5bc6e71a0a27e5a149591f708b6e7c1801e591db5ef5b82d5fb236a0bc151ceec71b677015212b8c0228031be727d6f2e07b66eb95b5a635c41c8ba72bffe489bdc66931147ca22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6063cb31ebc85d718f4b01c228df62a8bb4ca6cb70fa07073297485bce04ccbc474286f61f2a87650212c8b6356596771a5e52b8e842d13335b313210ce2916243864a5763fc35ffeab68382045fc6b8e14fbe330;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e1992eaf8b0d598eb3fb23ed9b759149e22d59f0b3f04515911115d8f501b5c8524f0087d671dd9f2f273c3e34ed0190b244ce9d4fbf985b1a393bab853d984461980128cb84f674f53dfc33a8779708ef699d74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1595caaa039456cd93e392f7bf4bb79b3c8b310e68b70720f6fd73038dd94e31de26a0767e023a9a084904d8cafd08ff8708456bd439d27c4d7ea4ec2571b8e4fb34fd2a4a8dea0407e75cec5b7fb340d1b890558;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd301e0da4dd4b85490d5a05be394ada2c51bd7c35e6b0dfe7dd767f6f7b6286f9c2fbceff4016a0e42ab475355d62d8c0ab9552b670d5da97e222dccdcf8447a7246c2db121e68b0d7d72570094a3e58dfd928833;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd19a9d24ef921b1e695167f66dbdd3a907b0371c6bced6d8db3fa9b5af26d610755a85aed9c310e9c8c7613b1ed6c5f4f813baecb6dcbeca2829e68fe1ab77356cb5ac9b35279db36a5f99583d309569037a6bd0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b1b2822c6b1e39a77c001703c24aa33028ccba39dd497b8d7008427543abb68523be6fce5a09b869ec1e46c148819eed946e5e0b8ec6073f7d8c986d6d711d7b3e4c6b2595932635bfd6a7a57097f6ff7f7fd668;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5e2aa5cea3d1571cdeb00b39fff58bc6b8a210f0e35c1e363f6f6c460afe053c83cf0d6c5d6441b2056d82bc2b93eda691f9092feec256305c7491a799f80ff718c21ff451e9f1e9fd77a6cf9780992b8e4674d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cd8722a865e0b2b240cb3302114884b0edeec860b732e5c11b633c27ed5d0ec2e7c4ccaec8bf0ffe5641e36ed16528f3f4c01b396266721eada842c5bc61558c77a43ba4321ebf8d2e913cf72bf1317ac598b30a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d1d1005debe4dc98286012ddb52644616c050696bed6742f227e4ee3b7d4388aee152069e77c9784b416d54c1c4100783c8b15b4f17b08cb25dbddafa743e11f5ccf653ade63c974e9c71673c74ef42e7206273f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ab0b9139182de6438beb9d3a8d1b44a1b939cf0e6015e6f846d925a1a7f5e1abb8d1839b9984401b70f15f55822c39abd9b06a39d3915b80ba9a73cfdaba2d8a58749ca0f4cfea79cdd17534f4a84b001b188bd1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec5cafdca3fcdbe0d8ddc3af9f5a2229671841a9218dae2a8eb0d9531ab934937cc7d8a787b0df64d84124b907d69706af8a8276f53b0678e2d1748d305658ade7615a993f418e719d3d6c76eb02cc4356e01d0b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79791bf0b48d27eeaf97ed46746f890f9dfb188b83cbe4893ecc97c4810a7bc850d8a01052dbd16ec8764ab695bee8479d2af729549258b69d68032ab66225636be140941c3efcb6c8a3216422b66ffd6c722d9f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h285477791cac4215967b483127d4214b8281bfbbd5277123ee5995897ff89d24daab61d72186e0b42fff6d10d83fad63cfb73776d3b7631b17d6473a7e6135e40bff58f4562f1680b2d93e4802aa83f2d71fa5aeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h208977089018a8005579d200366361eeeea5add4dc19310d0cb8665b1088a2f8cd5a05cf292165d76a4ec0795c2a2c89b2d420e9be2b7f03ec13d31783fada6d81229896d37983cf96a21823cc265aec1fad171df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h524f5f4af39602ea67c79376d2d5977b2d9a9d82a54fc5fe9b39397325e3970fb7ddf93be229d005078a3f9d155c69eea74fcc5e2608e4d777ebd996ebd3858dcab665dfc61518dab4ecedd95673370f79985941b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47d4ee8bbee1918b05a556a13e21d348d44f00a7339192b9b9c0b7ba1a23577e3fe5b8e61983fb369aa05dd6a889c344f0b25b50ed2701090c0e5b56eca2ad47379dbb5ce05e745c8e46cf11f3f82671fa71718ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h438bdacebc281acd91d4b8eb56971d26de1d4922196233385fafbea87ef67b479112cc8898ea3712c1a1106019d2269cc502089687e4c6633bf21a609f89be5eee7dc42ac08c1b30515ff59ee499703df65664bfb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800b113bc2ece5f146a3e7c6ea6f47adbb8df51433c99d3212bcb3ac83318445039089c27c802be4e57d50d39066e2bcf650a97f2b7220bdac8b8061d64b5fd115ee06a5452f866c734770f4a0e34d838a570b534;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24fb1d5093c62f6d63bcfe7a100f2f2035212de20e487446efa86c62333e6979747713fb1d317e1cfdb8c3d2fa7e70a6b65018b128e0f86bc1b81ba0e458bc74ba47245bd71b8e5060a446ad139a74c3f220b45d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h773e92859be964732e94f4025b0036ce10b1bd1633fbfe5fe070c0bdf2a193194177e8cacf2887b175ad123f87f4bedfd9525c8acbb8559711eba5a7aaa3f3c7d4567bea0e094bf31bcabdadd165bea2b8017ea97;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h169769fd1048ca8def376f2326e23f573ae9af126dbdbcea5085c0c315a8c3191a60d689597c3ba0597326062ba5f19def67e1806534792a05a41203b0923c830f9169271499e5cb738730c7bf939ab4483e6eaad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7499d5515a891ca21ca011643bfd3944f6459475379df134a2b1d3600ed11683d339a27a822476451ada832964b2eb6c9eb56f56bdfc5d7ee9cf8d04f86e7101f2177e7cedcb26aa26c3d1e92e7a3a5229946b7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82756f60054063e5617ab935ca6216f7fe5dc0a14580ea1b07571829ad95c41bf4ae3374b9326a241ef5fe7aea383af0642efec4515bec3414a16fd124332c3a59e4c1f96b94879100fe606e2643251d1ec3fe7b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8efa4e9f51bacc7b85678485a98a7e96e05c05fd5ab5c9e9b4ffa2061085036110bf2ebb76287d15a1aa044cc97714eeee9ced4c9608975604a435d86b5418c945c1408d2b52d5688f962c4e34425703fac836b23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf23711f0d35e6df548530b9c1ee9b975661f57d659eba536f4dd7b4cd24bf7639834536e10ae632d3b0e407ac6f83cd7c2a794cd30172c2a4dddc05e6764c799ab87752eb1c1eeb50cf460c0cc9dc4758e2671a6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16db9d975c8df031be5067373da9c63436ffdd72e633940b58acfc5f3d5b012c5ebd2748f4f796061e5fd3f60d7d3dfd7c4cf08ef7f06a8c78ae67bf0ac354bdaa0b8a09df7bf3d30167faf4d25bf7a6ab235f1eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had091492bfcca34dbe80632864f3a8ea8f1b0aecf1b37e63d977638f55da1a6acb7e374544c0815d2070818205aa6e76f15dad95badf20da71f5a89e6d98dffea1298d800eba955ba62f01e648625d78e31f06b38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc74a8f4d740dd1c64eafba00b7625d5a93f1b356afa06f4213573dd77a1f9b0a4cc2199882329b72cd60e94d2e6949e5ebff946d89b1902e83f4ed0dedfe958ae4b07099c130cd6a6c44c3d40616cc2275c57c9ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5afab03b4fb01e99b4bac663f39c6443c268a8908458c4768624a3704d8c6138a2859fc477db8f77a08fafba995e06576690705bd135d515674f30ecd0ea36b3dd289f05c957fe0373e0ade2150891249e011d088;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc86fc5ec523da84603fdcc628a644d54df97a8e37c01fbfba4f7cd0d7cb2ae3975061684cf194c4cf84ff6d78fe7dbf4ab96e386dc0f51b12b7ffe2fadba44aff99f3ba64a5e478f237dc32647c6444c9267f2adf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53217c7d875371200736747021e299f6ad19cc3e36e7f044b966182da0357cf0c494a463f78a75eab55fccff57ab9b27eea8dfdb0d6a3533d4f43b4c664a0931e9ca1247fe6352effd827a80487f5bd88ce5bdb3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e98d97c715e07af8522bf784f3f48bde9b6514c11584ca487c5c27e2dd004d541b6c4f028c25eee7751a45057c292c2262664f0f1bfa0d2f8de1922759384b9320cd7ef7a4a97c93a54c291f4f127d2e44f7a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26ac08ac630f0cac8bf570c4a30a92b706eb25f539d64e4c9285c8528b2540c966f11d2b5ad8eeb2cce5bc6dc56e3b065d70ad7ef78af15bc15666db99d613497d6b8e1d3d7e20f6439b19293959953983b8e0b24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f51ec60603dc8dad7091a6be8d8f1cebd4a492ca6cfcec825513b97ff3c64dc1d9bf8706ccd251cba9ec1967255f2cd89945c098689e1be30c031b24a2d540db15bcdec2a3410d6295dc709fb940e4fd4fd65529;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26df3d99c6b47df930c14243edac51d603501246e11b4766500a34ce9f1e189f2174a0e4aa736500f37bbe7239b5afa50a205470c8ec7bfb1076991ab26a0622ced26b429038e67fc4db1a92abff52483743ee450;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a222764e145d62d549b478ef2be0d19fececec3cf1b81b418e4bb698653ede2f8d8b95fb78c2052c3c55ffaec496102730f0f6b07f46e9d0f7d4165104736754290aca480e50fe8f3c1a670bf2591a1e2d5aa500;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb66999a1e1557a6b952cf0b881e8e0c29f0696ce223a2f7bfbef986f20d4cfe16fd6f8cf1ae3b7faa9edce27aa68f6b13e12edf7a31e0a75fe2bc93f29022796d43c71a1773e9b17ae00c5f185c91f784a6ac4934;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h693619a3594803b9ce750abd2ed7096d70e7635014155d188c51afc385d725c5fc53f7bcdf332249772fcfc422f324852e8c2ca5f64c6f008c8b6005fd30b4bae52e6206c04ff973588bfae145c9f40af4e5f6d0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4ca2a8ab8220510ada0dbd915287658cdaf001fbc5fd3a6d226903ef0d01e0416772644a76396dc2d4cdc2dd5a9170455e85383dec267fe289fc83e21bb6888948f404d13c392e75fd58dd8dfa604c897acfd8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1623e322b9e07585c2c8c488a8b47b702bbc303e7260ad3ec7cf404fa986db79237b2c029ac316d71007bb00360aa79626c81dc06142821acdb1e7e43088f2e00c7c0b07f695dd885d877cb1b6bbb126a8e5f4fc9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a015e1f21400a833ac2829e8549dac8a0d65d1644c6cbc5ae1b6330a42726079bd589897264720309b17b7a3eaa46fad76d0cd5fc50baf9a113cae636839f1cba7ada06e28534c5ef177856ebb4c7b1881264709;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h693cff5f28cd83e59d119f413915ddccc44581405f4948185d501155a836a81dcbbc3ae9861d7d8b4f4a0653bc8874d54e3c8cf6964fdc73f6f8969076ac4c5683ed663b907bce11659d515aabdde5e90f692a59e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6eb22b2822d34197f0e15441b68beb7033c73c4ca525787da0d049fff19a23c22461b5e9330aac89b13aef72d35f96a265e7814a722be47cf60b36163a36176c199bfe497f77d867fc45e1ff3f912e2ce6207045;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1a518ee2a45c13f9fb444c02d3fde2e4f9e6ad7589efe7bcb99f2ca69b42a669eff1823966a9c0da94c9d6210f65fc65aa1ca626566a8914c2c4f262b36195ad48e1bab98981c776c84ffb8318d6323b030ada77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3d5f1dfd14ef962562f38df57583ddffe4c5a42c197da3c44511794ec85a03b123644ad2604c553d1be23138b27dc106da8c617733e29d5e68902a52c23d9a45fea524188a9111696c2f3c81e6608bd1617be8c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb98eaa0ac2e864af64e59239e2d7b5bc9ec1e455a87c811199e845f5779717d22894737a88bccdff0879e34cccd973d49ccf91dc06a3ad1a2268ee25356b4cb55bd8fd7fd5540c2d45531dbfbb08e45a138397e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14d8878473eb3d3eb45364091dbfe4113a0bad7df7b4016717a8a96ee06aedcb610e6ee1bf71aa9382a200db4bac2b5109d65afcda6b4b8e3f68383572f66b3fe9f789bf04fccb85cf048c2408c10e06ef888ab3e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fe2f5c314c2b9b6622606116f6340af8213bef322a2900ed7cc5e10280f3c9a6acf5e9fb908e594527f26faf89daf72ccddcb9ada6666cdec62a24231830c40008f15fb17fa9fc016426212c680a33952e74c5f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53f555ba2f7fc76635c2c818c8464b3f3dbebec6ebdfcad55a4cd148e2b3c61fc60d3a47c9b422fc40eb3187ed7919d3e583781111346a8e1fe633cccc51aec656a626a821c7f59c0cb68c49036dae6ca5aa41232;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11dd039987f495cef09fbd7349eca2a54a8f2801566510faa50759925e1030a1cfa38b669b5f257bd620aa3244b378e5846667ddfe822d9c1f72e3c4aaefbec12aa6571e9ae3066ef97d34261b2b34a0cb0c4a030;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h187752bca3e2d928c2caa0e8aa10b3e5639feb3e7e260e64383e1ea1ec7dea81a7b03c26779d065405b40ea192ca139e4907c2512e6398bb37f1ac17487658927da6a9ece4e6da3b82233ad9d892d00d262169851;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e3653d6857a6f25ee38dd1cf1348c0de099aeaf98c569316bb0a4f15ffb6c6c8caf9fdc850374d793c7ce5e3047cd452c9bef7b42845f17e32437dfc749cd2eeedac75542cbada6de62dfd4fbd1696dcc4a9277;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb11f55d50c884425e1c17dfbf20ee2a787396592bc54e438873ca91d61b5087db9b9df9d9ab0a14293a1d9cf678fcb1bdc7a0004e86bbb74f58dd0d5dff1f8c405393554d415f7802a6acb13565cd0d74983c603;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fd95099ba80674a26ac058931533e3d0145ccd6958062b0effb47d47514f1245c98f5191d65491c1759d96510da84a23d0b47a13585cb123c1a56b98ef92bba3a0c93214881d999f529cfdbec8bfa100441b4554;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf140d4584128278db9c93a317a3817bf94a67fd3a74f17d143c3c6e020150ae354ecb0ba515f8e429f0ea800f6b0662201ab0075cef680e214e18399dd2f15c9927d77d8e6a52e587d29ced2d0342fc46ca951171;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a4c8df2402e68523e21e672f091cb128d9fb6811b641ab921a6e0a52c2db9105a687d5a1f89d52512ffa2aa1afcb4d016532cb9673fc052a624cc13cc4f5c58ac6695d0904533a9202c593503b934feecd5cfdfa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc56428ce0cc8c12185c838c042d2b548b653d781b3542ee815d039e072d61f068b30c3941073c3cecbf9119fd62c1b7ab96dd6111b1a173fc396ecc7597ab49b9e1cf7b43cdc59ac932c7277e82d3c08001406e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h308a0fd17aa353412d932f8d47060cc4f96bbfb18caee06265ae3657ef5a803125c433e17884c5f9085121e3abfc5895e994a3166c3aa10d182d1ce258783ce6f9badd1ed4c89154c2f573c7d54e45340512320f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb82b9ae0f0b986e127a8f60bf53d670aeb8be6dffa1898ab1bdb418bf5d6b7ab96fb992896ffa154709ae0ef0b74e4bcfab616eee72f9868b68f70efd402d31cb611a99bae4373058c1d37b31027f9c643ef2bba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46e82dc1975db7c845831efd5403740b689bb47ec4d896597e7b60f331d29451903c0b7d993ab8022755bab8fd60bae96e968a1ee30885c7c6778fa605eaea557f6a67587f5cd19a5025fd0159892ed33e1545549;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h594acbc2db2696b9e179046c46e0427a396fbcc9535e38001e50ab0a19ed4b58a5d9f329dee95287b80c2b338d692e043021231fae1f5cf1b60ea63b3a8f6fc4e419a0d18f737c6839f6f988c4049fba65b9a7ceb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4d15d2e17536662029a4e3de52410635d5ac14282c647d39616af9d61f90d96a03157b9a3de342ed00726c695b8631e1bc8638207e207c365b321a802697d2d3d251f70511edcc7e53728cbbd2a0c891ddf3610a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa3f5b7bed974d80da6a1e80d119d12184f8a1d3c2b27dfae8d2d3ef18504da503b82fa14c9bbfc48b2a820397ca2a3b0a08a75c37a96ffa49d637a61492063695793bca9c28dddfdaf08e6ba50ef38f09cc77697;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c55804e0daca62245083cb15710f6da37da9495cab7809e9be9916ba50c8ed51b25c63824a7ab20f422c0af2940d79026d9c642b0a4a39a77ecbc6fd56bed70b43bdab841e04079a3e6b5648408b6278b0687c3e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf5fef2a51dc86b0796f4132ca1afd34b9afa2bbb6b999601d9d5c4b5223a1756492b945084524a8d70c7ed91b2950d43a7525059a1689926f0db5393d36f9736ae8feadf6d9b5d592b36986c1def2f3c74642594;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9168c930ad95bb6a56bf4d6e0f05834eb48c0718b3bd78bdf5cf7d08169de9eb2fbee1af1b60ffecd9241a2ee6f52454933d6b477673fe9fe8b001f6cf8a4ae38b63415d5e35c5c4871615c5216d8e9ebb8b0663;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf4084a3de54a455c04f0e23a387e36dff7299f11c76a4b98af1feb62d55428ec6bdce100ecb763d8eedf889820cbe6893d816db2ee08d92db78d86e0481adbc9b5c218b16681d608703faab5230f3e2a4104f963;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5ccc2eb46675af3360799cf5f61105321c554129b0e2408259cc37939ce6eaa494031f91905f37d9c95d20ad86c96ca4ec8b9954b6d6018aaa5895e753b97892c5dd13f9753bb3878d9c9f227bdeb83471dd9ac6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51c25ceabb47c0e972675014549808f648b43ea1221b441c563922a9561e4356f6b7faa4f8dc988960fa994b282b7dd9a070ffd56beedd725856167328704640ca50ae37434543ec11e76c222fdfaefc36b2efea8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa4ccbf0da5b6f71ac06649bd01cd2e9590c2aa150e379538f6f52b513894aef5f82c373a702f41a04ce9aa295e9198eb6c8652da6fc5069142b8d907769cd3d333db7300ca53a5de2852d69d6c9165c0dc540b4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h817ec962b71ab3e49ccc4b796847c47ec77493c01483ce1c6162bf888a452ddea98a12e59675f4626c288969ff70c5aafa76ee675f6da0283b24244b9ed8d1e382826902b914479e40eb53a6ddce5aa0b0708c575;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72b53c02889111265570245b5e286ae9b7aa5b364d46f7d499a2da8e6242ab1606803407116d4ee9c5b4a021fc8d14233751c1a942c7184828cd68ef3079f16749352dfabadfb2aa3708c5458047bbb35280f5f7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c275920e405388bc5db6a8519bd070351e3d2414d1dd4e3d69bcae394fe8ac22f64f3cc44fd2212420dc1aab0eced8851fd62caa95edae828a237f5be5657e2b106da200d278ff97289b458d0d19848096ffa338;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65c3c3ea7c42df919c178568700c11c8379e24b273e01335ccd30941f975bb3fe5c187ed5465f148b913224f09f73ac8184ede327200d22ffeeb5d759ae5147d03a1738c7c9ede721a2de62cf40737ed9fbec8936;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd24625df11cb2d7923831280b08ffd47f5f45839a7c43f566b9d99573f1f8b26acfa2d8f5cf88b4aaf1c4dad326c2fbf34b1ec42b72b99b9a3f2cecbe7264d1a395057c63e025bfd484b769019bd201fcbcd74283;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bfc6215c635aff9183d8ca01c770b028a7d448c29df49a7165ed5d0258da82f372347d5d65225a69773e8350b26af193ad6f08fe567025d72ded705ea222e701cda51e9b9299ef0132c361761e8c24dd7646496b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72a00679f4882bb9ebbf3ade22eacd99aa1e015dd5f7b41940ccf2eefb0e739c79a258375740947e1c3cbb1049500bb1f0eec6eff5cd61ae57f29a17a2c91d1db565a80081a9f34d836f34fcfc9ae09817612d6d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c66bc085868ae89aa294f9ff1ff5cb52ca85ba17d89aa3f03d0f0dac55a68ad5b2460e9175c6cbaba63af28c2246e7803e6fda01cc4cd666402234d47ff10d4a8ca324c2eada035363514d36a3a5cc380cbf24c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfedf7b49dbdcbd4920dee3dbd2797de99bdb4de7c01856184de71d8e93c1df4664c56fac8b56dbeffe34b9bee75fbb8f32beee29b806e568547af936ff961c0504f43cf8e5fa444870c4e0089ad2cbdf8f460a10b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5690597867f9c6c2a64738b1da6e64ba6fc8c5575efb1391f10dc81a957def81b8cf94845d570cbdd100e476e3ba88764083d88223d241b0cfe78c7398d2b60ca2aa9a190b031e347bacd51b646d07604ecec41dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1faeb5ba45cbe201b9c0c59a39069f328089173d1788790334e6ec49caf93bb7f071ed62743f058709dfd866f552abfbda3a12a259e926b0caa881e30396862403bb887e37573a825208b87ca3b87e5546478e033;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0c6f49488f97c426e59f602b215f7e895e3e69d00882d545de035a7c033e07d80335271166844dc59818f43b48a119ef323790d51dde58de3d100e074e020ddd95175a5952d54b42f2c29726115947e203b16f2f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7340aa14d3ff2a7566d041776ef98992fbb8172be581384845ceb9d20604dba15b3836e236cc92b13fd14fdbdc6ae8e636a626905e89f939c53ec922f7887e6b99ab137ea7b6da130c819a5870a75b06e510889;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41ef1ca44b1593df6399b5dfe717bed6cdb517c233b74fb580c8e1312645c56d4d57bbdd6e868d471185bf3e2e9951cac1616934090749721d6c8379067532c1b1ed1b3d7f7b443c833b79cd4f2872590c0905130;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f599849b49efdb9d771eea106add09dc7b4040c0c9d58ab5be3b2187b6131a414d200d2e8d9560d24eeecf019212058a2e0b1e05540f60485f8b03ee8dc7bd3bb7af49b5092c3c775c2c2ef94c2673f37862937b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbee32f5eee5c91e48b1a62a8f3cdcf9a7999b4ce3389548b3c10fca9064f5172bcc7f0ee8c6362a7062b9c588fc382f694660e0c0ad914bd372addbb6102108fe07b5c58a1d70dcd0418d3e36576c216767e255bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h374866cddd1527fd2f314be14803a65feee7e2361b6aba5b57b1d30ccf3373d798f3b2d66c9e190ee3a8a33299b02624cc72d9302314792b198b1f57496b3cce328b04cdcbe9f3422691d17beee6d4bc60f7fc119;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e91df6cc6058918b0c057d6a5ac86c85e40f4da81472ddfef9360bf646fdb1173cb6071eb808870d7814b29eed0331af34f1cc3f13d98e4473b1579f46ff35b2e00734d19b4160e12f163b0b2e6ffbfc4e3c2ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c47a1866b02c5f5f7698809b836932c61d607f302e2d822cef1228607b172e6df0b06ba40457df5d9b65f0c9bd7048f5ec1a368819efac8de4049991967d9f798559913eb865d94710818e827cc22165ae3707c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcdcbf0854dbccd0591a51b494177c56236f1c2bbcf22f45a68715f1398fad4ba10fde037fc6d218a129485b66796336f0172a2067a9129a87c7b485fc2e417e87ff33b742965a6f7004d407f3c2a92ec49ec155e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6ebda39caa5aeda43eb9d67afecc6156094c60d36d18cd1fee3c99305aa05f93c6df6c10c9181e6fdb5d71397393e1ee3596bf4eafecf23d03fc3355d88b3f01f84bab29f468e4abea5eed445099300d63c9e521;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdba831893e878c05ce6463f827c4ba423351c819506439a95cc07d0fce397b60bc86298993216804a7502202598491338ca16da8275d6c7f47c32726b00875ea1faec67cb9dc8b72fdd8d0a610e92a751f6036dfb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23e1443e45362f9fa950e0b4a014ee15ca9d0f95776c6307a495d9e190559047afb7b0253f8a4ac9dcf345af480e4551fdfe5a8c02124ed63e9efd031e6a150a5245199092427279375983ee48ae9858cfadf28df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefb44fd32cda421819f3de862eea4874937e9245772bacd676bc6118ef58029c2fd92f1d2dac48f55fbbfd995b6e4111b9274266f2d3a267cbc40f85e0acb53a04c6b143ffcfe5c317bfe35fb4f82af3be373f79d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf0de4b434141d5f605c2bf33220bc04648757e58103fca65a44300d376a27fe2346ed54e54adca0c3eeed322e2961d84fff8e5811835bea8e9770ae60ca2b71f3f4081519fa686f91bc0fb7b2c759aae0622620d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8318db6fcafc58431fc0b44ab24710d239dbdba3b33705702ee976d662bc61cfae0965136d5a35c687071867673be8be34522fbae058e69a216643df2cae5402a4e6b4af9138d2a1ffe090a5c49cc944e443c4db1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6164dae5d0e14ca3e9d7b6f041599eee7a4fc1e2e725a30695bedca2834fa3649fe03c16501dc9111ac58449876c954e199d125527ddb8156b5e086c0049c55012017de74190be7db6e7ec5ae685baf91c43fa9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf22cbf8e91dd62a7774ce9b2513af19841c9958ce82c21056659e2691587f7f8ce280d9cbbbf394cd8fb3e3f64e9ef244d6774297fcda3ea0f65fea32556583d98361db02bc6463e6273ee39fe5b4f0931c6b7c60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4256b2cccf94811624ca617c1d2030196b9abf59d7a8e9cfc550132ee58d2fc6c67dabf17a813b419b5b73e86c310d367318ca816f95f9e7dcf2195cdbf660b01c1b26e39f8a2c426cfcf207f1fbf17a92ce729a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75f02bf28a12a33e5f7120ef832c847bf025674b39c143679bc6d8892c33b8b7311a36ffa344a243c6ca07d6f45a08c9a301d4400ff7eb7629eab4a596fb2462f34187e17238691c129c345788cbd3abc1dd56a7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h303a6c45b04f1dfaddbc56a6928a236a6eb76023f73469ec7e3fea90d6a085a153a5a1c233c608f71eb1227c148d8d3dd481b23de12bb1dac8713818bc08a13a1e7e2b4641d90970ce93503fc30cb4b7f8c50d457;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd57850bbe2db160965e05d4600b2c75d8332fc8abb6a8fee5e7e5826ec6f3e0d63df9790cdfa9c93a8b64d4bab6a42a28e05312ffd517e1d6a2ea5734a82713756f4d5014010fbcd0942eb012e5f5807b110b09bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h786c4d16db836e5b71dca850e11eded5143131ecb458db8688290608e5b58f1b68a4df07d316f9e5810265a818aa4d86710dd040ca7de7d6c6537b6c4a622f83ba2bfa79525222c53afc370fdda429f19bfc96e24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17d719564199b901588d4cc7564fa9bbf834e59884b6a7a4705a46d80df91f7ff0527e46e417c8a3b7feebbd1bd8578dc83d52ccf14b929f2437aa042fccf49c8ef569950ef97d176347ac379ad7242646cb772fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21d081c9dc81adccff45bdf5993ba468ee2a4df5c94f0b744bb843b9e111bdda0ff8601a8e76a0f4c7c1b23349f9cad6d567b7371649d83f65acc08c07e4ba36d20b344a8d2acc820bb8545e5f81d87db4e82bff7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc3d33c7ac3674f3ff662788d79aae43151895b5c128914ef08653e3d25de7fd3a29f8f9d2c7ae5b93ebc38363c240888f4dd0bea742d359da5ab92d639703e8ec414993466586a2c989691ebb22510c71d9cdb8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc1c4927432464d63448db16a2478c082beb4a742192806a32c75631d24afde7b36f1c535c863ca10b780f776ffa3c60400347fd72a55822284d00e1251cbebf7aedbb2f9553f3408518d2ad21f51c0651b4b6d43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31e48fe3f122cfc39874cbd160291cde6b2faf27a3ad918a1cb3b18c03d994dddb95ac4d5c73eabaa3a993ef6be9f48523dbabbe209cd7557dd26e5ca002247b833645934d631a8426176b7db805e6adbc1c75f7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h868fee20c92fdb43368128a768f8e81f463a820511aa6fd130bc80a75fb8219bbe80ff369f6cf5a19f14b49532231263d4cbf1fe0a4c57cbb385a1e965e7c1d587410edb611c730a59e636a256b99cf6ffbfeac68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20503eed2e811c879ca53ac6250e984c6215183e423c59d51074677a609a843caadd8033d3123182a380c629780a413452b2ce0b05c22e85d59475170b9b5a79f7fff1b7173897c0bafa16846d28bce603e975378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86013ef1b7e3aa685450a637cbab50bb06f9fc8b3abdaae6466f6eef68908fb10283dc4edc3df82ffa1c3f95f27406be91f7523885e32efce2de682f402990c79a4a76b8fcf1ab3ffe5afdc6cb74eb40d56915a8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had38b4d21165160bc81ef925b751aefb67046d26220546160eae03f27f8684d3c8934f5bac9ab87cd80b8edd430e4491813277375abfc264063e9a58c0a99e7d7ff789de60077d7006e29b607585de4ed39c40a7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7533f8346774d2e18a997919534c723911bd4c3b179faaa84c904204d05a750b9618c392c7bedf28963a6d9995c26ecae024a7aa215aaaf73be32e14caf417c93e4d04269592fed4412bcde7e667e3c3f1d5fa70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20b9c40c0c8308996de1d9b45f5990b9608436f21ba7cafe5cf9a88e5ef53a05ad3772aed7dcd1be2b11117504857a42da3086048b703b121fe37a4b446f50768f6f5f869c7b356dff880c91b0702a6f1a37d27fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7370526228fda36443702fb07f4270dcdc4affe5a224539f60213ca61dab559d8abf2844e8af8384765ec79687002ba26f8c5275d19f74341bc3684e45264b66555c4ee5125841ee0716d30b244033c772e712a79;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88f00bbd7e04d5d26529cac2162f77eb0f9378e3f51c8674038563667e6e38f03e40fd005b994712ad8afd797bd14b87b504eec6c34e9e5d417897c94331e77006a5e2a2a45a5be82cc5aaa61a688687e04575d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a6b9b9547708280d1bbaea7426f37129acfe421fb619c52bc9dee5ff85aabcd9dc2e24050a174f20eb90bcac88ee875b0019001117fbe2a1278c8c01f126f1f5ac144c5c56a663324efdf2fabfc8dbd6ebf56db7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7332d62f17a34fc8ce47669dc5b7e6471aea89c09e9fe40b4b5d92bba55f8de0f2c36a06ac80bac91e38bad52628da26afbf966a77996d4471179bd89735fa8091e28bdc579d89a3baeca29638082ac96db15f04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb171842d4f0fcba99afd08172b1345019ca693b2aafb6af7cc7e9d7292f3a9731441dd5dfb5fc1d97d4389f56d3cd052469c1203cb35f35c32ef320b3974b7624163a8002874ce5ca8a93498d2e1df75c426c49a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1db7904c15ff18040a8c11af8b17ef189531623c6b3c8114c5320459cd519a3240fa917e1e074cffb1df21e14e5a80d1891cb6fe33fbbec0350c67e93cb9cb82837efa59e33c1ae71f5103dfc7cdceb97fe27d7e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5898ae425b398877cba294d6fa91f9f6bfc525c8f51034d52495fb9b377ead01a130635af5816c10f0489b9be364351ee815852a3ac08f08b34de8d26cded25cf2aca1f1ad547bb10e1a6f0284ef236288e7a6c88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65b1c73584a5e17480a02be83fb692424e3cd23d385d5d9606c9930a670c3f64a938c24cb076b0727f7111b827b7740c8dd2260c24f706efa7a71b06fdfcbbe27130c9920876afd63b1ac91aa4db814245e59efcb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e7b07f0f409f866b424561d08feebdeea0d73064443f34c2dcf636222e5a3ccc91d881cca75ffd66a179359a1901b38bf9c716e515d5d634af4c89a2638ee80108edcb87db8c3398e6400335b7813cd50c688199;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87d952bc29f5af0b99a7dc4cf0daf8c1ac73b3fe94896b743d3d275404d9da20b557a106ff9c045fc7a3341c2944d2350bc2dc7755ad66f618265e5477a2fecda9176b3fca601d481b3650d32a03fbf620d1e6912;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17f3426e34ceab420b8d12d6c4a11bc95867bb284694fee2bec2f41437e3c53c2f3b15bd8ecec3758ef690faa30c29d03148fec09c1d21a7b1b46e1d104c96b955e8cbd68a2382f853311c55c06bb6256ed767203;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b09ec9e395890f4b184a0308531311bf1788c47311a6a3d3a7c5451de0d8d79defe00ebcaca8f4eddc2c9ee77368a805f9826ce024b78744d0decfede3f2b299b6aa7eb7b394bd99c93efb88b88c6991ea5b48a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e0ddceb4c506ad400505641808fda85193f6b7e1882d2caa0c5446769f9740f1a17c43701b839bfb756d076cefb96260fe61ad26e4a4fd724b8af419abc40febedc74c61993c43adc7386fb8f1daed16804335fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1f186f7c7cc11865c20a749bae9b8947cd3925e058f1675e7e91cfb2b0452f3b001a4d0370c581cc35d90df9d22ebe053690edcd380697583c21205afe99a8fa6915a9e89c5d124f86e46214c56ae29dcd846d01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d10e0276b7ebfdcf9b2e6e58c9d8b4be2a443d7c9b7b82091854f9e685d675800523759d5c951d7d54483bd08e213ff8b83084b9c9379bb545afc29de895d27a521aaa54dde9736df628a86ace894f90280389aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5676dae6013c36df1b1f56cba704e459cd87d773514fb5ffedd863435d1efb0dcb85dd0ded31b6eb5834a43b855b4b87737ac8f968dd68128ced8d7bb9785ccdc831ccee5e7293d7b1dc8fa32140b04b411536846;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66c485c3b4a7dfafc9f9b2e2bfb5da11a6f482bb083d8d5b0ed10a49c1b97cbfd3752380048c17cb7ffc406cfdd4a9b32561d0d1765eb64fde3e57cd6a2dfba75fe3249c878b92b672c70b5ac36c0b4e60ab2294e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he600678b29f2b5453bf6d41d68e1725e200c095e42d0b529568849b795b9763c48f127f72b57b1d258c52a365f59208c52072bb15f9bf27218af9d964ddcc863770ed67fbf54964c54f9cb7acab8a3730035e9634;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h642cd54b82893d8ecfcd4366c4bc824e5da19a55eb69c12bb5f8c0f04d65745d470b697e40820b9c6c004d5c8e82aa7d97288e05bba36bd0187270524161a00866c6480b9e51bd5c57a043d92bbe1e60f54eee6f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h615262073453532107944eb6c5f598cb31d172dec760866a9534fa103eb73c10a695d11f9ba77b3dc4c54ceb27dbaa8ab0ec361f211fd892a2c1e4d547d0b958f18aff75b3fad8eb371843b3e8fc380e221865975;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4084fca959208355a9a198f2b3abe6c949acd53723c01a115a149712b17dd3a5359ba0e198d2461a39a6f694e946a546767517b0bd59f192169a16be8f63fb5686217bee6970609776d335ce6580f776d9c08f937;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11650e6b57ab29669adfc176b280766ccdf700de6ca83e12f154d8c00766ddad2a27d985a9153b26c7780096be1e8bfbd0a010d1a3e25896f0c81defc1ea1fc4e82906e19c8c39399e3ba6901538c8a89ccdc6067;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd9425799e9ee1f43ded05e404e200d19647543505fb2d077b27f9b48c1bff619dd2806fbcdd92ab7ab9db0b8d23ba1e7014f04a64a0e52035cea58b4440e46dd989575a10abb216914f613bfb9a2f7aa56a78d99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88c21c92dd7068055308c84bc471cdea553ea030cba43b66a9bfc2c9303b54978de82a7186182df575c1650b2400727007cabe74eaa054d86997aa02425d19385d3f0ae1abca2b924b4329915e5a857e5c9b7da44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd3328ade459367cbf578f63b673a7d75051cc3db54a74b00f2c48c54d2d6d25a621b8840b1bb5cd4bb249cbf2c7e51c95c3e11de8a08fcdd7e5cf49a948befd82ae6049406a969bc4ed3ed83b4a43cdc042410c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h629b0b765b5b1beacb293e1c0a536526a9c8ce35c499e6b7e0775acb2c3b1e9c4fc1e136609b4fe6fb2c7ceba633d8f88e2259f03e66b76054110961b5c40dda2dad3bc3e506df67feded2c48f014511dd92ec082;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dfad4dd665af835962defc8543b8547caae4a05babcb252bb0a349189fb3e37e014d099d70c17e0c1847b3f3f2bfa139e628c3d4e7d600268b1b0d93f10cf968841f6ab54031673cbd3770483dd5862955dcc085;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e290e3b111f3f37b823e2509549255615b2cf5cb3cfe9d988f989dec0f48c86ecac857fa4a13ccaf8e7e99d3686ef62bf77f4edfc89b830f7a7b23aaa8da1a57ef701fc403ab7fbbdcaa96172813791ac5e59238;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h259103d358f4b7e257f9f20b75daad480726cfcd9210b02d2b2d40b536a514df20cf2161fc8a74dc2fe2ed6933ef68dc41ee8db0d0a55e7c6eef84efad7b2ce103acf709ce3ead7eb2fcaae0f100a49a6783cf8f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7e1ab845fe0bef1ed8b064d7076b4fe5e237d605e68270c1a4db68e048ae6e52deb92901bccad70d8a212d93775db986a6d1e37337f3a810658f575739e41bd820cf0c25deab872518cf3cdf3898cb2bd9f35fc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9641b8f8a20763112a65fc45f000fafa339a772db9c4b861860d13fb679f5d0846dd691db1a87ffc6e9a6b831e6c5c9bdf6f6e382713abe1f40e493196c47fb7a201c12a090c22dbb4b325aa36cd4a0d20a90ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32f710afb0b86023e48f0072abad2d643635fbb7747d7d4da55a8871aa7ae48b129b610289e520d2e81f1e10169cc6c90d26d582c6d71aebd8f3076aab88e4acac71d1969fd5c588a53ead0777a624bccdb7592ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaae82d6a0ce460254e6f25375f3b50edd118907c8edf070529aa2a36981d43f1909c4895127bd3e89343599bd01d8233ee4ecb9f8dc299800c0b7a94f7cd17cc20cad78868abaa83a12c239e6eca9e5dd9c93d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74ed3fad0d23fd5de4f34d54eb53a100d2c664c959cc5f98c56ec076b4cec71ed8e7ae7a3150619f42e810f5c2f74bcfd77e0d8c8fb4ff665fd88c08d70219022b30a603f31d39cf8125a1a2c1084b3754599cb08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h706fadeb873bcc9213ae45d357a3cd533cfb27ef5dd255c8b1f401f0cfbc2c0823e3fb6f3d270ba2a2022c4d1430b153f14a5b136dc052c98cf1f5864164ed5f9759b4621ad01cbe0076bb5c1c9ea347c36ebb0c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd724f3dc8b5fb0acfe5d4aae39c500f1cbd0181b35fffa9d0bda5ec26d0dbb8a2a77d3d11d92496e76d513f77bcc7a6fbfb02bb8dfcad3b1838d614177a36b739ee156a5fc474abe8a213d5a51ae38e5f6bd59fa2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he39d20ae1cc337bd32c3a15593680be5b129ffd23a04dd237aff1c522bf2e7b303ee0357776be2d7e5ac8df41c525e723eaa418dc304951ecc08456274d6355c96f68da3b39cb4b234d252317af8e41c2da85d440;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc19e38c295523ec9f616b23aa1c9dafdbc1c6ec1e1cef27fa9d49e879170a71ddd862b7df4bdfa9c7ec0f96931b6098b38952c847b135211385b62cb0d4dcbe505c2a949d7c533abdb32b9987f9d20c567ee5e931;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h592b8989074dceed705177fe00620a683a35305259cf0a2b31dfe42c4b656a2f3b4a6ee3c78723173e04f2daeb36faefeaf137bd0097435e4c849ba29efdbcb42cc7a522403c5dd78de1578a9dd9061755e5d612d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d3d2205cca3322b8fcf273d197abeeb58d1537cc2343ee55087c868ddb2e0ea6502fd989507a6e2bff4058cef8763ef43582a409ff44093b4fdca5195762ab8d1ea21c6d28d639a4abdefa06c3625a3ed0ea299b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h962b0d21df87d3676eccb6e96ebdc9835b60706f587d4a591ced92f2566d9f8e14fa812b8afa7d11430f1a69aea5925880fd2e63ccd9a5249baaf9a41a00b8f69baa04aea8b9f24b7ef419d44d87d156ed9270b4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3a025fb4576c702b5dea6acce91baf2fa6eae68cc8013064564aa909a2f27f4fd8ce16103864143d6ea33a4f3f7227ca68f6e9526130a856619b126a6485524e554d6c51ffa31579d6d71e09e9b528421932ff5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24d8c869968688af214c789bb7dde46f0e70646b221f4c572d10e6fda6f029165d7cdb752d50250db506b3e9bf311cc2ca5c9a5754a0d758b30ed6fa8a3099c57cb7ca7a1bd0e7e4836c5f11e2f725d05c7a649e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he58f3afaae2d187007d016b3fd239a5f9f6ff282a24071060871e36d59ff2ff98458d08cb599c8435694e0c65cd85eb6647361660289e63af8f34d9401d44e244e5801ff7d505cb4fb82255e56191def1101eae61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eeff01ae138f9abffc67c1ba9c0ea35092e4c2387fb94224c72cacd7151bccfb50273d85259f4060de4add845a9db7691690b9cd00ade5168bad25c5df26e20f0a86027a62c978f67faa74dde78aa1fb19cb22b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7148ea6927f1197f85c69d1fee60324832424e2d671a8380c8e18c61e961514e0812c3a7d214d7a767e3c5cbffef272dd7e76b536ea61a917a5f928dd2ea4829ba5900e35c1316568c07b434558494cb9c10e590;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h685f112a2828e3ce2c12cc6fb837e9cc62673d7729bb76e19091fe5a4de5a4ea97c7a7e452bb8ce3b4baf8b9d162c9878468ea96f2ff40423588fa8b0235b49bb119edaf5f84c05cfd9b9c3194510923febb88dca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e3cf926355bd4dc6edb55e255f21652da48cbdee210a6674431591fbcedac4407e6f4be43bf373b6be387d272e8d5e8ba0a64751c1a978b27b0d94ebd57dde4f24007cba30fbe76e764ccc66d0a39c132a81b9b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7a7f427b36f24a0b92ac1ad62decbddcaa8b063fd0198d19ac5bfbda1759522a1ec4e8f69739884fed42fb80ddd2910d0bf55eecfeedc8c01d49197df5db29c96b6e2a79070ffe6992e6a83a3b965795bcffb234;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6893a5020fccbf5edcb37b09a674756accf3d9f55046aee798f66ab7244b09c6f39e545d6ed5a7a7135df6abc6fd3acb625450cb6aa6193f7bdf7449be30ce6bf9d41b3dd2bd0d81c8e24b3dee3b5c09cb12a521e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7057c3868cc53f08c0f4d498c77b07d8bc9f0634736f331e853cbf255a86019bbd579572a3e324f3e5fe7a6bb1759e65ef545d19119bb6baf7ae2cdb19a0f47908ec966dd9b0dc229d9ee1841e87baf36d41e91bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he49315dce256964a60743c92dd99d9728acc645778c5e62e8f12835a2659c9577edc1085c24ad3a40cc2dde3f3b6e76030a559cbe05ea5f6e06cd6fc23012f4d01fe1f6d6fd6e07042af276ae8ba283d5e1db5b61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18c1f734705c50cd6b1c10e7a97defb4d035c4709c416202a5a6395c16b01cb6433615d85929250f01c5eef3ee516b338a46b9b24e871686bf4ccc64ce122d9d554ff6d981ce6cb626f72a2f8c3bf73c301a2bc8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h259ca2fbd8919d33c4288a20b8f9c81aa2c3e5a3ac55e41d3368c6f4ac61808afbdd559c4965164fea238f02fdbf75b783929852f190febaa3cb61019db368d44e743e8504abfca22e066708f059844a2b457764;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bd555ddf10196d0048147a978728425c91de4f73f3864c048537f5c3b8f652e5754ab6ce2503b0090057777e240a24f077539d1ef720e653cd11d02cfaeaa27806202b7018834dad08007819a510ba49f631731f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd11a22b5b885a516821634d6db46783e1aba58c2075d718e5d395d107712e26e22a05088a9bb54e61f138aae7f6678059ada9a685c45c5608613a8445b3987abe5f6b55689f5f22bb2f1e06e0a46e0dd758816ad1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d7610740b49b5fb4b7d818acd157073d2eeb6adf04957be6a7fac2232e2c850a896f9c829e0fe11ff94cd86fab69443afd5b01d3e527436460e28a7b66a60e5da051ac33a2b22ce9c2ed187bfbbfb86eaa635dc9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba885c337271433bb784658d8dd921e5356025d2e06d97d63923ff300a09f3badcc6c56a7594bfe1da500f8b2b07036e6ad23b1f81b8857db3ae4d1ad48615c2a384aadd4b89e07c81fc05fc0ebdfa909c9262fd8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30e8e6cb3469696c307769d8ddedeb23e6f433da73099f8625d08b7aac519e87d85067a84cb616ea18a0deaefe8873fdbb33fab8ae5a6add5c88036c094732f41a0caf25965a305940b19a20b6164b4289c93476e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f2f40e74afa45cdb0818701d49bc32e5fba0610d3c928518ae8e1af93c5666a61232943e6938f52050737498ac37b01384cb730bd7155536b1f79f84bfd88dd7387599a169050c37d913e394b36bb6adbeaedd4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98d85b5eff6ffa830cdbcdc7ff3c7f9c13967ecd6e7bfd901a2adfd37beb0e7a3f69df69b8bcf07bbac72409839e6b6490cf83a7af75d38c5c39e45bfd7803c547f0c1c4305001fe9fdb2971f734825bfb8439205;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88f1c75e102bad4da0b505629305f03329b3dc2540b7f113f0a4d5e3cd6fb08ce4f85a6d5f122d63c5b1b7f253ae2a71decf2ad037749e3fc78ec09cb6a2b0401a8e64c582afd95bc7e4cdfa57f23d285e030968c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4faf870bba9d814ab3f094611345a0f8a1e55d9fbb7951af5c6e17d2bfc6df37e7feea4e89bd90dc76b09761688eb43ca9dc80fd98400a2dead58b98122dea5cbdce9adc350aa6be2832d5928ed83da176e6b173;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcca881589e0be66194c803dbc913568c86915de94bdeec7a0d75135ef7e53d6b6063726c3a3b1a1242d1f01f84ee420d911b8001c0f18dcce65992218f62ffed745875c7f326ecbbfd4f934c35ec0b2c7b0a3b0c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5140cc4d9a773dfb73e2b488727840bb5791530f8dd2417674f7a3278c38e858d13bfc9034259450f79e7e351fb3e63fde89744aec8613ffe7e1b9b2d73e6dfed35198be995e598ff7da66673c761a0059da4fcc4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h392b1fbecb6f4e187304abe4e5629fcf2c9d1d51a286533a9cd543785cabb2e13d6f38e69a73970b1dc608a4cb3bd6cd181c374dc60ffe5f9ca4d629db6820c04fa8cc76982f35be0339fbdf3fbf84abfcc4c44b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7fd4cd156a7eb3ec459995cf3a3fc05dec29db076697429b1c367241f2515e791b37b99db7eb40cd468f97609260a01b66679bedfc420ff97eccda5e8d68684b91e5d242c5bc4f9bb57708e665046410055c1ac1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6f1bac573309f46a344492913648712bef589be4da74839feb6dbb0487c1747240060a7fd9faddccd94b29a13b5cc371be4c0408b2414a9ac243ef1580d01af7f38d1e55aa7d796f4be70c704b0b79f40a4d84c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c9acf2cf23e86cc4b54a5aa19d589fa24c1c34b8cc6a14172ad0e92f3f008d3ad1cd0f80cc02eed6f66902542ee91feecd53496d675696924a8ae010d90826552a8f0390c36622b60cef270c62557eacd5ceae89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h339612bb88f5ed778c7d3d69e7ac9f1a2b8527e2cfd085b1f8d1d1be820fbc80d0009efc4227950411de70b7080d58d202b9a17f4ab7a0cabd7d99b1c46c80081fa23f419ef108286d1781618691a31f27afa43fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15dd11c65a4047022e34e9bf4cd9b6ce9457ce6922fa693acec9db537ee6b3550380db7ff1bd07edaa215e6f2cab45a39d8d73b0091a5758aff708045ee10fc9dda6a1935f0e923f5512d2a085e0443e54cd9696b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2447fc0717184c9b18b39259509b9904a084fce4d768112f0857bad1e540069921d910fac292dde68bb320d8e5d888d356d6243ab723134bb0dc140a355178a4e8037b128f3bf56bfb583f77190deb68905a35dad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc05319c3619874f24b569bb4c63f9ad83e728717ca87fa86114153c02bbad2b4286736a248b3604f72046d7f9c56b6124e82dcec3894f9305fbe9e6d1721fc9d5f04ae6e1e33f5c1545b6793ce7b5f39d94bf21ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b3c9e26513c8c9821b29eba24d899e01e982295d08df457c9fce205f8b17f399e8c0c205e7339bba3d501e642271598c8e8a54a05d381a62cca3df4a134a9debdc5e01ba16f835b2ac8b4c0c1db9da1dc6469306;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54709197b13a265b228d3a58994b593413d833d1204ba202081eec8c8f2f27f13aab7b1c611cc0e3194b540684cbd4ba47b639b1c1b2d6d51a9f5cae6df8dfe319bfec4bdbee8dffdf688fefa2fdefdde074cc098;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h616e56bac3f8c50daa42296b06fce730ce8cb0569433f3a857b7057d2a40c94c22798153f4be0ca95712449afe03a5fddf70bdee006a9e9f01f945469b1f94db6d4906aa301f7db575b79b99dd454baf26f914eaa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b4966d4b349d3b4882ce1164f1436233033e00a91f5abebc7d32bd5a28babca968e0a6b0826b4ee0cf028547fa993e0e169d7f68afb6016c4164060499d59998ef04c77ea8c1c0920ed623889e2804dcaabd7ec8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4632656decce2e5ecf39a9caf487ad7f1283a2e5725dbd9e377f83ab4f02a36cd9b926554644172e8842108bcf0d15d1a344f3f1fb7045912f49028ab3d883bf8a62922d11644920531cfe01dd56a0de1fea6bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cc3ba8abbdb876105a378f456f5a60c05694caea3fb04a9f99dc863af5eec97c150595901077de62e069d2d773040d470c8b551e5dc725ebd2e0f845ca63c6c4e74e754321aaf08ddc3144e372dea9ecf450ff75;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f5dc7def8ae32625fd430ed785fcf2ae3f6be001be4dc09baaf16b1c43383ac0bb5c16c6d4331dd920d692788f124dd89bfc98311612351001e5aa3dfd04bbfd8557f27c9e896833fc6952465a9c7eb50ff5b498;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdda75930c16988e034bd34c630ff2375fcf63945fe0281ffe6f5243c62330011492ebdb2f8be09614789ef52ebb565d694208a05b6cc7e379cfe1acada18327a61802dc4113d22900c73161615cd4556c3ac3f30;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h554f90b0d606065a909a57778eadab71f8d77699604253fd35a79df35d272a251cd9b7409d89d22c155a3cf3dd374ab3be30e84c9d31b8495456977399bb4cc0cb1a4f7b518198ec09f36dfa3739ba11dfeb8a26b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80fcdd1fac026836571e934a9d0b708207e4a205fdaa186887f1114229df70b145cebadefc07b74031ed972cdbc263a6b40be7c7b2494717649d6bf9303213863e222fc7176ce48f9ff42affd646d5c632956e616;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb887aa009fabc0e780f893ddc9b2ef57a509feb60b2eca950e1ac210cb0280211d9ef119821e413254934e1b50b1234fa98859a895e781fd446c9b0b6cfce1adef1215110c2fb1295b43ea5bb88052da24e47a418;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h224ba3216dcdd3e4dd8c69407b5a4dcc1d6604255180f8771e1a7369514b3729ae6c978f8ea0167be031cd8f4c42d5d236bb708924145d156639c817d5900ce6ad835df03553ff23a2610c322bc0ebfd94b7dde2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46b59b6c22ce91928a776b3409ebea8ab1c29ded79dc796cc1427be1dec42a2499f4c8d8b17adc4f2ee77abe0f033a9f4a8fc62cedbc1069b14d0732ae470de3a00cd545bfa6eb507f524cde91be4ac23868f5c5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78d28be66740687b69580647e0f82d9fb27fe06fdce7b36c55c2bfd9b10bc06f8408652863eb781b503bc2163727e89c1328e3b0c0d9d824d44b3dfda01c3677b416d1482e97c32b556f697d1667888a19dbadb47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1156b73b01c1616dd4398ff462799261eeec553cef01429bf917a9c4431719fd42ac0b4ade4685b35c77b6c0c20bca55c0b34039e5ddebd8e38bd9408fbc30764d7ffa7056f4ca4e782bf5b3fe3acb75c0c1fe969;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39c3fd4228a83c44837c0c98b53363fa628fd1d2c008a7d03688a792719cac06e5811a20b3b4e598c300b0cc14f97c6a24a8cc2712292594e7025ff7892ad23fae9f045b031e301be0df893b6bafe1d5ec17c01f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c5fb87069fee8bb029280317b6535c8823a483861985afb02c66221df74d606bcd00517d7e3e775585daf0c27c333604f78948f8fdb6516b49567a434c6df9c317e85334d65e1cd8ba2fc26895de712408072aed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf665e63960455dd2212ea7841c552e9bd1fabe5faf10da47acd390d72aa49260bd8794c988b1c19c6a8196929ad838ef5100469cdd6b8534d2ac718319f3dced903a66402aa3aa5534baff680cd51cbe690e0edf6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7817d0ca62b3db5f0e1caa7078806f217a50ebc021097da78553f0b59a8a63a55472c80fdf9bf8082f28763e696ec9a2a9a3ec6f6497b530253ffc1e37862d743ae8de223c5edc009f484a741a26137687370e868;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ed5e27b04b53a3f729c00ee5b005a9b91fca49bb49c698ee8c30b0559e4136468a9ca34a662a939eb81364d3a240e3fed430edcf30df2cb225b89ba1efd1d35885f41f58b621c63f650c134582d24971f3ba2cda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfdda3aacfcb0c6e7da832761f89ec4d70a227b4003edddc2d7a360c860f8fd017638d6e16a15ccbdffcef6ba5c93fd51ce34146933111cb56df817f60de10a0635bcd17d8e86adea1346afefaf18fb30ce7245dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h878f10293afc73570ac29b717a45b3a94457bb6106934a29e30a3fe5a58b8c2e6e46dbe1bc3ffce58bd684b3dc46eb95844c66a8569cd9bef49ff65055424a1c4750887bb622a35788eca1a388d67ff69df78d96e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd77278be593eef6972391f32eec315c52b5fbd7289b1dd6571030341ea09cbfa3243b457b158fd784c72d27ef80366f03d31fb2547327401bdea22a66c77cf64281f2eff696c4a9cb8760b67882c40d9aa5b5fe30;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2da8043e0102ec78cd139ab4a54307d6483afd5856e9cb6d65754922428b5dbaa645c58d95c63b3f2f6ffd2d28b3de2a7f74aaf41bbd8e1fd9a98cb4a0ca669bb6182cf51118db6915bb0060fec9d26f34f2f40e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha55f0629fb205a5aff3bfa3554cee28f2551c9b6d040578b488f966185b39b815d3ede4e1f1f4fba61eef302814b486de42221d0484253e738172039bfe7e598ecf5f89672be5d90d5f180580ed6b80145c3fc4fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ebbea0ccdd4ccab11fedbe7847e249282782a471029478e62e3618c0b55f7a06ea97a465439bbfcc5d7f74df5aecd5c5774aa70ec6e62e9c1e4998639fac62cd6d4191fcb5a59ead3f5abb43eb67ac6801ecb03c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fd86fa4d03ee69a67a01ac2f338f470132780690d4ecf5bfd976714375062a56658fa0b4778789b592de7ff950fd89a3aad4123e5b5013aabbe627de14419c618557f9de7e0d39872bcf3014b504f8c12c8612f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82dc84a0c8b902529405e1217e5de16e6579fbaa3fbb54c8a9357378fdd7fca3ef26ef1341e0aa818c3d9f28016a7876e15aa159cafe82f6f9c1578a944a0b6b7827d76ca28acf020031721606292aacbf0756701;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86f6e666f2836b30f6f375902febc90c8f1a981e8300b9ee5962c79225dd3102dc363ce8b24ef561aec1146077084c994bd668d50383b396d9be0e70814eaf16bf9a325616662ba07e3c3565e52eabfa86eba3315;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h644255e22b60a4ff6d930fb7cae46dd4938202ee862a5d6248a2d12cc84997be89a7c99fc5a9e11605233b6d87bb21a9b6399d9774f01b3b424ac68890ad0c8eee3eddb499ab459338c0a3baff63267411d1d221b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7699077dbe048b0810e4b9f0dbdae363bba7d25e76d26e18bef5341bd6ca975d2198427ab4b361fe50b5c4960d1c9223626e904242397ba295bcc018bdc6bb18727b8cf882fbc6aa1eda2af58d48ad0fe493f332;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76aa8a625a3b94601c5b7995c43d9bf7c3b76d953d04860f25bb9943b3faa45c089eef5040aaa59931f9797d209757368c8c0f11dac66d2ee9107c22203be1c48866fcc94eae0f777a575da43a92cfbc0039e383;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h563382571f02f695aaeb472f238769eeebe38738fe2077f27d142d61f4b84177c011264801262522fc7a576b1afbaa45b35d4fee6ccef1cb9b0aa0eef89c157d1f4094085d84af17cf92c577e240424f0d13b27de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bc489dc967772f07d6d80953c27d90e9fa9d1b72dd2f850983826ff2a7a85b67cc8ae9e29923a02a02840a1957f3ea4eaf73344494b07274029277f78b5de778e05429d502bcb9b064a31551bb54f1bc81046fa2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe222f828f29f7d3122f3e522ab0ad3869f4a48d8a779b8342b95070138003ebd3d49b75620badcce47cae460d45f33ed648e25f09255c4f7410514c3e1e4097bf07f4c349c4476d66793ff7f3d0d95341080aa8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99853e91c908b78bebdd29d1f58139fd65beac9c1f224cb2c729bfd80508ac4f93cd2329102377a24c8224bc7d0e2c669a16e992472ea8ba39e27ef80d18c62aed6c9822ea80cfa40b35778d128676770dc9105cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29f8062719d0384547da8ffb1bce94cc3445cdd1a09257c632202c9c52ef59912b0673f7cd5d26906100d0c787c4e1fa1536ccea4f8ac1017ce2db9486502ed9051e6507f38c7eccf289fbe86ecc85b9011e011f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdb31c9dd565a1a932a99fc0517439a99bc12c5798e2c0812b92e77b5eb0e421c2e570437b003085b0ca8f8e3a2fc6d4b226d7cb2aa2aeb4c8555ecb35c0ae8abc9fec251593ec2757d336990a3329c66de1a7921;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf14abdea440cd9b94b4c241a7e2c769b68a5525132c8d8c7b51a1913cabd5525043e8c49c58a6d578e1b1b1c3951b398ef325184a944b8be4b429c10ba29b551848ca1efd5789d1f0e1645800674a078e554a6d78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8d6ccd900eff4b41ed7e21666ec36157874aae510af94e1200b8fa981d4d605a60eab7bb377308acb6a0dc3fe56d6fa82ca2a86ace8bf2a0f13a38b3f3b4ee2b5898e4737822a3050bd9ea414189564491815d4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48e4f4093031444e183d30aca439138686d8ceafbb738044d0074c849daf098b5e7a2d3df90dc2110d065fe336e108b70ecc77921890b36c3528d40a4816e87fbc8c59dad45b5b9ff18e7521e738656cf7c29ad15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cfb4154b7b544859c9708125c2884ccf83093a727c1714ef78e58b12085b0bdaa7123c6fa280eb108281ee4a0e9ddb983da8816c24d4b76ec06ee0899c2f6aa01c4221d194984b7798a2b24e30d193c9bab20a8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c61ce220fd77b7592ac016cb410de5cb64ed7b74692d224dfa311a0ca5967d7e2d12134bddbbd724e3866ef13660e9726457d8c00030f5c3013a7469e81ca0c73021d035cd2559ebd3836688eaca170e59243131;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7c4ebb2d9f157f28c476f3242ab6b4697040bac7ade78e298fe26d7d4350950bb736a92dd199f368f385090cc38ea1d8f36688be146a3fddd11613c6b5f0ab6fe5a6f83380592f6bc9bd92c42b88474d49ac0ba7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h656be246548d55afea0f1303d12fde309603586223038bc8d9798e4118f7c696dd74f062647584ff7bab179b2a26d0681bece72f3aad5a4eda79a48bfba0694192b4ea974bab13876ba052e492370b34762f065fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31eb8470c4a1191e19f7459727e1f3f2d79af824ebf22ae8c7acc99b40f9fc4a0290ab117edcf1bbf5bf17c4154c73d62200d8db347c15f4772f2c660842619d0414e8efd40ef7a80158eb5a5148a6b93a40b5211;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f261b72c456a3da7d666360da0ce2d347c015e6eaf3ef77cf92c35b5aa0271d6cdd775acc9cc553b2ae30c7fb5ce0a71fc04d25aef04c82e78bb91526ee8f149f74d0ff8099e3549dd17e91b1f0aa38727800cb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8deb026ce82fca70f8f2ee1cd9b89b4fac06e8801d9e923da87689952928c29cf8c2066ee51730bb1e51743f2a8362bada172533206427053cd9784b847c24922035b0613c1507303aa5e0d1bb8725c325bac9c94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7f37ee3daa6987fe76ab0be5cea32e2d1db7935c2ebb1a711297b1750ba2787334715f767e21455d8f9972c57e37ba7a42a86a4f3e6adae25da7bc48ad2916dfbd8727b786dc0836c6e149ab0142625ea69a56e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b72eca85a34c2eb789df0204503b24cc4b3e49d1cf40af37a0576e0e6c5ccb304402a94787916a2d5215cc4bba62362546962a8c6ff18a0c6a067a965281adb9b133c6360866c989558d5180789fec4a88e7b4d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f7e5371fea3939cacff53d5fbcb1b06be787d4810449949d0709f97e86f3656983a5ce5613676294c4052a14b0e1d1abe9f0c9deca0ec55cf17085067820a385ccf0f7e4256722d3c05f1ee2846e5d778a5205bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he17b598eb76002d83968ba4e3ef32f3f6df97464acc4d9ee4b8e1b8aa00d322d9fe35f06059a8253d033fc2ffd12b8056c00658737120718234871acb5415d26816d5d6c2caba089c85a338d9c8ad5690eaff61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd93376d6f22105e8443b74c95aabf0192efabf1ca9afaed27f07882986d15ad759a2df61fb5224e7dfac853b1e2ad8e3e33da72dd4c3f7b3278b9f2e404be4d77dba6ed8bd63c244dc5fba7f4a8f070759ecc5258;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11d51a835261614b828447eafca57a5b77bb4bf7eaa1221ab5267ef5acb07db966aed79b9b2b14deefddc8ce967e4bda6acfda0cf545ab6ef725159fcefc30c5d2f8762e35bbc39d3ae1ede037d93ec83c1c5133c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8da3c5a12d7f671fd78ed4a9e6156c70ec0cb7e63fd7bfe08a5ce4b87ddcc074b28b1fe5e9e8ac70fe95bc9d6a45b39cccb69665b90221dc4044c09dfeddab72af8dca5fb95c593c1f77eb859954fddc55dd3ae94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha61e5fb399e03e64cbd7fd4c2f10122e0709770f3ae3f948350b903a283c16977e3e3ac30fafc60aebc130fc7d64940dcd8fcfeda5fc88219e11ea4da82f2ff0fec4d6b1edb994fd2f0ac7ce6046511809876a116;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h262d2c00dc7daaa935aa21e6fa4cf82fa0df9d58669f3334ecd9b69211a5eca0a15bb8245e7988e27f09fc65217d38ea759d6e530918f14f748a3cc8837244878bfcb66be13c1fc79a861ca8cb194f37bb79d41f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c11b0b3e0cce140997a0294ef193f8824a21aaa580d8ae263b07b8bac77874034c0d5fe41696645da8b31a1199df6404dbc55e6311a3ffa35a57afef3433cac9f77474dcdb81fcbeff72bd9fec59dbb1e882c515;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b7d61cd5b83ca78eedc7a7c989c6db9e6795ce4d6e41aa922bd9bf85f2d922080f07105e537111f2a4c05be16ff3c936e230d4fb4184daf1e310eb23ab5c44f2e75616784c4c1de35c1873b5d577ee6df1272e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fde5ab2935bdb12184163fc76a24a31dc8714b2da028f9c9c57db40b3826cda6223756207db9f0e80365190992175f8a9b0a3cfa33cf6172372829ec875dbf043e11c57671f1832b56bf684cf5cea892c7e93926;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8c613cfb2aaf087cfb1fefb897dd01bb2641b5c8cc77655811ce418ee19d6d6ddd7a4456eb6f822991d8e2f171a7ababcb6d1672dcd2db253cd8d9c9f6aa9a178523db7214b9d2845d10878eb24d9b7ac5e79a24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f9698f083aa3d8aa135c6c05e9256093951a70f2e98e1239669d7c2f77da94f842ec99da214733bec3a369110c6f759a62aaee04998bd2fabb4178ab46616de50017e3ced601003c76d7e292363d5851fa3dc864;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h109089dd83e8eadaa96ca4f668f6ffb084c6afbd80bdcfea1f97f18d46d297d4d2d8395e5da1ec28252483539c27874bf8b07ec781955caf55dfe77205ae7888cd044e712db352d3d6e347f299fb6a9e47c9534d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92db472fd267553e96e531a07c0afd510da8b2313c9682b65c09d4d37492221d4bc4784e45d1b227fa57c2fe936ce676ff61830d81723a50d3df6b4f724a9c6c8ecb939b2e3e4f5e57969fc77301836382d6a524d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc499a8d47571c267142fda00a68d7edb4f548e357f91884206806ae86d459f5a3177c6b3e523d95cd4b03bfb9c355b8c287eba44be9234a9dde6996e9d279feb00fc64d0fbbd9f1076c068bbd24af0902fbf39a59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a34982d0faf47792b195b2046f3b8526f93ea5cc7c6dca02ce622830b7dbee9818b6efb87f3a64b9cca2083950be3fea955869ba261aec3cb23a85be73f381e194926e9b90f9deb7c460f215ef8f21ca6e47903;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94e8221128c7f226250747083eff781995bc5ebc4dfcc29b44e7032be78d841c95ad633217a894d7b4d57b626ecc0942a577ddbd79981333938cda430c58b6595c7f78f8d19135e06cddea3ce0b1ffb23c7c85056;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee21b6d4f77196ce0db5a294553bce33fa606f53e8b9e211a1939f93bb19561b84453f00ec28753ea634b6eca9342542dee523dba71813dbdd360f30ec06748f5a37a0d7b93dac13f882df776d4d0fca702709d23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23ab9e2aa6e7f0ac55fe53e1b784ba258846b3b48b7872a875a117ebcbd7af89e33205fcb40e6cd971ebcd306fa2a5c83b22fe84510bfa77275e5ddf06360507d8d65281c32ce85638bdd9e1c753ea985e45c5908;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1fa19456862c3dd73f1eb0cdd234934609c28f47f3355127adb83106588c55ba064c55e0433819aee87d93dbd138b7464e95dc522772a9fba0adf4f4a87bf0961568bd41fa320ba4d601efb14919236811519873;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc266212df22c80e291deb1b98cf705d76db14720779016d7cb33b329a437df0122c27fb2719701a6083fabad703aa46c74d494a4caa47e546276dd6c0ae664acb11968b9bb2d858d1714e712f9ba3b5c68d0013f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h863f12b22923641626a5dcb5c49623bae390a3aa7d216053ea38dc04ceafa496fbf4e92c1fa3980a8d2418a40db8ffb1a2d94a886c2f42e36dfd1b39983c5f4b427366710286da0e579b4e60d8fdc013234098033;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71626e1d37eff761f7b095e1c32885461e3159d1f838ea0abee91db5b9cde08ed3f71e841fe8c6b010517c70279b01347fa0c32c6899523d80dfb2e9779e176de4fc507677015925b67a4dd51f742d7005ef233d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfff372b34a61940ddc5f36dd4315f68ed61c5ade93036c19605dd32882c1c403df68da5bdb6cbe3ef8c40686106b8e697857b519a29120a196f7c8ca9cef2a3a2e3cca93340803d1b39090203fe715dee1e28f93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7088aba58a830fc5c5dacfff07ec24e8d2766ddf9b686fb161b8157c246e92d8c7a12530579611019eef4614031e22e115ffff901b2439e38ba6ecdb0ff97ae1c7f3928128d4d75a41e7c1a170988333ced0b8a3b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3404a7f7e8524f52b6c0cfbf0ebdfbb721a45013ce31dfe585ed4aabc2ccfe458893a7b286264f924a0000858e2fea2f16522b4e5f1145a0a2d847a9921ce928b014697eee4e4a620c5dc4d71b2788b1e9104b00e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bc07e7e371765be64081bd0319512114d6bc1f338fe2217626747e90c07595081cc1d2616c87184817e3bf35f2f39a9b475eb9e1bed7c39d37dd4533d73ec95afdc7f915f77cd9011dc73e3eb4ce4670f6a24660;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h669329dc3e1d9cfabdd157c35cdb7edbad32d287cdbef87096004906ab142609815467c4e7dc0cb769262ed5369bd2ab31c913a13eb6d514c1ad1ff6a18cc1d2a316c6354dda805870171c227f80ed23532fea231;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f3a4b66a790a878bed328cfa5bf30e1239750e5e0fb8d3919131fe8c8c51d2d958580ca3f1be7714ed3eadd35cc4bc2fa628bc9c2735fa8ba17558dcc97eb2951fff47a5cd770cd5e6d044f8dec016e243779959;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0cb22efb7ee3f3852f76881cfabc0945f4dab424872a62a4eb5f67250bad928e04b5bd540a0078826f4b96aeabe36c6bed9c5d245c0fe186910b996ff21b473d180cca2208ec27bda4059fefc88c0e6fa86754f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h232c6c801106382bb66c7c05c72d50b2d6bea1b99c13cae6497960b93c46a605b0770210c089c511e1eff21ef71b4829af975595f712a7a87ee8d9faaba4b2525973e0b43af3628596f5efd9983f15fd9933639aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a1a5e1e5be7817bccd78c6cfa4ae633682754aa4ff554da63ef1ac5dbe71480faac1e07786cd38d7e00650f503783e6feb46bd58767b8ace6460906df91db7e1bd96641138f204c16c692f22c9f9ff89ffa8a2ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd914d9e8ae9943a0854337a7429edb717ee2bd4ebedb0bc87a1a551d292cf95ffb4754f6e642f92f7e3e23a14a095a4230b5b0233cb7043a3874212c9d8f7a3f5c4f9144fe247936b5b924dc0b0069d7a5c7f8d3e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd977f72f74001f51716e703a1df249c16b5bfd9beb1d017ed7d1805768ea4ef3a7a47289a715a52f252cec3ff47dd15392cde58adcc958864126a7931b312581208f629f30b99d07cade5e13c9999d728de872fa9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6842bb54b123208c0c3b7f26f858cc7541778af44d3a2ce8cea75b00800eb5e5db75eb510f5aad0b419ee6b675af6aaa95505e504a03b93106ff17a1f51c2b1b452b5ea14ea0a48caa178382c0ade87a9ebe55138;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc69d95ad4a575f7b10bf7d3386931cc5052898c6696f951773fb58501b44e5f83863c4c3ad10dd1ad3c112853f35d29d20bcb4744e0c8cfc430ef0cb75b6e6f84b84454fa1c8558806a91a6136f4f3ac11481a58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c1ccb7c28821393d26296707d090928f24c4fe9c336bf0dc1861b3d901271b3984fd869d23ddcf3e452d8eb6517da906210d59c662cba6c461fcfb76f89b3a3af6a4d10608a8ec69b827b160e90d341f5ba38c39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16b7fcb68f4fb943e007ccee385fb4e209dfa779a5c53a7ffc29c6a694637564ca411e8381b01e27ff5083059a12087651f415e067cc75c4c9b77d2cb1abe745f46d2fbc221fff872cbbb0e05afdfd93225dd0f92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h146ae331e6b7128a2dc6e9136c4d6096d3142e0dc2bd4118fb4e766b712d3b60d6e749a2a94a8e28f61ea6650bd505e706708074cc53fc46b85b0ee0099749de8b72b1bf24738c2659e43efbfbf0e63078a2ef331;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bad8e34a95720e52ae9fa45071a3414a959fb007d7aada19b08a66685a266e3f108d355b248bcc3c4b46036b71e3b787ad57e364c64b2be6b845b242562d8b96b4aa8be65e90297263db7a879a05d8245784958b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce7e58d3cbdf60727619f5e33b6529c421d17924bd5d388fb01ee86ba2bbaf5ebab0eb7ef8cda852996532dc30f3bb9611fd658993d61aba20ba1b642fe1f3e32da1645e11ea060ee1d68a4b37fec0238cf34af32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd4a04a1f9d2aefdc094f4fdea7ecef21c5d3dd1fc43ae937fc9c703ef7ab0341f9e78da41305dceeb8eab51a6dd3d21e2f7a241e4806f5aec94adafb9de5ce4b7dc650ca702345f29484dc07bc511e8d89fa5929;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc91bc8a2e3a073da83708b5b5c1bba510b1deacfe5d9e9a7f31f40555fea49db8f9073a3379548e752d19946daf4c5deee844384eb82b6f0ac48bf256b1c64914ef51f876ae49ba507aedddd369d2293f2af2cd00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d9e4304f021b01e1fc3380aa47c12a42bb6e1e66d1758fd96b1591a42071a2fe120fa9e7e1e441e79d09fa8e0376cfd48af466afa63ae4ce2ca5d7da4987a6b6a63815e718ca64f63167823dfec1d3359198472b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e1e8da6632939f44147543316fbd622ba8b6eab1fce29ab26fa0a138caf8963df7f8ecdd98c1c6b0bfddf212b8d4c18c18e5ae6ee471af0b49c0e62a2b02f05d4d9025e6ab67d93bef0c65d9503af971323fd6d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he99ffd9b27c7238bab4e156125913879ed53680c09ca4f52604a59363f9ed89582d11333b20779f6f0f26031d67ebef84743ef1f2dc710e09ae914e0d6179e2af1954da526b78bc92e034fe99f3789ca03cdc52f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18004416ff0ff527328fa1cf995ca2be0bfb4bf9db3fcd0b981976517813856fa6d66149164ad5d292eb29edb88f578f89893a1d800fe57c2aba44025ef1df302134031dc6bc109c8aea7365385f44d09c0ebed8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h971de28dca09cb9b6db32208ac228bab48093dd4511b97f8c9a5b8c815814c9ede5f53b76b5d38b6833706c9d3729827137c9d58bd8d4568851747ff8c60f0d05e8a0735d698baa114f0cb529df37f6881800a6e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9e7287ee58de7c4509a084051edb9da4d9cba66eed5a7a8380fb74925316f15bd6ca482143068c9d3851ba17daa5df47d7249fd1fcf7e906705ed97ce319153c50b9917e1a03d92f46864ee92f8ee77cb2beb7c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3679fa24b60dc47c25d814a1ba2f0d02ff80bb452faa8d6abf34522ef6b139ec453e27fc0366671688614111ed85b72a704f6cecc9d1bf1a4168fbe29c951fe8959c565d37c52892d8bd147e785a3955e8a46020;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8f3e96fbbed548201a035e9ea87994cd528572393398b84d65823403c7943142810f5687cd24b311a8cbca2367fff7afc5dca7e021d11ec65614f0555837c8c7f1cfa0186ae2db8f881b53088ca9a01669a22c7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h809ac98dcb2e01abbd252d890c95f0bbdfab905a5185fe6311dbeb84297fe679e6a25685badaeed6faa57ea4c5490d844d713783ec8fabe1feedb9a5afdc536ba8696cfe4dc4b067f65b56185386e49cee66327b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'head4e4325a1d5f562fb3d0c0244d3e0e1ab3c71d4baebdff0db128fc40dbb4e3e27b70cb28bd2774ad4c844293f84cee6d26006cd82a97bea2bb367f3376a6551b1af7f98a5c6c160425e4f13a82a233b3eeb471d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8ebd7c1085c84636d3d45194bb87ea6e95d7dd014216282b100b246118d96c8b6a7c471375ebdd1fe0088be0acee9271cdc4f4052ed468b47ea53710ca604d9d3dca619381a080852a36297417d61e8233de6fb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha47b48cd903145b29a9324987d8a753f8af3218423d596586120e5e29a94b3de3e483bdbfe7bd1b87bf7c4fd107a2475812accc2bc5ad0ca064539fa4297cbad86c1a2769bbde86b4851a3f61176aa2c852836f08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8945cae3eb321dcbb45400cd170a80ab67e8ce444ffe286ca3ce646285f9b1ddf325e8adc4f54785fe24e85c8f91d4ea5c63e9865eb95764b900099721ee762d6286aed0f1b48bdf3b60b5d500dc534401fad81eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bfb13f961b92b2d957a2e4cdf0d3e11820b188bda96d2a100eab4fde603487ccde16edc3cb3a022b25f2ace3401a95555e2acd08a323fbaa062ee367b34899bc6116a81e1a4f7760a10062f9372c40980c5e64ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7545855b0e0d5ec27c1320abfed1b48d0e1abc0bd439c93e120f9e4cb5faaa1b4f38449eb2cea71dc66440a12e6db97c67b247a110bdac5bb4eb02028a8463c4e1ab225351904e33ff5e222dd13ccf13646990b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1e79c3eb888469878503e20c102bb5e6c6c596f8fa104e9cacf52338318268588a1dc1c107e9672fd43671a92dc86207d792d13c087568b6da4fa2b28debdd825e86145c21681264ac7222717996761655bf1f84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ac6f2196f964229854180e6342a9fc1f293b0c623d14030940b4624416c9cd7c016387901b984c36702c7aa4401a5ed6ce494db9bbd19ee3261a11adffeeb47aaf30db565c25374cf8f3d309d4ecf70ce806985e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d8a318957958a8314c6522bda9ee823c3124c98dd8fa04ac640a5bf04be7178c0523b1163ad95ffad8a8ea858cc44767ce13f476cf91767552c2f1f9ddf79be9c96dd816223d815747a98f35b006cb7612499249;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61040b133466543cb4b12c78589ca7bb48ac22f44a922df4d5906be108a1f0371d3ef82af91a6857596ae85ebfd3de37f9320a3a78916e4544d4f7b0023af7fa71ceb94489d446f0b1254ec5e32235c2017225345;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed61a69547f80670b2e3499e9e2c97f1fda5b0fe71161b56de57649c812d7e23f30429915692024dc663c78a909a5baad35c16b196373291359082189cdbee65879f210f50854b4e52671c9273a2c78ecc6879371;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35be61b5c45b17515b5198f9925b7833eea1d2a7bf0ac3e19f360c2a6258a7da5dc30ea3a9b3dc9c5f84be1af4f98624d1b3987357fd01cc5155ced564de26a35a0763a0631a132a705572af9f447e9b834e062d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf30fa9caf2d92fdf1c915baac1fd476adb920c2fb4ee748c11a7546be26625a32f178c2f82cf448fe5b367d2a761fbec1fd9980917f61de412bb0812e192a7aa7855980a0b0b2361c6b40b88d18b4ae8fd5139c5f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd06d2f7acb166d8868c3cf2b4f90eab239278bb0e41d7845b52fee1237e6a472eee1d9d106c1c6de709daf2393baf77a7776316ca36e70a16c97d30c128307e891959723294f59a271d7eca868845b8801dd15441;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9f4d6904b05b1aa429f37ca9aef8ee234c0acb842e1f3d70480bf11fc16ecea96bcbd93e1509808f1ea7a148a918656e871640655c535f4714edac58061678d76edd15dd1bde8619b5fd234b72eaebdc545fd734;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b67873f3299eaa75bd2f82604663bc49eedddf99c98f16d3dfc7f35f420fa9f75ba06ba75bc4ab4a507de8ae62b24f7ac6f129a6e49345ec5a4735c24b4db53cd56c1170769911aad6e93388b1f6b9a668cc4cb8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1babc06caec56d26af918cb764e6f67930e7c3c8708141ea85b827728ffd68407407eb8b6856991940cd046356f800a2cd352e8e211b1b963607f5895a8dfe5a2b1ad1e50836423e12cdb2ef790efc3aaa490bdef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9703e4abb7db9ad51f247e02631c25ac9d994ba84cec593861aa014c361ee90388f9c38cccd1c8842e8e3852cd626868cda72dd64c011c437f74caf33a928df9b3fee5ea296686dd816c1a6e94f93c03d7e9f6d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haacfc6a4410fc3d169f2aed3df046b3380bf57baa32c5f706124ade67590572db7a4aeeb571879a600130abd4ae1eaf09157a6fbc94f059f383bbfbbb47582b259bdbf564fff3d7d338a567fda241d9564c5c24f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68652aa816dfa232f4a583e5d17e83b2322e3cbff42964a1330f2471dace0bf4b266e9c222b0558e424f628f80d22956cc2774744d3cb4d776550047e36f434e2b7ba462cf72940975e15822ba12c0acdab20c94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h850adb1d4e5f1b06e19447a4541d34d14499ebc79199a5e059ad209b8aa8f1f5af7b08369071eecff0c370484866243a076b2a4eeb00367b5abc00c768494c37881e6caeac2dfe7c729213aa76bbb73ecc9573259;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17e5a2b047401c319b3a6ae67c2827c3ab3ed327d3f0ac77295b1f22fa454c1928cb05b8a9928f87fc6b7146bb898b114c83d52ee4764ffbf7d1ed460f653d3515427f78364ac1e210dd65f6535a9bda36d1885ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1945afb609571bb46cafa30101d3795696782572ae4fd39e67ce70c091b8f0851ba4e217507bd69a6d8e9a255e9aaa76bf1cfd8a901de4ec36a8606bc7b68f554d50a5d976fadbe613392782f11ae6dfacded32ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8f466f22df5de9f96ce3de679b20a4ff8064109edd724ec310f791ee6adab33a27413cdbf4eab164b93e7f241d848ea57d5daa51a738c91ff11aae64bacb235cccd75af66759634316d5444b5880b12145597c04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55c584d900c3d530b18d1f35656156006a56a316747a0e82f8bb8e3b4392c374eabb4062b483d9d233b00e670ea90fbcf0a44fbae45f66e64a191baae8e5031fe257d354847ae538825e9619e4c82cf0cef135da7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h316eff49632bc6fe54a29fbcf042cc339ff16d522a39eb528176cb10e5b51f82812ed4779657032bb29e0979f7b72c7bf02cc0dd5779ba319882fc7d629ed947ab6d558cfa0125255315df7c118afdc98d6d1f20f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a831fab9087d61dabb56e56e8a404776a8af8248904babcdead446d225e097ffd71d31a45c29b5f061582ff195a61ddc978fc0376538ada5457bf8d41ec4ed19cb2cd92ad24fb955b948c398c2925811bb134b6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cbe8475cdf1629d1ed09d8515cbd85d03ea4937107aed87dff54e151557f8a042fd6f2a11481ec0752d12e9fc8bec80184b9e4cd490b5d73cc28530281afac53ecce5517a9bcfd9413a777d71d7fac94d3dfc56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3864a4b257ea047df9fc46cecc73044ab67c08deafdd9b93903930b48e3ac51a4fe3477af2539823b9d66324a331af6e509e6080d721b23894432457e9d492e6e29ef2dd8fe9940245c1020fb7c42a114c604a9e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33fb322617cf7f599754909d0521563b6098e5a114b226fb1f90a6b1cb87a7316028969c479a5b97abf2f2d89ba547e75b1c88033d79ebe4e8b66616f57cc098e12687ba3be6f3dadf703d77d49fc6c87bfd437f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a2cd5f682466e1a28757d3e2d978f7352e41050a363498b58c82d0c994fd90205f18ecceb652bbd7550e53f593cca7b11feb0a7677715e1743fdcd0b700f38986a3a270f7c08c92b7c864f0ff777cbf35c877015;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde6fe1b29fbab527e8b94b215f840e6a067c901b2e3155dcc446165a06a0fa6deed0b12444755ea5e98f28f1aecb018da3e167dc6108c272bb70fc010422353c4b700acb8809d289e1dbb2a40189cb536b07cc21b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd12844c5cd3c522a3ab0e6ef2ea58b3de61b0a36b43b2cd7a35236df50b19a4f5e9a04efe31d3d0dc1e47dced824069e05712cc09d3ec633b0a2b1359016c13c1aadd0756ecfd5aec1c18d08eae662a9967ee1a48;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h802c874aa18ca9a5e8e18aea6bef81b4633f772303ada4e248d4670fbc2ed691259ed0d0ad995e8f0bad66e7f97356577afa0932cabf49c59a1f8348206ad0dce8867f3f15e65b6a25cb83cb1505dda1c8375ddb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52c19755488618eeb8b2b759dbd645729cd00373f44c6db5bb00024528f2c9dd84b1e20429a16f089855d2ecd18aaad04bbc2f98f960272b94c7d17c49263cc79164fa4f8e8db68f549051f31a6ea4e226f29e202;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97d8855b7058f483d7fd0148efaf6228a797f38ff3a72775d2a5cef0e0532c04d0620e7cc6cc58cc3c89bf4b1662065d55fffa3185fe49d8eccd541c1270bac0e92aed50e06f1ee4fde47669fdfb5ce381928ca49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80c29ba0e5fbeb218a008b89927f4c5b228848269aa37ac73467151aaaaa99cd73f37265e6d7405c8697272e744668b93d87003ccc34d4934a3560f61dba5859b2b12ebe4a490adfb7411a71252fb4682987a138c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9909f16559dbb646ccf076d3d631d7d87bccb3672fd1d78e2e76abff8754dc2d270954a26cb195a34edd6d73895a2b5fa465dab036f36682a9d49030faf8f8db3a6da1878f62a143b08c6d95116c18683dd102899;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h898c60c6b11f632f95adb3f68d8f3086df3f9bdab7e22fb6b54b8b2e37b33cb376f82e0a05ba425f7309c11b7d7932385a39aef6de630bad0c97c64c190c5b5331552acd3a6658da449b96de5a35abaeade30e531;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc12951162e07eeb06dc39d51ba39eaf0d267cc70dceb2dfd3f149190c689d78930f70d80f1ea97e32daaff242d4d70533f69db1c543c2b6aec80407047bad02da7caa6b0d322bca5a41edd28544e6755a371b56b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8615b4bb25b4bc8aa425ea53b0064af8d67d0f634e8213f6d4f8dd4eff805502ffa4ab66132596976cdf2da7062a6156a067a71c6328d88e4d585945e248ed2c8c8d62bd23f343a42fbf3875fbae50a631378a42d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h999fe886adca0a5098a343b29f01140aa2837e8490bbb1076dbf24dc0b4ede5ff4e8268724bb6598972317d25d400b1e3d656577099bc212bd956f568148d654b1bc954c48e74d31a0b1930a42ce2a219a5cc8b8f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h356bc917e78f3bc8654d441047e204bd0670e681667ae76040fc7fd3fdcdfda6665d70a2e0352102e158f9db419c91d658211cfe67e140f43ee65716c09d57a5617f0cc43b423c47e2a3137bc0dd4d895c8c7e61c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h164bc1ee69bb7a690cca6da8aa66005778ad5d9e0cea33c4a871649c02f27d7f1ebb74238b22ea28e0f13ca91789eeceb9975e4622a3e1bf571ac3f4a5a9e3ba39a35324cc3998e685cc0989cb69a28d001b878be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf87a56edbb87d19f95d8c27a8a8f559e8e339c6ecfcd1aa0372cb1113b528e7706142b33a5832364fe46b34e423521599f86efc7bc3a584be9e4666d61f2bba14a28e7ef7f28898156f758a8c1cf6ac9d2b742e0e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h308a0fca430bc9014f1f11e262c87d1740e7088f040706243f26877008dfccef5b4de000a421bd0b5456ef5d13aff7a08b87df7f13c016fab123b65dc73973e5db31a948092031f77aee3976e34a429660060fbb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b53a619150b81cd6732906354f6a4650d2fe9435586306aa4360170ef639eb11038ab3a3be535bf1ef709ed5f3883caa6035e9165335ac7ee1db503ba3a43c5d2f1e682ec1cff22c9238427d785c9707ba97a972;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c4133aaae3bb6ff25a01317feaaaec54cd495a120e766e27d32372b864349113835c3b2db0e079b7afa65f560f2eeb598eb66a652ff953c32527898540dcb82a08eb59f1f5a6b5c74add2b6e1f0ebacf2eb4b0cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd17055127c4c1fe02b69ec03ac34e037c942ef560e221689b9cdb1f8ffba611d2b605057692b0fe3643746029432dbf1fd23d8f74c2d73f40532ab4ba1744175cda1dbe1993552bb48afda4668bf2dc54e0ec4e6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecc7a3401adc5b7c9e65a0c5546b91884e750f9abe3bf9e1c0bbe4dd9b0f76fd6491463dc0eac2d5a18d18cd3c5a9cc73713a589eee4c8224268f49526a400eda81268afa1aee3d7b17c5a4d8f94e4f24c9bf3ef9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1c9dcb470659ff12d1ebd2562beb3bd4f0b72bffdf982b9c12ddddef312decb9e56e36d918da355b04142909a532761fed53ae12c8d8accbd120c57fa5fbe22a1c291673c762ad09148f0296ad72b9bb3d723a45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55b6d4e294f693364dfdc52440af627828cfd0fa533d2bd0aab7af2f7938c13ecc6e11d4aea76b3eefed20d77a9cc0ac93bf982136d148c6eaa2621e020a834e7a1b71ddc47e77fa0f9ebf9e9244ba1003ff7c0ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c645b8ed32f1a1ca5feafe05f5c2e6d1aa10b33f45be0de893701faf2b36837bfb2be883baed61bedbb20c8752c20348b8bb411c4492edff56885e730319973ac62b34be7b8f051f58eaad8c6f112dce6fdd40ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c2bc380f134bfdbec6a93e702596fff342c2a35fd054153d17d422a9023babfa7b3efb97079e68cc089321c8fe27b30f2e50df1e2103421efa17659a3055bba3fe04e9e7a2ead8f1ab543ed048effdf1e5665804;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0d74daac31f13e3785b0f540536e9152b76cf77cd405d6180906f415f1fcbb345193c2986c135bf27de973635f8790b885aa551b44ffa884bb619dd22f1a948d61e75b4e55ae7445f350c6f31557ff0d26330862;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bba7794796775cf3366f7703cd9ef51217c61bdd2f49e9e06695f4e6bc4e692376ee4b09c77a08ad0cc641768006e8dd411471529e1adb63d8c7a3eeb1d15e2bc5a779d381f44bc8483c875ac1a2389045679ea8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e9dcee6eef699054e049afb6076242d51f8d652f6fed7432765ddd8d6f83593c8672aa20400a5110a0a9ee37013941639628f8955a076bb5b74e5157fe1e75885a7f98003c8916d4380e6be79747d6cb21ed381;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he97765792bcea9f2da5210f1f8bc5d9b6f82eb992c2b20e4723937e2b728008f50365ccb18b2f0888cf197fc4f35a886ff1612ad0bbc8441680030b0b87fde7a4ebff1746cf957c53132886dcff650da8d7870ce1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2abdcc42dccbc8b714ca09ba7ce127d298cbc68f1bea7860fb433a5d8e1771fb7a2d84d88acb3aec89a6a8da9286262d34b0f6ed399d54e51125a62da65b830dec358146bcb7e6ba0bbe004efd78230c3c8808e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9f68f9cd31142761b4b056d475252bc017ee2f01705e095d9a7636ec3d8dfc88b52efb2ff984124aaefe4c31d8638a7fab6edc68cb17aadedefb108d991a1ec92d9b35176e08d2f97ad4d65f391fa2e7057883b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14c4e2cbf9ac2952e7396c7a1ce835210bfe08204ad84749b4835f861eaecd7bc55a3a0b057c7066cae3ddf2a37fd4f29264dbefc9be852e487a775b70ac259b428badb75b0b7caafb0cdd512d910d80808f7dc64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bb65abe52981f2454e04336270b10cae7e13b58a1cfe2616cb6a76aaa10659b72a3110c6e75ee98785855fa6a40d82f42136f61b078b4f0da189c3628467c6b80ebed397bf16f34c48beae456315e0ba98106246;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heddf88bbc763b71e0d29bacb7360473dca422c3790abf60d75f7ed0e63f7cca2d5dbb698af42d7eb6b32049b540b3081b0e01626dcb680bc6d9e32dffb5fc24970b5f1964a34c02af837a3ec12edd092d8e3ccd52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf963db41ad8eaf2304d14ac40c2bb2ca3ed7f47d88a8a53cb42cd439e1897a7d6c4a01ca40e8696780474c037b3aaa05a5ff9b9da15d8341e3359082efb8baa4b8a80aacb3e456c301d90b666db89c1be6c7f812d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ee34c5efa4e82ef2f7cf634ac59e6ff2c0e3e60f4a4da3162c0f26fb9d494b828484303142d1df55a15ed041faefed9f455b4ecdc893190e61429d20491be340358434c94ce6ee76fadf1e1ec150b698feeaca1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h414724acaddb46ef0adc8eefce733ab443d23c196cf901416dbe45318ea1b58c491141ebfda3abb423f3e97ebbdf49ee4a6cf8ec28e1ce0747a1011f4af69d1b45faeb9c535609d59c93c991502bb4cf84494c6c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5004b685480eb88789caa978cf41b838ecb5ac24853e9a4c66fe00729cdeb1868bb2579c2d329c547112982ebf1544ea583f25d79fb3d04413e4a42b639ba721d893188cfc313e771e7733a8d43c23f31a08b09d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd9109f8312ae52959bad19d6251dbae8bc358bedcc8d4d23139d7c52cf8a5125dedea8af66ad322e264c696ace5e1c11c129b4d1679e5a5d93ea34b296b7dcdf1afad70f3c9e3c660fa202ead1bdb99af48b7a25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f9dbb6deda0a15230f64858b2d77ef82357ff61386e5a1cd89d8acfa4bb4b2f4f985c97f8b186537be35bcd2a2ad7cbba3414409cc05a09c397ebd6aa8a7ab7cfd1b52b37f86bd8df549814afda21d344b0afdb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12af94c18366bca3fa2a601f2331adc5b9d841ec1a27a7efa103666794f9e565c13856037c35406875dcd860f5cbfdf49317d9d0676392a583e609795cc303b2770f5530cd036a23709c03bedf0a695fa86218a2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd856c107809a735d57cd48c812c39cea7952f11ac053b14103c5241d8ed8e765c7e6c58c693ff6fe41873b3b63c6404f26c72cffceed48bfbdc69c3544b80d5b815ee3f34b04b6d34c072c1ece7b522d5ff04c1f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h651f0eb36ce263ff55c7c9cf8908a18c1d05291baa4ef546cd1d2da00018266ac869be150c7ec45b71533010ac520bade4e50dd9b615496ce19b2189c5f50c5e60ffea181a8e587ede407ec16fadc3dfee2f804e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd79436c8a7d01da6c0219ba6c58fb3309b7d7c5999f90d21aa5a7fd7192c4cb9f1d2b39f6c763b5a6c86c15252cc5cf74098ad897c03f4067f10d4de599f564dc11d331d9c260d3ef7935d9f796d938150fe7acc1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30eef6570618fcac99e6438224ef013bc9aaea7414b8404636367625ca7c797305bed0a4edaaf626bc0056b80345caadd2edfbd9b056fac807dcce2d93d77c3d775ca17d53c69d7aa4c6308a674bd11aa8df2515;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8621e0b9b1ad8554d4646175db60c3b1bfeade5f7872c8dd0d65e0ecd6918dc57220b716176875c540be0dc1ea8a7d78ab6ca0621f552feccb02f714dc4421560e29a852776a49cd138ff4bf37408e24540b43ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99055b40f121f6a9f3f2e67cc6a129794ff838151841df5db1927789b569af16497ff8fbf701a665620664c9b41edf6e08fed5c299effa0a3e474e401c93952efc463e49172f0dfb82d05ece387c9d6e058cd74f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5ce0404446ede451c7a8981b086dc4bedcfe2f994fd2d665c191d9f07db20168756ed671eb9c1fec26f32117069d4c1923159a6e484d3b0e0c1ee3d1a336e0538be88c88deebfb16103561d93e46d443c0dd4471;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cdd0e65017013bad3e178017778b8e93625e041c802febc3bf0808684daa1450f2c2b92bddfbb37672b656c134dc9b39aa42faaac92833be5b8378cf98775981caf7ca3557cdf57ffdf7c7d4a135ab5a10e4488a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaf1d433cc99cefe1cbd55609beb39672cba6be2a3932af8c59840480b2ec4fdb6774bb684b59bbaa2875e5c049a5edca19305ff0fa149ddc2e4e94b7cf98ee730e46228e529df813fac7453b67acbf40b995b662;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54060a59488443c11fbf617bf4e18515a81d742ff45a26951f244842ce3cf89c43575f103a0deaaed96b594b67873de9babe981096e78a7cfac3ea2daec4626818705f81537975b204fd431a315cf04410c4f4272;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e8b61c7f22ef845c138a998c936431eb07974c36e4c07c759250db8209bf6b8886af68d05a56e0fccbcb2c43cc00a1fb4da1051604a24ec51e617dabd09bb973ec05986712ff9202aa4265d1bbb8da34b514de6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd582bdeacebbaed1359760c8c547dc5e324b0654a81637cef87d8288996269034b6dead8b3015b327bfceb5c9c6db9724f15382900c2d2363d1891cec2b492936523b131ad7985b2a17a2ceb157e5d86b0224d6c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h299bb2a4e585bcf60d46b46fc3a368554aa091a1989a5d7ec235739b748f006ad774bb97409815a06b16b2380f30c23ab9e790f301c876be1f9b9eff9ce2e430c849edbebd4041e09151c6972983667494a61d907;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had0b5e651e0e1b78f5af269aaedee709b5a72c52f084889dd8fcf7ba4ce6ac8bce6e50d0d143f730ab6551c8fcdfb7111e253e7013560f2061d54847af104b4e3a4dc2b2419bdf1bb14052acdc23424965ae97bc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf71323e7b118f1cb28264cc683cc81375519a0b4bc930f2048ef1fd324e623e5821d96ee8aa10fb91e9a8f151da4fb6a9beb5d9c1eb3633f0847015941f3bbc36f563ca480d458ae01c4ea189bc78614b6dabac5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55fe294c12a166b03188da224f0b83135f13901e2517e22d199c21977aebcd1b6e68af1352fa08ee977d2c337164927bf0f3928ca712756b613c4aa819f3aa86c942e07c301cadb83e6baba2640a967870c3602dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ee343016252434429eee8fdd02cc27a11257c6739a4ab2e0602d718e4f25d8f3fecf276154bf49bd7558685dbb014381da501de0b1c6c3997c0a14ac7b6a0b3e365db2a411376268120e589bf4d10bfe3b31f16e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b2b83866583ccb34acd452dff224340a8703f394490f8a894a9d2a19e2aca31fdd2b0b22105c8f250c08689d2a33ae191416296adea0ab262eb2d36e6b386ac7b3828c6fc89d9ca478b4d6d054e6fec76b60b3ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2c598dfbc3e493b35dc170b7327dc48c2c3cac4d528078db53272abf9801381553216a580fe5299b0812513445a82c1b2e55d1ef7b39ff668a763846afb9bc268745d1ca13bafe27b6b9183a88247a281dcab61c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95507a6acbed15fe8275007c72ff427c8c6023e1edc94626af5a444b021d88cb92c5aa23a0048fa8b85da92b1586cec49c1a86fbbd162076c33b29b22c3bd614dda2e08e21a43530dd8b3ad3c8d93018539b0510c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb38b602235a87b0b2a0d5c41bc51fdc0e99f17f01ee8c4546e9bcdf49be8fbcc06cad6659efe2b9b32eb5f558c2aba9a8866e6008f42dfa225be2ed69445a429e61121288b0c740dcd993398cc5d493ca0e04241e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c33f4eaee50aca3fc80c1b7c2ce117372d7652d628eaa8772f5b5b1fa80de54e93688ebf19d020ad014ddc54983eabf5f36d1341d0961377db25d2403185f2ac2a936461e94a112b5b36b2b9b6b793e903e8c3dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h761ed1fca74f4e8acb1b92421ec278b50c13082fe7df5d83ae7683437ad9a4749a850da24163395b87b7c3132ce4c031500105ba760cc5dd1ac500c22e1150818f70c0fc897d7c9b2967ac3abce5c60b426158dab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbff27ffddcd601b6b2ccbba66595c37a1dcdbaa78b4a49e75647d27aaf3666bc72ca49f018e6c8bdc7e37e56666db4eda4743cea9e01255aa6c9125c8aef3e155673ac9428be9d281639c2d44966ed9f5e6d8552;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a8267fdd5f69f5a02b097efa3aacfcc118db3cf1f0dd954440ad678a3ff4010ee8027a31270752648a660bf9ace3f792c23c4c36abbef7699ad6384bced9cb864bb83ee6a07bbe3bb1dd49877c8bb60f04e36bfa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15a3f3df38c7321c3af941e3d1d6a237495458699d1fd95e2bf312e5fd8bd5b822c670462b7dc2e980d32f7154b08979e5d0fdbcd07a0cfae9db3813df33b65ba7c24d343301250af609085dd6feede4799826a62;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h973fb98d656b07237d3ae12bc9b3bb609c602be7652651f15446821d80038657b4bcf0a5348b6ce54c093ef23f3bd4426f0eb363ec15b7b8278697bba586bddc101c87ba41e868791ccc1b4c5cb0b00c49952bf03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffa27c574e366db66ae4ded5698ae97311bc1c03d83bc5f73486dcb4e8cb9f6e57f80ca51c6714189d64ba6d0b43c1ae4b638e81eb70323c1babce9a6052bcca9dd1154bdce470e9860f6298bc66761044c76532;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3ebd21863a821dec1d4755ed9e82ab86e77f327f4fec40b552b5a6ecc64d738c98d213098fb85e61e0e8acd7be07e60699a85271403473f4b5b638f54caa201e6d22af25197f86acf1f1498d3b75d7dbe9865288;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h159ca93885a3eb9c163ea500c3fd88e80ddd18fd68c454ae2e433b54017bc08c824200ea37298a8606912871f85d8ae5d6522d4de4cde9e0661b5fee352d5ae4c8219c0a1b69ec8a3694339f287e7e714098057f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d1a2f38f0cd99705626c9645fba7af28c8cad59685531c676dab98b195669aa527683e03f7ea2d7d87c2c5363f66b8a33ffece135a118ef8dca5b5426898ec497dd6b7064d0200e6d378b82cbc5c0ddd96660f1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3219acec4b22c2ae59b54cf53e1ae0af4ce2950643810576ddafd3b491a4d06456284299f852dd4fdfad2d96c7f64641819181c3bdfec977d24843c216df11fe2f25a236a2dc7dba6ee494546d7f4d844b8f9ab9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d6eb15a3741e650639f8ffa432f5ac7d978ef10e0f7262b232623d505859443fd987e03a3ff847070853ae91cfcdd1aaba5d9e93567274e8e6ed769d092f3e04c9c38024fbce7797d1d58740c599534c3fe40a34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74796642775c9b37bad3290f5c16b78c4bf16dee7828fb5b92507c4612837f6549754c53d9e60d3171e3dcee8dbed5a343e14e7fd00a970c6ce5b5a894bb12ab5cc0ced06ff8cc0363024a8959f0810495b8c1cf2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fc270da5dd3585a04a9c960693ba44aa23594821a151dfeec0a9321cfc772c8fba851d7f97684937c6b3de22fcd66b8579e7545d6c89732e62ffee3274e40890e9c744917791ae2d2d6a1dc92b76576a98a85882;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3619e1ad81d108e812ffe0365f55ca4639e1ff7b1e5990eac1e36641c1a6b785c0957dcadfc6d9cb497427f8471afcfbde571a42121de63464f9675f780e6edcfb671edd6f12ded06240505a74e43da75d8f752f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49abe92ba97d840d147d431634142192c78c0223512575b0518d906a235573f7d02c20ca105cc21d12ba43586380ade726e1357b1e662bbb7e260765ed0b0ba8bbe31eab45d274be9b36768127702898c15405f9b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34da9fd6dadd8f6d758ce1ac96e31a4868ac782e940a121cea820ed99f192e618713a4114a6f7734852f8a086248e662ce68002997b608e2391a6a4d784c5e2c8b12f74e9f6d24eb159611e0beea7e1a3c218b8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35760bb66b86963d623c315bf66a8d3578d2e26f2398cc93e00bc99fa66a75dc7bc4d70a519b16cb66adab28bbd709bc4dc2e990d32279c599c5506fc7a08bfd4a355f8abed0a1b6f20a61f179312db66ce5feaa0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40f7aab34115846a1cd9dc5dc8ddf9be9c6eead039fe883fbe24155adf2f17601308d80c7c098ea8634d8b6ae08ad52c9793d5652a6e2a698c08c9a93c935c5043fc05f97e4b9beccca8f2cbf14bf620dfdf5a838;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74401b8ac2820f6ed17cafebe0840e786f5a60184ede146011f39d238f1b62503b56c306d36c42b73c494ee8267c4964459fa6ef43ae6e722107c7cba190b6be5166a308d781dffbfb68d387522be59927f008692;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1f0709d427190b0f6813aa9e5b509dbb0de62a880df68d51a566d338d3956427f154d226536cb4066f9c4a450d1bb3dc27e4a9d51738144cf77b732ae98f9d8e02afa32321680e268d7df190e1c95f8e674465fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a14f54702b384d8f4229f0f5136e75c4143110e6ede0300f2ff27f894d0b57c65c011a820216cc2065e75f415fffb3b66170141ab6ef57c8cb08d101a80b3c6647e983b0069f465425b641328f25e8a4b9f56f09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f51856f0f211b64b27fa39a3462796e45e4384074eb1eb771820d100e84d3f48e370b4c3cddc2ef918d546c80aaa898ab6275cbc8f72f9215e96deb5823e63d7443834ba391829e1bb4053654ec03b6bd2a8526c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80c8f8dacef0f9f5458bda9ba8f53164e96388d499f885a69e034f64c2bc71c3bbec2361240e7446e2df4c06d60b9e99be46637650f67633248aa98e91dcd9aee7efe6d30c3ccbfcc342c09a3bc7f1db07bfc3d09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f0e7bf714453b38e8d71409840075d89e3a95870b136f93a04143e14b878f16ace819eb4803337fa97e0bd6f81835ce3a4652be53d71041c686b57daac2b1f2267f71a7e83649c4621f31f7e0bb2236befda3699;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57f9f6d0c7b222512b794a6a786a20a2c8d81c2191c49d9363a2ef51eb1fe778b46c50aabb69cc4b930e714a179ca4dcdf585ed86149e1f8c1912554899679ea9c8ea02ab34601b01531404086a3a365f7f09607;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b5782bb1548a530b68bd68c049dff4ec97392d840bb7c2db7ff8c74a91f4b6ff66d6232bb8e9349208836dc386b6cbbe7ae32c907d038f5db4199eedda07e393b3e1a9b31a76c502e4c08c4b5335dc41fd3d19b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haeadbdb146f3b45c2da49f6137683ffebbf7fbff68580b86017c847aafb845d25526dc6ce9ea82e485ea104eb215a42f9d7a73b494dca19f5de4f8cd6292504e00c8a49db17b47fa0996b8015eb05c1a4a15547d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c2d316bdab8e82726942e35f43f3c13327341761804ac6d3022f659dd6f4f2581131fc43d5cc2c3b1253c017e24f37b10f0064d4679d17ca73dead81a2faf5d8ec8141812e627d57a5121add0c285d7fa3f568f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfcbb05b22283cd4cdbaf69138666a2ff7317b36ed77a86b8ddd8a8fb8a41e823f222b737e448adaa6aedb71c3c97e51964b22ab1f8f6a2298f275d3d513ab2aa7feb921e8e454864d4136966121c75fc22f07d6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc177d0be9e5c41b44945e3a0f58b5a41c7460c8b0b3a9c44d0e58d6ab8be370c18dcfee8ce87c3207b1f1fbff280c18a14faedfce074f7d4842066845af917e20df443093fd05215f6d2adabb728a43a5a626e31b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf878de846997a234117df6b913567b46bb69afeab0a85cca500c42ae4e8a621d1e36540a461b2add62272befc09429a0035cafbaef2a401d08f7ceee56d3151974c31c4f466c7c64b5d1c63b2764789bdae480107;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb01dc6b8b0469a1764322d815861a8d7c0a7cd0f2c2894655a8fc146c28eb37b569c913b1edbb54fbc23abd0301d2da04893c6717a09e3f2036f22535ad2333de5e5133141eb9acec9a090083d593e391e9c5d9b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf633c0845b4fd5c5c177edc1333679351de4190dbe30f4faa93efa7777bab7901870d7588d6a8fbf5f1e55f88e821b655a0432b0e30907f01ea3c6f235f5248a87bee5128a703d3158f4c04d6a75f074b8d32e89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52596763bfa45db4913d77ea8364ecf621a7c9498afe764d89a05703d0c44ad759dc59ba0dc25329df4c498905547baa70943adbd2ae72221d29b723d380948ca14b682b53c1e18c9b7aa039cd74932f85b0f12d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h536aa8ff2640e8f82c3624f25378e83b7506cafabb5c6264967d8d21fb4d4f3a4b9d0d7d51042f4dd1ab9320eca250f114f4b0da9ec88fe98e34da24aaf7030910026e9adbb0f05893d694c6cd68e1f487a57970e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf55b8589e5b1af682b545c526c45a12688797622e07a1759087261f652937d7429f03c7976a15406a78e3358496bb0737d933d9c8259f9e2cff906dac63b2999a7ef57c62f85c5ae15efcea754be6a7a814fbbeac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9e0f0780a980c8895f14fa724826c788a74ab93c792f30bd31cd64232095051fa9a204d60e54f8c9d2f9e1831549f63ccd6b667edb1d042961839a31132f94d535dfdb48238add9b216f846ad748916ca99c2226;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6070440c9fda9d3beac4ec2cb269ebb9de698b0819639756558fd71ee437b1258484e2237fd0ed5ca35f8b80dfae9e88b7c414add3b1c96aec358dedd0174c74d3a12a5e3d7ae9c4a740b128966a2c1f3c82ca850;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24a8ef4ebd72faafb63065dc7a1c48e3ed6639d972092846ad3dc56553e5e7027e750a3374540ef6def09721e1ff1506d38390d0a3c877b758953a4970f9a9aee0f4d6e54139a9d64e43438fc719a28e1cc616806;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82b81eadb2d2b3e7ed1a02316bf424d703863156105fce18d397d7890981b2125db6cdeced0b75a2a838ab06479b95093865ab9416604547d882c0615048991f56895a3c4b675fd0a0e77ded85aec72767d6d30f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f5ad38a5e473fa660fc86a52e912e768a3acd4438ceab3dd156ff3aa13dfdff926d181d23561b0dc1bb6f9c066619b8c1bb3fe85796ec1e2c92544b9f2b83ef84efdc4971c02cd32871d314fd1c5bb7e55a1a39c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1b2490fcc83eec56a776150b1f4a280f6397581cf9e35392ce5a776b5bd0bb936f5ec103ca7f6d6465e6585a805f06c003032cab5401cbce490612d6d91c9df4adc8718ebdf6f16bd666232ed289cd80e08f9251;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha31e308554625c03ca4592c814e4fad374926f9d54749299afd87a9aac6e205bb0699f1b370dbb35fc43e5ebca576d24d366ab7f1f2cee0f94532c523f51eeb2e1913c062d84fce82298ac710b4fa53dc3e5db026;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdacf124a75314159e3dd51c2aa03662c772c855fbefadd0a729d355e0bb60432b8e9b930a5cdcad56b300be6b794444ff8e8bc1f7e3cb04768f91871eb026c4015e85bc26079724cef1a2a2e579a45e80a3688862;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4965a1ed00bc15ab2577f77aedb52ccc91eb6a6e9e6fce9f0077a39953f3c85650249afe4786476d4ebff322379108b3fae5ce0d281e67aaecdd48b2cd449ba7897f2c0d1e7c80b432ae74edd0d598083c54dfafe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9321149b00f10a494ba0b875085f06bc5b872c89c067d9fd5562e7820349d51cf15b22eaf82167f0759f383ea42de1195f6f073153cadc577ce17e697b2c3b450d44b6769de948e685f17e57c2810ccf22a12d93d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95c7d278e33c83acd4941029966338139ee2ac536dd8af018f65ce50979abaad023816a68e48a1ce05ced8fbb8fb7972b30a9183c03dcf2d231a8472cab25e365a382589237d4287a7af1d728352f5c7b19d97d69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80b3c0fc664204df22ce4949ad42586105232ff1421096a00a45e313b9a72d6b0fc74d7214e8d708033e7b5375d0362614089f7f637e9f92db2cb6192c3bc5db358701d7d2cbb795f261b54f8722934570e075839;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca777388a0edecd5b790bcdb8481e037a368e82a2f54a791ba20e62986796307e9867e81629860e5970a692c6d757e38ff6875b0dbf4dce59317b617020f44ff364622a07295546eb76a09be72020d846cc617470;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb35dc272743f7656900ad3821e7f974dfbd691daf16ea62fc5ffa1369cb84c901efe59b3bdfe59ba66d82f2e258a3c4f537a84fb4872385f7dedba7c2edbe28384496c433186f655afb0712be3cc26812a55a5514;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h679a88ca56eed6a95a7bb0207cbd63c6dbb11e3d03d8316582ec3f29b688659e64cc75dfdf483c1ded127513cb689ae938881eb9894cfc814455510815f4feed94a0ad2c6420842d6adb0906382cd2b711939d1ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9982de4547ff2822a08af784646bf9003982c3745254641492d971e8f1758e5ca1080d6c25ca3fc19a508abe212a072875f00b125554b39aa28a0c13cad536939648bf18e80c6478c3a7e6b582c76775ee5d75f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8766641b2f4770892c5b938c6479fbeff828144c259fa35de3ac0d9fbebea25ebf6ad445ce7a944560dd3cdd54b3232bfd1276f9a8c5d4b9c9e3f13c29693d38bc76e4d2fe01e701d423ae4fc48b6facefb54100e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe3070f0749e67a8c3fafdcffe5817dae18b32c47d201c6fb35a04a16bda7cfd5052846af3bfdf2725772a46855432b16a6a51aef8ed11fd2acb263454d9832ba555c3f154a68c7d1a0d46403c26641b1cd073145;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6eeaf8b1f5672c8b0f95f823f6bfe05aedbf34ed81f4b8836c10d9ce8ce4e32570c6e3cff10e3ce1cd26a18501cd020571ab0b266b1b62e46fc02b10f8a296683e03eb9cc3cc11bec5aa93ba642433a62ea3a6b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5dd30ac992da5e4a8aca277a8d8afaeef150381fdadf9fc0fd41884da17d461f946ce36a4d46e11a6beb58d51c6248001a8f2625eb59e33dc500284738c4991ec420e83dd5af2103b68615fe60002ab4b3ca51ac0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e8696c4f309d55d404822ef85f74097a502946bb8655adef5ab708608c0987438ffd929208fe12a02c89047232d09a5ae6c48cac9c93935190b0b877b6ce866fe9152a3547b8c74db6fc88b6e4aa662b5fd7443;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4edad1ca09567540ec074824608ff03e9d16c622cb47dc80e5fc08cb772dea0f23d5793276c940c9d69a5bb29c11b93f4f8a2a970dd04f6fc1541741e79a849d1347ad51fba4bb7b724094d1b106d8bc6fdd005b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff31dc843e657a7520423ba5d959cf2ccd9eb7435bd1f549754c7ac827ba89867d99e15470a404ed64f0e43e0790f14417fb0822cee1cd9cfb34762f4d707c57d9fc9d2c2f9557cfb1e1d3ef0f246be1c1eeb5fca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc78e34145e4e742f35919fabde1c73b4807510a767a8c350b37f9ebea192a2df4067751f19f91c95d8b3303d9efa5d25ad3e9aa3adf541fe768eb72b45b6f650c6c5416f7265fb9bf3f1756f7f315dc3f439738f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab161781d5ba5e1e87b43325be7387d058d5ec89e1aa9b0c4b8a74d2404478acf99cee4824eda2adcb0c33b3624863f78d0181b7f6eca63aa5c780550798a528aa34f7fa96582ea0761457dd8b87deecaa06be944;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5d7c846e5de6ad107da58d0fcf686e42c0d904b1f2c44e8dfa66680b273f69ee1413be302007ef3035be38134393f5cd0d2020b1527c286ed19523c531206241427cf9c4426f26cec523732a66d543e3bc185a1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h687d465178b862af25ea0e1f48b30607866cb8abcdab758605b9250e1facb1e35df6d061dd121133bb961584c116180f0660b4d564d853373526b63c6635768e47bb0e531dd658605e3cb3a9288e64837061940ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc908adf6ca5d05602295d70a9dc3a3c402e1fdf8eced6cc57d3a3e9f505c19a19cf978a129274845fbc4667ba73b7c61e46c2ab3e68a4e3fe7fda09b0327b2452b201938db5400f48c5b42e042315c787b4f3914;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h865751a56232322125f67d6661d657b2342c9c88141eb7928ea1122406af58e52d92e39ff2a6f499ed273a177e9fa803d93b333e6612b56fdeb6ecefa74669554ef570d80b7c356c16d9e6114c10cdc1b2f5ec87a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h985c98a753caa8072958c2d7c2463a9ffca587534dce1043b4ce6065e8716466e011927461de57ad78093f87098db144d067eec7494503db962498e21849174d035a9f1308de997f701ed68822ccaeba1a118e4f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e409232fc9170bc6fca0dacd703b667205904c115174578993c264ac42bbf085b1cd9a7d18cad6db04470cd0d813067399d4130f182dfcc4cc660f240ed720b177908922a78cfe5ce63edf4d232b34628a2b7f60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3741bf8496afd4a16c65a62e33e6cdabef8c8c90481b32595aa9f1e2b39b3d157918228020b6d13882d7b3d9f22798ed4d199a4c75c93dc5df600b776191246e937abb9cd2f437562fb9e25bad3c9aac43281074c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2eaba1af21fe4dac1245a1c3552fe50a94154abcc11c9f2b71fb754e4242e0f268b6a1f7e0844b4aa80e9bd31b85caada6d07e4ff0313913ffbf927c0b80ff2e1ae08a64276f040d6b51ab7f0a6270bc084fc0c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc2a6c6e0a7e26861ae9816dad7857cec80353b60a770fa525b0fd8be75c95b4d9630cc138c1839dac8da9b005fc7fa5ad26fc46a570369b94de87e6000f9063d8e836398be49932424268617aa86fe10a1245c9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b67752aa2326a245aad6077704cf41478e307ebd816fd081c7c841a3e1adcc396c7cc2ab6bed940824ac1323eefa5515b9943ab44f8470ab845209a2fa60fd4c6d0443be7708f521a08a5c019da9736fdab72afe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he32b543211ba8e1cd58682178e25c6929ba35804587485a59c1053ef5d339a9b3b4bdfac4361ea9f2c86b2c53a0ae3ff1c4d1d5a8636483555f2eb585421025e8c894bed7dad66624be0793e7a5c624e7106a415c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33dbb47936fc81305c06db1b5eb0e8bfad9fc489843d15264adf5aff0c02f04ba217e416df7f6bfc6976d5b34c8c2c09a3090727e038c1caff7c432c8c44068c3cdf45ada0953bb5fde3c8b4e4ae4cd6fe816e80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a02ddb349a88401c69b2540415550d68a42720d53fe8c6413ec40d2c38fc964aaf3d57e3cdd230f6341fb7990b9fc24befb150e18e10dd5e0b7d50b3007b5513db5b3d90713836a54384a86bde30427bb07675ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd46438278007fdeb0a88696b4569ea7428c14c5bec69ee2c316643a96c70cb954ec4bf203334e4846d04929a41078a3f9d8569880a4e7fadfc01874b53147ffd84e934deda7627b3f3513b8facd5bfa1aa7b20b90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6a90c76e1c946d839529e17c80161d6b4218a438128c028144003a7c6ceb1f56572456b43cd74a5f6e9afaaf72d70f55e91da7ee9bafaa4734b089f0aa5c3de0e6de38106e98c35460abb4922f5f589bc2e24081;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb48407ce709a5837c79ff816d2a648cc446830ca218a480df8a99472109610ad81839939b9868711c04894369daa0b9cf10a0d8bf946daa013c085e0011391eedf3e0f8cd7ff33290774e7fc27f38218c50b220aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7292d7e64b9de23d226774c3f6e70928d45701558580e8f5d6656c1f5c5a6b163dd41f20fd1e6900c05878cd538186d3fb16874fecfc9b53364b1a2fff7ae4d1a3d491af655a0b8ee5fa62816647eb277d7e98305;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ca28cc5d5c0fd45eb615d4db03f719b3d8cf79aba330945d93e2e4d2bc4fb5f78c31035a63d1fcc4530e214cf3a35d8c6b81d949117e830a8bd5bd730de63ed153b5cada37ca9c282f3426a4e4d70d35afff8fe1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he66daa601e8e128f6fc21474e93e7083daccf889ae6f6f0ed6745f2bf61de3435fc778015e8e6764490e680128a49fc4660587a5b2a40b837a3748193c7cc2d2a160a8045444ff6bbcca5b94dd658818213aa6429;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6114a8ee1ccfc9404e0ec453f3518f554e2ee954e2b21a61026a00778be12d9553c78bba8f40b90b90274fefd2bc0710ef9800b34930d7b51244fcb5d9aad410193eb59356c5ff4e21336ab0191bfec0179a416f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9db8fa8756a62150243296ea6e10a26ff0b5df9876126fe2df3da3dea29111756ff4aef6d84e309234f43456840e0435e74a0ce3abf4d6a1c39eeb4ca119b3cf17139db4b60ea0e8e60756b6741419432e9c9edf7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7333dc673232f34781ad72575ae98d338b20921c9717499e1e7a3e86a8bf27ffdd9b2a85e65339c95c818406390c10ad8fa5ed84b2e507acd55d8dc6b070476ea18eba145a471f3fbdf6ec732b6fe15d46989dbc6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25f598b88499da09fd3aaabbf54f719c4707b39f7977e43bad4e9292c476c3b14a84babc9115b9c1377fe94102b01f483b1b1d729fbf8405601cae2c52a91255e6a5b4be03556dc118b804924363885f86cc97e7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70de2c5472b798786b459beab47ac7834934091d22b9fc8bbca36e0aa8994b9b097499bcd7296b7394b528ec674d6871f7596bf0f09abf4a65f8b2022dffc61943262d08555afb758104f7702ae98fbf6d89246fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63518d20200106121c00977ed958e709102c41617489a2a19859e07f57401a830893a05cc028c3447a85b1b2b33e46556c93daf2e37ddf9622abb4189ef0b82aaba4d2077d5b971fe9f60d26deb421e8f4c70cda6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h200735588e87798663eddb861b1b8c3a133cd10c89bcbcfbc0fbd8d82e8dc24756b1653f7a207ce057df6ec9aeb251d17485c5ea648b2082e34685198a1c9553836af85bf4822435652e5583e65658e5aebec1455;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd727436c9bd42fba3b71a1f828dd11891705f41d238113f1b48eab314d8259520c6233b655c7ab543da4aa910e9bfb4e635089edb399b58c10504026a79061a62ffd657677e59b2aac7e2932cda0d4538036749c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaa89da841cb29418244ec9d13af465c14bdfe724c66773ec422f511eeb4ab6055f7e4a82c3a96d29989a6a397a3f2e32100216ab65655a0410802143f68970ac74677f2327b98ac8b3d03b09221a383ecf91dba6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h551641ae4e59f485adad3455d7e08f841722ebb05adbc84f0331a0188458a4273d14f348c8876fba16dc3879546095a4436246b49025c3a877118a5cd5ec0af9ee52d1e9fc2061a777a1a1eaafdda3bd9dd87a390;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3dba81929e59c4129742dcd4362e7cab50d0f668fa6a1119fcbe0a6af0fabbf6cf25d7f5bc35aa58a33f217735101a45bf5dc09ac20435d6fd7145ad1167ff750db38a1197411f572dad6b96128425e69a879849;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa75d94b3ee7205ed56c95ded05c8e6b4df7bc5da1d7b0d195c4839f131d8666d95133f8e2d00e06be49f6f67acfd469f5dbdeaaef2d79ab5769329fa2a12cba580315dfad8e09e4c8ed9e43a0002b4304094238b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd96dd0038538f1bf753d261fde5c10d31b5add7286089c67f177b3d1c826adf46aff9e9632142b66a2389a37e9aa44dc8fbe4a7cb1ecd326f87d00697b042bf2d0ca1fb1062a398dab74ef9723b5a2a2647214751;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4ee74d7e2ed3d5e91f498e2ccfaa6bd776b2b2e73d5493ffdbc12a9bcde1339adfa26e9a4a32794a5ba970f7b44ef6e2a6f8b309bbc213a884a43e0af1f296a8eaa16963236700a7b96f51ef830a09ff090c744c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc67af4c5bd0d6ab6ecb1d254c7b48f8e266bd5d4a850147e6a1aa97a055c1a9dc7600bf8290e110cf98a1970a6cfc1268b24ca27f92a290f838239a24f65d7253f08feeb0b4a4918dc0cc8668e889d974746ed02f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4af494955511ad8c2c00d6ea2ab379f528bb90f1f6267b93096d03f45faf867698f25febc59bb58e46b2a6e8836a2fd1f2addeca624a3fb82396d7c704a3bc0136985e4fcbfd5e7dd75d481cb7389f13fa7a50ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8933c2d0bf165d8e0372db62d38c1823ac1ae51df5c88949418503d313a172931df7d882fc839093d26b92b21fbfe33a7f0534c9f94b17002cfe3b3743637a2523088f492d69d7d020c053d64b4472d13be05dc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f8fc38e1c4e473c56848aa35071e2a9f1aea8058573512b01fed842225d3327a716e894dabb3697a51659d6d0891ad1749d929ba0cee7a88d8da3bac693feb559c8028dd8d95a88257ab3925c2d43bdb10c14d25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef3ee4a6154ad54d3160cb63e053d54e7c35f978c51943e91e110577d505d733fe4767446351cafa6dd606f5a86ed56801422c9b4ba982705b9f72f10e4bb2241bd4c22a4caa374f48776738befeab0574c738194;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42b9c4608eccc81c7225b3e03bddf2fead6cb97d995af2be0e5836765500b4e17bbb6440c60d96e69342d62419f67687f2a3f356ee0f1a3b47a2de7f4f83797ecf84719321190cda1c7ae64d7cc43aab9c33f6ceb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ec4fd8e2af0c720c12cce02900a12c0646e5758e8041aaff1827db154dc8b12b092c1f1cae08ebbfad3c6304fbfdc94fc80cb776e29437f38aeb5a31da2b858e9ed3739b8ef8941286ad6e4ddc7b29dab7f34f1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ab4ee25712e0dc8b239a8165e679484310927655adab44db87d20ca65a30a9b122b7c14adbe456059a55ccdbf11000915ff938a60266f6d2bc1b35d567eca6a6709707dc78f378ee4d066fe73af0a03af1db28cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he673d9eef21abb5c155c15151b8871cf8dd6be0c3afc82ebe8e0be529a58dfb4cb3d93158e1bbe0d33734e66846a21d7bbb7f23ee9c98ad57ebea562eed311bfc510c2b768449945aa53bfba2d470329388428602;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fa36a01c6fc5ccf5483379065ff2c3968ba466d61a6c4293baadb36a40a966fa65096d3a9b38c296a8cfaacc77cbca08c6e6fe08e593c05e49b0a7e27b2bb17eef0300624466cb68beba79171b3758798a084228;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d315545fdac9ce12d1a30709f38e66634a4863b7d46d1a5aab3533688da352ca0c70989fd2660a35414eaa383baec514e5e9b984d37f8f69aff02925af165910178ca5f4aa5214766662e069932e79d616ff6fbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fafcda49779be90f770640eb012f9164cca74ee4c640c3f04d560140b64fcccf08eafc6034b45f2b685b7b8d123dbe0204e9b4f615ebb2539469885163e1a8e644b92afa377e51db2300fc97ba91eec65b02b4bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5d90476ad0883c4cdcd49483c15db88bfb58656009293f1be57f025eb70a8adac405ec05483ac8e8dd578ee85774d9f5ba11a65120eb882af11402b8654db3cc98c04e57364aa60c31b14ec9c390e6b23df0338d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86da8387cf95417e96f7e6b234b44a6e731e420acc9feb24c5a1c6d189f90e8705e10cd6f3548ae40923301e271fe64b481039814280224df6ec8ba591fd950532d92fc3b77a0b9b51965232c0582102a0d0c86c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94e1ee448c5ae58f6b6783a9cedfc5853514e5e18d997585370f11e09e66d0845bfeeefad238bd3a2f2498e14054a2b3e9857f85884f0a4198755d76acfb9a4fdcf04b77b7acab1510db8741d00a136a68a2277b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hceca6ac8b8736c985db18be8d4071f87c5ad66436ed3da5468c12bd8e22d856bb02bc3eafda89f7ca43e653d47aee6af5be7f9b75a92deea01dbd3763bbcbaf62a8f415791492703027589dd6ee5e410c0736ae67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc881c7065fb3c033f135bcdca8cb97294bbf21ce733a3e0881eda9afd6580db5543e636db3ba5f86906513462fb3d854133428eb06362b2377da19b1deffc40c976cf01400d59b75f0e91715df4cddd3ab5d4b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he354431a81c980cd4ab700bfd2a83759238b20c33124698668e7b20bd20c5281e2d6efb80925e4ae7550e815336f2daea012ee9820bdf47b9eb65e7fc7fb2a51c986e9b463dcbe7876588c1f9c1cd8230aa83453d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h254db4c534aed87b4fb9bc8c226d9f99b6db68a92a09057add1984b08fff807a127903046c7bca90a566954ec6d5c702cccba02273ac6d00f5adecb8f3047d1778843c115c25d7fa9747fb7007252fc5746d2f7de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41bfddf28aa6996ca605e6f89da00a02d2c1b0d0b183a44ddd1379a42592f272b3ee251f099c43290859d4d0dfcec7b300cd798262c2bb6d30574de9cc9c76e2521d2df21e6704a40397bab69f927f54fd67028c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b54dd8c8c57e578ceb7287e5a53251a96f23773020f7f904971923eed00d1dd64c3f13fe52cec1384f4cb8436ab99f380404664084738d35ed428f6445506f054ad57d73ef71aa69244e3fe2ad6f92ce11edf7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f7c0acebcbc9738d14117e7e9d56b3f2815cb3d72c10656c63a6da033aa1aa80165449f48e6500b2c4a603d501b5e86cbc07e71e64fd03b960691e4ad672367a6fc398084fc7a5095408b4ba7edd7e4158ec9df9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7925e26e0a10b9e6a45ad6b880f4c1ba8cc628c1446a17aa9b8b4a4a074250210b31b510eea6179debe4dce8c04d8425f1ba1410e9a6be40dca00390aa5e4afcd721f6c95f5a86b6b0b6899b47c4c3530bcf69019;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e18addc1b2db79ecc79bc4fccd3370cfe0d28a72d2de4ded82c30b4e926366d21fe54618870529cc5607d80485e780d756c84d4848460597d3d76f9da5896737bd65ef4ae86b1afaa4b9166b7268be299fe7c8bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99a6060b19820b0249133499d963da5d32e416ee8a6219d45d302d091091372dc009d2a395f2f9db40ff47ed12ec0efd4f74f8000c5b5d469127274059b8a97f10bb7585b194f7216d21a18abffb33248168268c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74d694d4d1bab6073c73e8e2acf0b89d907346c89c7c8a265ff065399cca260c8855a00968864fc39f99e518f901abb3ff0f355dd929f6322226c8b8ecf68cc72e8fc5b72ea4f0be7d0dd6ee19cb92c5fd90bc696;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5df4c5c9e19ce661e4c0de47e525accace99ff2a11521d46be1c0bfb1b0b290190584bb884d06026a6fe0f336d3cc3b877ff1875cae76b650455ffc053ecdc4deb3a2e6bf9228e8568866c66d9df5c478bfb64ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41735d3928659a882ba3475f64694e65102f270c6e7d0f436fe1d3a6d335b9f24e5df5679150bc78404b3c7a50fcd81b7769bc6f48bd5dac7e061d4df560e10928cf55ea24db1089c5afa1d3950fd64c205f5e76f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacc808084f8f20896e5bb4eb6c58292026d3d9d5a0097cc595abb1d69b15bfd712d9bd80f5e774cdf06a252568ae12b1283683f87813aa9b4c184abf0d91a9fe671fd99835ad1d3f4c3360cb41c1344d95f1ddec8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d03ee07bfd17ac1e0b3306cb65c888397770cc59c86def6112529e48e757be7024b18dfe1151f7e02de82d8b1b4435cf2f029261d405781f5df71a114e46a25ac98953f769a3a07215fbea8e5357abbeb08fe4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb91071f1452713a2be32ae2c25906c0061bb0599b9946d3486ceb9ec6a7b051d480171e24d58c591079fa4254a6f7aad6116dd9d63f41f91d79a98b457e77f9aace34204946d2841f83224504bbd6f0e0881a608a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab157e9162ed27def4aeddfd5643ac7a6af55cb5c67785103a477eb8bfc5854fc7ba2e23477b89e87c8ed988565b843ec4385df11d98aea657dee699d5d3f584ebc0adcdd9c220da34ce320cba238513180f2d44c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2836199503134a213b022f6850fc946c0bf01104e839451d3ab489f0e5827f11939c4dd36ede38e2c65b27b69d8f5ae2ceca65fb81ddc092d221ec1e3f07d9410f315eb3124c8c232ac017d2bcf30b240746c61c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50e573e91867339e210814821afcbb8c080056c50e54a9c0c154e728334b9862b75b5cd11a9604050c5b71d11478eae5dc33b7c39ccdfafcce8419d7b11399e0529f677591586ddfb27536650accb3afce71d04a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb26f14c4cac1f2fdf260378c2dff752ee9d805c8d5e12308aa74b5157913d305681379b1608fe1880a7864c739ca202017343f8f89fa479e126da36cf915365249c5341ffee27178426c9b7a79844139fe2a3f2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4aae8ef155888940742e92d270b5c5a02bb3b9d39bff43a551100481e4f745332cb3c7e8beae76245a0bb535c3c368251bfec821f5f1aeaf69e8ec098331a1f2917aa9290b366399ccc7d93498574c08d93f0d97;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc867e03979a15fba3e694e86e38b8f61cb8761de0ceb9f481fd98bf638af111cb50b6d2f6378d72afb8b012305804aa9a2b9dfb7ff7482c834eb98c9bcd057e6e34d77056c089c1cf7256a5ed0d0fe5d775023557;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haee6890242bf68bd150d829d5b01818144cd24f53e775e3bde8dfa5a5424156acac0aca19091097b7a519e37e98055553a1c2dfc52c7c430ff358f4700ebbc6fcf3895a6c5d3bf6910bb8f7ae3c2e847da99b1036;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4efd19e926479d50ac89bc0b939c89ad5a1b9024c207d3d13294a82346126a2ec02e96903f1dcd1dee4984e1855e6caf8d7fc63ffbf086dd289364f82144b3f1e7784b61af7545fa2a2ad09fd658856e5b125d02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64c96ff0310c59ac543127dac6d22cfe683b5b6426886284b555d306f6a6269c5dc598ed43437faac346b7d7ab710866c4dd4f7bbd0d70877d32040592a99d239f7f21657bb6f787f2be290fb4d316c1ec229bba3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha74308a9c2a9931241d131beac80d685d1208a89b88bedbf8861efeb90b5c9c0c3f4b9b2b91d3ffcfc6dcd0f2f4f445257efd491a68d163c4e74f0f055251dee4e86d61e3776ad36a2c2110461f8e64500bf49bc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b97b479a2135bdefde8d83b53b33e643aada197c7c25fe08a57076f380904cf0884bedcf32acf22f8da27637af51e56906cfa8ca6655284f58f23875ffe4420a3f9a159e8cddfdc16c1986d14a57505acea27431;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h773149e159bb15ded810c8d73fdd765300410cdafbe293203c8d9759a136d88c46706bbb2e87bf00e87fb855a723a96e96d89f548fcb9ea3bfad556725302e2c90633e06d886adcfacfb48ca9e3b281a0cf4f3c70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef0db426ca467c494e6cea6cc5e7e868883c8af8089b47c35a250cd48694ad2cb74b74cc31f55e86ffa34f95a300f43088124ec759047be6bae8370e9edc4d2bee3cb3b354184b61c170ec1d13f196dab8a3a36df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4765416eca7b7366dd7927f3b50dfd8189819f7e64b0f5ccdb8700352648d80656aeddf351ff03fbd327f2b866971abb331f20d553886af5da6793d64652e329631f91b9bc0fb154c133eafc1e2dfa378ebd8e3ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h216d9cd91dc459b985cc45fc334ef35fb48870bca8316cd176d4ec574b948f3811b6b1634f75e4a26880ee69fab74e1271193978e0498e7993771471dd7c44f4a474067acfaefb60263b9af7ab46a0e3e693355b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haddd9cb4a24dbd49624ce317fc4e9b143ada0d81139180de8d405c5d4ba28f56914e8b209af474ac7331613cac516a0ce012e072bc8e6f45accc9d9ebc130aa80c50135881e425a36fc79f8694ac2a92c4bda4e14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a53a38132ffe855b965c3ffae19134dba34b4be42626644c50fb98755e40f5b963eb9d1896314746481736f5bb4a9a4557ed78b45321e44d93e1ab50abc5ffd0247ea2f184e2d6364491307de14694687feee10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h456a2ecae87d29ea80f94d6372f8e78b55fd8d75bc0a2a5f140ea202d3f864b9c855ac4401680e26af8bcd54f0f28c2b885cb730eca7de0c9c4b3a25db4be970669ec233c38be54e67cf1a6d7ace1bcc016e0183b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a2125ae89dda6ba0d7263f6cc071344f1fed229c20f55a50e4674132531b158bc1a46c382041afed9ee18a35f4660682ad089e8276642e94fa7c248a2381e1134ec32d3925cb289bd7a8175ef9226f8cbc5ee22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9839079018969bba78f48e0d90ea749e66ab8c92854e382422437ea45fe29a35f9ba33ebdb0b4d764b52e7aab0f34d7a4adca6d190c1e9f08f9d3a222d174fb69e05955cc4a80605aaf6a42255c18571123ad19fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61c06c9aac2c79677df37b86375e70d3dd4dcfdcdb30b110bc18dcd4e1f3467030c313dba3af73fb02c0287adf5287b7e94eb78db775644c69234a27951fb7a33703e3d04d8677276a34459157d2e40e0ee0708dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc6a9469fb0d4674951300f29aff4d184cdf70aa70cb05b8f153157a6091a2ff12c0e728f00733a486190035158c297373fcb2807e57a5027f7c69befccec40649671f159f08b6c66d689c64e1cc7d13d79c9e564;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f511f7eeccfa1bf204b78fe0325cc924890069120778db7469267f5029bb3c4f69ebf29202219e72cdb5d6f88169047b65061b00ba06c857a26918cab4909e7a2970ae4374cddf73828d667aa91cca34a97bf7f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda8e40531e32a7fd324e5bc4aa6ac6da87cfa6f0cd532a751d6525f7772718e2edbcd0c1bef8efd504a89ffce39adc6b7dfb53276c7ffadb7043ab8f2f9a148d90e133cea6a2e7ec39d73bf516f7ff28e32ba3786;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5cb949a375572f2591ea20c823c57baf85d067f99e8f3f36dd8a4c7c351af3dee90e496d8ae17660ea714e3d5f7e553c33f484273c9c140f68753a52fe1abc98d26a17a45a30b653a73a0a4d7b63b17247ab371;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h102f848cb57bdaad0a448e409160bda3c91aaf690db030b0ef5d5b565f51126f49af83804acf1a6d2cf2e1c3df50acce8669f913ee34f4fad751fc4121964f8f587ee2be7ba81adae6cfe5abaa0acb539709bf74f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddbf7a8b96649d4c2abb01ed1e3bfae2c07423350771ea138fa94fa4d4ab67923524d30ad1cb2d9b871074d049006ee2863fec77e820d06a7a600f4de9d8a36bbb99f95176546299a5407cd7d2385b6ab49921920;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h253032770938c42ed6186c1c42bb66b9f8f892827123452a6068a75b99d003ded750f017d0b0bab4b8a6ca9639b21151236fb0725935fc7473907bd4aff909cb67c298e902267a976992d60d2afd3977b5c163bca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he22f9e89b28a5c4596f49b86f904e228690f4edc71daf97c1c25898102c6a13ac2c29df772ff133e72c66c84294cc373740d035450803a0aa0d1796cab7b4c2a37f8613c321ddd937519495a081294949ba197e1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h517519b2558ec9c38eddbdd3add5f2c1e522d7e824b67d6a5b0dad9e6067918f233d064ca0dc88ea10bfafd7061a32af9c2ae473d0f0ec2423b1a9e37219ad1deb8b2a9c08f3d8c8af3512a721910a0cc49540dec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5080cddef0c5df8b3a8ce0216fd5e7df4396b55f1f0921e17c634565263fb2355bf7736b0b1890923f29a1fa6ff04767b067f69746195ac7227e2cdbac944fdb39d83347afa55483826cab3e0f57c73b7b389b49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe80518e1bc74ec0888036b9802a99240a619c7b16501c06f37ad13a8982aeb1c8728e4e699825c0ea4657ad8740748f2a8de5961e72819971d39664538b5dc1e0313373a1ad64766573195b1b6db280514256be6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f8cb15d2e567be0aed93eaca0a41c6d0139516e59ec6de835538fca90512fd7794b8f1d24ea2aa680a3734887ea2035809f1d39360cf62ba2a7144bf5ce5483b864fb53e73287bf8a3508b17b0b4935abbf2eb66;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5812ada57b425b1b4d27e5b4a3e2e9862c5dd0bea4cb6746e3973f011795ef3996a79ad3eecd80fbeb1ef5c5998586cd9be77f84243ec27c5c8b0c64a466ae3c75b4d5090b1ecbf7d2c7d727bf119629229aa9b6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c4444b309b43b804462391d24624b8cf8256974f6e9403219c719c9fdebf6d3ad86f13668e787e7cb142e257f3a3ea3a7014e99f63022fcd367024e662b18b393383764c5c5a89fab31e2257974cd03bdeab3cbd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haca077c5e362554306ed2410d7c293cba3c83d22f09db1876f2cfb46c2d1ac683165508bf08744c5dee95cbf330cec8608d95e5b0ce8c43aed4d70ab3d0ec708a6c11ec27fe67eb2c1d47f865623dcf8d39e089e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d9bf8983003868f78b40972d68ee5dc504c0d0f86c40fecbe843040b705b3d779a5b43fa6dc96fe45a56bd6fc821f4aa7144b30cd36f00fa9fafaa598dc302034909a9e94d882e0868e21ce79f8bf4f1dcb41fda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66a25b38159f45c4ca78734602ab49b3fe382c4193460be08252d376611fb2c7734d180dc5ed33fb27c400e3d1c1aad584d7197758f5ab639f499d865d4c1592958fdd635136424eb2ea3c63e1ccb2df8b46c97f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92bac096da08c62a80de00ee08b3b097a6e4a695a3331cd975299eb00261820342b4e76f4f0e3851597b142eb35aa90cb5f2717cfd47063e5a53542ebde7b51723c386ab25af368cd14ffdfa897619df2726c3097;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72a4105bd324b92bbf48b89a1b9caf1ea638b56583d933c1b48f890cfea086a022e149b2701cdd8d9b8d196424621a20e5bd0926138e30223042a3e89706dec8b632115dc0b47ce9f423db0ae825ef0f07aa23d1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3331e738768fa279008f9e38ed1320a61076c6255b620e66d9a544f58f58ebaca328bbc1ab4d2764b8f39825f334693c526219c612a5b37ba0e8d32829ff0a533f970e16f22bfcf137fdd626dead11624604a0344;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc40fb334b83caeba05970bfc2a1d040faf5bad3f59df18b0dfb01d35f5a4c7c9b46c089afc0b74a2fe38c6de2aa96d2951baca1dc61bb25c4d71891a50f469457065aeae8aff5ba9aa5dfd5d44148a1e6bbfab799;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80a875c0a72b5ed398a1da8d77eeb309f4d32ca47ba3646eca1b849d8b13dc051b0a7d23f38b91227de90b57f8aa6ba7e83d8d2b9feb5b81a86ed2ba34e55bbe5680e3feef1d96b87eb7e6e24639b7e6ec7d3890c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f355483c1d332e7953a4773373c5c8548de2343e1ad5e7353807ddf2660ecb606833fa3cba6ff60db8a3538b184e380b43fd14b9f04553a45703a691cf0f9976d5c62d5e8fe2456ceee419723d63b785aa83bf55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c8e58eb4c10a18836c451fe09f9e3e3d63ab71252793435f7fa86166b5858c432e65f5962d2bb4b37ca63a4f11071190d8cf502e4ff0a493a95593c6203d0badf7450835dbe5bd25e0e1f1c21a7fe17c26e33a73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef7cbf191ea65235c56ee065e7a0ae3a80a6dee5d3fef4d04f9a1fec24990940cf899152b72bc8bd094724170c1ba734893a4b5fc2e0bb2f862fd939acec050897a2a5163d451d66a7b7c84d9b8c4214294e2dea9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40afeb15122de833a0ccd4e2673920091ec3390f2b275c28f26bea06461b0fc1595fec8cf055f2cb4a58b8626da72971c4f6bdbabcd311786a9b6322fc0293c2a0a3dd76f1a3e91d935c6e3f61c8af2e902c4293a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e8786298b93af778d19e262db0763cdf084f09bf7d8829539aa68a7514019e712c49888cbd3d0e6f3e2af5756f5f6e1f6d5f62d7f8007a3591aec7b53756fdbd66315e753b3080227e4eabc2cbce00fe5c0746f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bbc28446942bfa10a31a1209873e90217c0b0059f6dfc91e645679ecbb94b2ef9c1ba14a9604c67552a8c4e15af6d043deb6b74f6d0170a06babbc865e8930e09ed7c831707d833fc06395f649509804cf2b1ad3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85a3d85e0ebc64612bf099d796f07ea6eca4c23c39edbe9549f6f10ae3733f140c23bfb1368480404725003608ba0745f0213f7065b613aba2dec3c4509c511d1b34356b6c487e5d82d3880c3656c4c03a833bc7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89c7b7817bafc2490abd1b0bfb36f4da7efbd1befd414a071822c3da8832181cdb58832056a82c7bb26d9c0d62161d36c089397cd9ecfeec854419273985eb5f43af8da2700f62df52ff89aac23ce30c83fb8ec18;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8169ae030fb0f2aa1d917680768941f7cd175dada1fa698be257b5dbae46c84d0b903bef4c3fda8a5ab52260ac99ba73069db61162272b7ea4917cd51dd1931e428d282fac08a2890f0d6692a30bf9ba522c38f2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h636957b991c488ed5de42bc803f3c07dd70b1cd3a316003d710798e86dd7347687363b049f519b673c85f9969ba5a09f175687015c7de124945760f6cd91dff00217b9a8ad86ff2dbb9eadc594d6756fde98573c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he41f4cc37a84a05fcd946dd93b08c00e9d91d7964b53a07d48a72cd2ca3a7df60f89a1aab01eaf21dabd1f58dc3e7fc40a8e20b79ef493a396cb03fd1ce038036ba84fd0d3b119599fb19c90f1fe302041a437bb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb63d61dfc56713e57e46a7824f04b93e66d1363f376760292431f221dba7969bb3cf2a8ed980f9aa2d1381c752b5d3bd4d10e6c0e6d555c369e81e04912ae8ae06dba857a1ad105bbc4945c64ee034dff8d8f034d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cb25eecbbbeb1f53284ff7a82cb5f7f6eb3c922f611f411e66cb35cd39c9e1251031b522a6fa18df35d4b7cdb5e5e6c4db2c8861baae893bd12c40f2758d1e1fa822d4856303b60e1b80492c17e1715e55f79d1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64d7aaae06cbc6afe6d3ee83434000e6aa73eed40ad87d8dfc58dbf4fbdb1162b0e578cff640e58b92f665db17a7a3b381612a3035162cfe8e452e0baf813249d8f309cdf71097380e7f1f9a46e558be8f71a9526;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b0462a3bb3df0d7b2eab9bc38dafbc23bb8aa9095cd6bc82823c1a9eb50fe8b43e41070058b86ee14fa9dd65dc1505d69c7df8f026a1982f40513dc83c02590e526250bf9f15a025ba4f2f4e59dda06fe3458eca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf18f75892a7403cb1956cccaa10890b6c32e20de1efb68cce2834778e03a9a57594099303b2062db0a0c8f80bf71b1c62ea9f76475401685c0cc300ef00a9f05007594fa2e4fbb04362ba0722194fa65257942b0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cf3657ae3828a8c0e291b3b57a082bfc2fca7582a23bc15ddf95ef450a0c6d94e74fd3712669d9d8d01adcd94099f3d905b9fe01ccf6d6d0b4d59bfb90ed20b36c16defe8840c60ebf7eebe5743f8c706958a11e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12e316afd3be1223a9f0b6c97804cadfaf27462a85df8c7faed4dc09ecb1251d5987596e7ed878b39a286e954e077e63780e910809b72525b17610f8ca23e72e7f9f37edd2af906a0f6aca718a4ea101581e77197;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7fe2153fffcff9acc48ca9e0416d885a83665103750e696a348540c1edc0a4993539be84b32af64649ae7fabf941fa94532a87b6df69b249b43e01a5d7b633f1bd0a6e9e3928ec52458f135a91805ee514396a08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59df1f186256c7854c4ce8cab566fdf4afc0d6ec70ecf38ce8eff2095a1e63df527e3dd564ce68b4a4b79110420e026cb6e467ecf60872f99baca9ca9ec2076bf31769522669bfaf148f1fb25918857799f396646;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h609720f909ad03e82058f47f24b0d4e80568b464209830688b9a72bb2fa951a983eea2e3861321c5604b7f661ef9c883ddd4a0c98fd7d309f1c977093b6a7a2ed569a4eaaff7c9cf0f01e61261d9781422a99efda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6e86bf2596a616e8ad6545c485ba2aae1e513817ef6a9c7bafccb597f89c99a121b22094cc1ed2742bc6d66ad74e64a1b39563670874bf2211f58815cb1d26ea86f08f52dcb8acce849c335a2f40a6cca8450116;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59464bdb8e48dbec9c25a22b988e921934cf8cfd3d0aa9ff4ad277e5643fdf0c5a3690c9d29c3531611397f8ba21ef87619804b1d4482177ff9de208aa2f5e0784980468e484ae03965ac22cff78fbaba522a5ac8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12e892bb22e436c5ee1ad9b23cbf9d217eedd92025b7676ffc4ce2272c1e3fe4eaa01473e85222132befe2c735da69430572e23504949ba1068c6c4c38d6144927e48399f253e1901eeed80634d3b96176342af1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h212191f43656f13cdcf36348b9f4ec70d8bb92b4fe913f96b33b91180df0102f45de1e324aa26043c32e8b6f6b5287de0864b2e6b28aa8f3faf37117f5eb01363d4976c3a9fc32a19e80660439a5bc1a12a3c22f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479896d7ddb9b867344d775dfabdc79ae40790b5aaf8667fea329c58bb83d6fa562644b63728fece0de26724115fd0eb8ce062675e40ef4c58a1e56a282c9b8f4ad43ca47bd279508eec3a9b00d9616259558914b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bdc5ae9d3c6c0aa232835496e9cc1e3f9ebe81005aa6ee402122dd32ec1c6b3bb571542ac9bc70c3b5213fafab43678205b173ab34d9a3f4f422f459840d1707161a186d287efe9366967a02b3071351828afca6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb230e0700c317ae41bf0cb20894136f40cdaac9831119b6059b475fe6755aee1197739144153ed3ab324823130a213ea5c62fe8bd41b9740629608ec90685707e778c46326e35eaf05e0668315d1162c25b15ae34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5347e7f46a6b0fd6364f3c4ea31cb6157763c21bd9c8e105d0f397bad190ca2487df1d51cbf434ca7b9577cbcf2138c8cbe5fd05091ccc6cabca96929d7673286eb48617e2112ee3c4b15b3431d8823c970ba6caf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a17044db43f37854e80fb1c330541dd93a3997abae67398c918ec92c035ebb493a43063d1523afdb51f8145fa156545b01757fbd465d08681a75169efbf13d77a49f523e8720ad8be8fa39349637eb6e708f5018;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b380e229bde8bd9359aa5171d45a5ac18f747bbd2ee0e4a369cedfa5b1ee730d997b3870b27a2d16d4eac21ce35505f90eed451f7e0ddf2fd27beb2bb0d1cae918002686b729d7cab69eb5244e64f9bf7d083766;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5afb8cf1d4220d83c8820b8aa3435646c6e80f4ef0617cc0df4d60a1d6a8da0e72bd37d25be3bf4f86b9d9e9644c21695647585d094c5be8a0b8855775b417f56753268e838fabed54f280c269e0681273d66812e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d2b772b082ab772acba72567b18d6a6c0d3216d6bbd934be1304bf603b8e3e64a770d04846e68c5b1be21faa425bcfeb7bba18b659dc81a476922bb9e777832701e604a15ac1e74c161f8ee768eaf3e8d653ab4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43178a5f2d17beed58e49b438cbb518b57990834374d670fd996dff84f185216b7a79371351c4ff616bfd78612eacddd5c4b25489107eba3d9034e1937ca573e389494139386771a7e247f160424f787ce2262812;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fec8041e18581faa9adb01412c2671d8ac5f6f8501afd8eda58306e794cc8e2844339a1d35fceef65efe1ea6ea9c8e91923c0a55d849067147630be6f993ad6ce6a035d804df62e70d775693d7afb1c2fda1333a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4635ca62ee08907f8e05c4f58874454808d9a0ab1709582ecb94ebbc8bcd7abb1aa46bb87dd387ecefd2a857a850b26f7222ca40d218a5865d23acd7fbee552d77903f050af0147ee921634c76cb54624fcaa878a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf9c3f272a3659df70eb1ebfc477d0697a92f7765bec31a7226c42b5885afaccbd87dd85d272b871f905261e292e52326d111e06587d1b642b0294004726814c69f71fac494fa43857ae9ebe80b4319a8321c4b69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2afed54e375b9b7a3f2c2495fd47ae888c02af72fca3dadf829cd6783225c48be8114af9958b8ee99055b3fcba0e733c740ee4fbfd6643b636b1741cb09f7d068e463acffdd51a17efffe448d505b98162325ff59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b3df16d110b200439f1f6d6985cbcfd8c596b29691a40a14145bf170891bfc7d815a8670fd6371f3f8f90050ad693f285e6396e50200675d23152f60fb444f06d8f6291246a34535332c00b2abc334322c24d799;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc45de771073f171235f701fc66a409a303c7b2837282f15d316eee7b34169ac977c4731d8081ee7a8ee4aa1395d1f273211474822b91616a06f3e3b1d84941e7432624a672c148d65e0609d8543e7c23c644a558;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a19746973b245312b416d3e55f3739efca8334f6e26c30ef2c182a3f7e915172d805014afb18a4910dafa4cdf3689a927830945a071fe5913449695ad4fbc9046a4f24707af8c778cdb66a84cf52aefc1903ef54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72319de8071240f2f7c9364a44a2f326c23dba0eacb30984a9f4d8857af30c2bd07e660c4bcf4e2ba0df9a41784fa9f8dfb41314e4493b7b9d3f8fe6006346ccfd3c6d31fbe20f72f484608da776e0a3d4b19163;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac38428c75cc0173b6f860fec5cea3135a732eae2c23b5372bcb8bca085853269cea4e1890c213ece1eb22b5ef34bfc357eb620bd72307b532f6f26793d1ebba9ad1d9f325fe7d525668b1c3b199ea220e714e0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a65b54e7bcec8e395e79c153ab1da44887c044d95b0168cdb1794c5b13879f0a873ac5d66d08367e64e8435fbb6058f209f91498c956888619ac722c323c686914b4d10d893d741160491da10f71dcfc7facc231;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8427e204dc1edb11b68c2507e782e1ab41fc961bc9905e6d4decde1f4993e4aeb424255a38f0c88ab38aa0328e08a4537563405e9d48965f55d08afaa892218c703f2d8e0523c14268fe059dbec0774b19ec0561;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48ab2c2b25b878fca89a6d0bee1458959ab0d584abb1b9035ff43f076134b09d1ca415fb7773bd443febd2004a92708af2d08cca6e9c995f8505ebe34536ec0ce50f8286b77693392c5d4da0b763cee7d36e0f05a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f95d2babbd13677199d48cdc009b2dc1764d2e3a9f32ec62944bb61cfc04e8aede70f1b1dc78f995fb6678cb141ec504d21107b864205268787faf98f41f3d4c1b3b124fe15ca366372fef194da8135b44ed9f8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cc767bae08caa793e5fced9bd5dc77911821c5b1e7ba5933ea16c298beb53a701d2bfcb09096ed0e3b9bff358f52cf74cebd20cb1359676542c2854ce4e6ac406cefa8a164b5e73aa0bd4eb96f76a85201fa4f24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h184725b79b716f40d12a7dcf97dbd11b3547af05e2cfab1b59fba9f9e53da9f85fd08c5feec4686152b91d436e79d9e3b9506a3b3eb8e0d73d0c8d8bcd3f22876b53cf72662217dccb11f6a479557be1f2c5fcacc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2e5ea3f6004247055dd1f9b9011baaa6746033732feff61090dfc72561e861f9ade6aaed190840711a0a0a1c42e71479d5d7a692f0218dfcbcc678d71fe4fdf02d2d1437b939186a2279e37c0b1c2c0f27b1e2ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h277b18fb4ae3a16ff1b3d1dafbb807157fdf1ae452922b0710f17d37fec5f16d26c2fedc44ac956415e1a73146ef7bf6aac0e6e356bcc7369ac09bb836f96ee11152d214f504ba0d088e9390616ca2de7aff1928b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7430c3928cec879f4f5bdc07cf7e95d45bf9a14a07ea7ccaffd51005105a39fe94362199b793af2af18828b4d8c4cff6b9467bdf2c09f6bd478d6c86e6b475635112d7c0e3ac0fd8a7f475464c8f39542cc7c2c21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57464db935b125d86e1c1ca156ac4116235bdeeb4bac1dac7c46eef48a0ed58f729979745c9709ec974a3d8e5a0352659fe6b67b36e9b9ea6d95a741d49e20cae5f9f9516a96e6208c3e6b8edc996231b774a4c57;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc295c0b3125dc16eebf00aaee12b32fc50b9520ccd8018ba5e3cc92ef3b9a749f3e1ec94b2b992726c5e588651a88f33cb61934c92ce5b845bbdb60f3d6f3e88b31606cb3a9cdcff7ab3c4cb7de3215a5c9186d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35479a9c1fd26d9d54bdadf5a045795cb5a5b9c370237e1107d3faf7da7b6965f05f55888deb1ae816fac93773328452e9f6f6d68192bc0d62063c269353cb08e8a1a08f47b3094d451a6587b92c655ad76b4aa03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64fd0268caacadfb88354c18a78b3445f26aa53d8e4a4302f5f14087289d0f12305350083a5e98c23886492a34a4dbe18f8dc485dc002e76bf3de64782e092db7972ce6b16af7141d8415081e464d6dd364f389a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb174e6969613c6d778051a6afc097515e682e26f355ffbc41926573b080fc0c30e48d2e1fcadbba0917454d584d8791f118699adc0fb516002fdd6945f7e420079871b8c4c380cecde67b21355fe3cc66551b5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14ae012ffb9aeab1402f46a08962e0bbd23b8d2e8b8bea9fd3ecab87c27f164fecebe81f01df8aeba8cfcbc51ad1234a309bc32fe18e6d132c142908cf2fdd8fc9ecbce5c2c26c7375b52fec9d4b098b73e1b5b05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5e9cc692265b7a24767ecc4f7b5c5bbf0b0e28e7124562d93242895d0b85c9c59fbbcb1604fddeb3e725daa7c1d2dab51cd4842f104c30cedd27089b54263c2a88697ca1e956e0c951b3f3fdf5c22da0475fef87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he69c71d27586ddd7f686a5a9cb72219be5fad526c18bd94334c19d4e1d45093149a812c9cc1b0a94eaafaa37fa6d7fb6e5dd008e9e1f042baa6de21ca8d5b80b3c52eb3cd63ef3dc9cf9789429f0d9bafa90564c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf012f3c37e84d6e672b91fdde6be612a4e44ed5a339bb12a492f1cba847be2c882c67ec285784fd3c5ef06a67ed59cefe5bb4410b40cae5757048ac92a0990d6bf7fa6bca9148b49f47d1c9314a255130170d5dbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddfafb9f20cb4b19c52219598d6c7ad246c5e69f42385114110e706ae32dc683e2cfd112d61d5eab04aec67ef1887f3ae2906d5297053d3869793f9cf1f717689886aa2c62a569a4e1ac74126067f7aacc78818ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h492847c15508ee34cfab5f7fa12d09b8f5b5b96406785e44742b98639755b3e66516517d0a237970aed3544af8bdf1aefdea16d9ffbe0fe45ff58677ede97608b217daef4e55ac1c7aaea26a68ce85ff1e1487186;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17134841cc5e12f2f1b20a7459ae8d88897f8e3356cad736f4d81684052abcecec24e8992af13915e2b7e216dedcb972ab9bfa152b535c6a6f09ec128f87f9374941147d1fc94573020e0287f94e72cbc32646f96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4b4fd823da997a94fa4b91bc9845364f6fa76803af9ee64b51597dadedc65b998a644f69932ee904358051d2b617c41538ecc8a7457cdbece909077071eacd8313473d775645cf69b586993df9dd33a0c9df80bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h219b04ffe6cbce9cf5c96328be714d1b0c2ff85ae8e9a9b23502099a90a1ba0e9b66a5565c542d264a9e7fed5a53a3a7a00c5123e9dadf05b36dce87cc6bcd690a9904ddb8346313d0b66e386ecb477584306341d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce0c5b146ca23407d7e4a51605fc9336624e1cef90cd45e6448218259df5ee51691ebe82483d5658b6a6ded2d750916d787d488e38724f7368a698fb86b83ed4a8d9a4323a78975852e8ff51f23006bf41c415e8f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d1820baf8feb86f6a1ecb4968d4d03c7f4188872b6b0d2728fde89c80cc0bba74d8f9160f4ad8bfdb29196fe0e110218e3eb85f005a08182fe304566fc7140f3ac73a2061bec7ebcb551875ad772f5d9650880de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he28092667997b26f9b86b642b5263291df836112fa245bba49ba6c647d3a2ac8982694f1091281ea1c5efe7b83971aa1cfe6ef15aed99f2e8a4ce42d22ae2e136f6665377ce4b336843f41be62c77f854e0459f5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800be4645a259d03d7fb0c2d901c9a13abc1e138bdde900deb681bc5ca119b977f3c98cdc2cf1fb3293337296d77a016877653f62b25aaebe7bf4d37fd9df2f97a62ce875cc30776b9b009acf267688404a49faec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0a05b87858c1df2deb3de422ccec19ebfa74b69b69177366af8e36f1ede87b6072a30050aadd6f3bb4ee2982aac9de784c859299f84bb1a42d8783fe1e8c6a95c99b3580cad14ec65f76d746bec1d4fc2533966d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fab53195a95eb1b4676d5410be0d99aabbdd75eb87ac18853d24fa7f3470fd6d05753b3603cd6434bea65c9a7db76409084ec894b760fe7d636fc31fddb9f01971e0155bd6daebc3289f0b8a68998483ae451c6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he55615268e0d4919d7c8ea8135483552811aef48aa07f5d5b6f4cde72ff53516909fbd3d8c3abae505b01c584bfe6f82388ee5a87ed6ed5aa88a369dd05f7047d8efbd1770e937574002b95c19d59cc915b6ce1e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23894da8c5b16eb9022a7e34080ea9f8f02a5817bce1407e37c01a362919e7bd7d28ec81c819e23fc30e27266d913e3fcc67d1fa41ec472ec3d7cecda5abe2677e0c01beeb5f059f5c282ce99a2bbdd3ac3be53b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8727436ccf1f0c0c693285c5b00c47f5ff2cd8be04097db422c02c241b9c5288a0e9a2907375c4523d8cb7d06ca8c03f0c3b0cc0b76a5ae9c9d71e9de7c40e0cc89875dd30bb3e54df70082b0884b707c82c547da;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79b7d8593dbd618df323100fd1b6c0abc1aa81f8de7d5e982bffaaecd625de54e14cba5091653660372fa81de6488ee5ef211935155b1c4babe862b83f593fea5bfccff41fcdd805b100ddaca813f56f00704e06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e1ede53a1fa524d1799d96cbfef59b26ef13d8b2df5d0317f9b8b86fa86ef305edba3a1f79b8ffb8da731e96de14da16dbc1cbe9fd0dfaf5b2c8ebfee3be215ca9d769d09d42a8cb16b19d636585db140effaf0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc71d54bb1190d654d1945e7a4ed4447d6ac9e6e57ca0e5af66e24074d1e29e35f2148d97ffb0f3d07bf435f6c58eca72cb23a0a31dd0648f7d7a8b09125cd362b61ecde714817b4b3108137b1fb9d68eafead3a84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h256e87101a2fe72f74215cebeac5e116d3ccea9064013af3381f73b54c180438db18af65da84caeb0019f9d1f3a9675d52f2804d0cd74fc739db6689cc636a2ac0b064d839cf4242b6dd4b5ffe848e58de2b18bf1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1593c5f8765758d1f1ec3743dd8d70d27cb8cace9ae7a9f2c353227f4989896cecd9aa1652e43858fb47abb67d39e25bd84850eafe7f0f09f1444e79916e6f0c62e02f3881d4af9b4b18b85c2829d22132f378e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd24ce7c4429b0f8b22e98c0061600bbd1af28d39ae64cd58170caaf3bca966bf8c5206ee74304874f51c50c190871488d4c10adebb4a068921febb2f0a47f46d915a2648b2ce6720837d606789fb819bb5c95e281;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29a7e825d05ccd144171d4e170486040928c642b17f00a6fcce116121389865b41ccf5f72effeddb0ad656ad014b35e259f914ce32fb70db33eb18e98936f95a8f801b90263c15eec1d241498fbe4bb66cbae898a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b611fe9ba546b364c9162dcfca1ad63ca5e922fdab72287f65e8484b223ae1bea5e68716d5b6115bf48af244aa6199078d04d7b0a0303bf566665691f9acafc486c18418e81a8cd18d8565e38b0a06c4377dba0e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ea9897423cbaabb948a2865d50b4e02e47912f90bda0a1c2704b3200790bb1805bf50936d70c2d52af0af21fd3ddad4318a48d2a2ebb819aa3ba55932d1bac285aca1753ece7b668bc05944534b623b31f3e23f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22d642b9b736460e9e6a7bfb66f6652abf2059fc056244cecfa901c981ac10b5fe6fdf6d31f2090ab0c89637f53bfe0d6a63e1ebcdc773a455000e5a8570789f42f760a559a3f338205ad1c51152c4ac09b975bb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc40791f74e662e10a163fc348e98decbd5067e86c6b5fabfbae500708b7636f439cf447e836745eb0139949fbffe262dfdab8d13f9a8463e4d778ee4582305332583d835fec5ee65c77224c758010d5406ee345;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h703a1a87166cff460a0437c58b381efdd08558261a0d1ef4e95cd1fdbe07099d0eff9fa6a3309421b4ed0c83cf42e8742e2e3aa4b6fb649998657c2593078ad49ab9a0330c2209c6fdab6b33be920957c20be99f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he116ae84085f29861232f555733acff99224fc2b2da53d303c1d4f5afb88ab694ac6f7550cddf56f9d7b857f207e2e9e0b1f148614a35539d7d31544cc622d84640a96382dafd3ead31cb48cc2aa6611ee04b045a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he875dfbd35e8a6225331ec2044a77db0dd0777ec1a128dda83643e181494598b8fb3af8dba35c5ed072d2bc206cf8e975b550a56eccc63661b0f6c33736cac242619eb71ac4f4ddb5b946c8c847084e965beb9be3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b888d359fe568a15f785f976498de0137fcb2f7e4fc57419a314b4b5520ee9256852ab2761faa2b029980503a7c78b8c480cb7076b3a06160742365029811d04072281887e131635a5ad01c851a92256a171beb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3c8b9577164c35c6d9e70fdbc6fd4a188434699e32318b8ae7ca3b42c4981f106674011fb2508be967e909401452ff78a10ef63b3fd26597a36c9d1a146d44b12cdf044778f53fd7877db98f743fe5e90321b8d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bc83f693bcd01fc5f999de4373553384f08bbabd76d75371a760d8286d7c763bb447a0215d55e884ab6cc307863afe123eaaa78f68dd8770910475fb78a5fcc4a86eacea1cecfdc99ac54daa89261777157ec1e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h828ef3b504896f3146cb364115eebac01f9fdb0cc8e2205cf230926f0488ad4a6fd139ae264ad6f03406c3ef77a73e5be73b1a300e427ea150f5463bca1f6868ebdecec1c0883114aa839747f69a08c671d52b8fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7783627c1bea5967b1766c7857b4e2af94e1f06bf3094640ce5120dfc30e90f723c22a920cb8c64addbc14ef05af985d79fe2ac7c1d3322289f12228135e019a6662563a658e90f3c8c3af5ea262a6580a7043cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1eeed68a5ae3942f96ae381ff74c8980d2ad76cf89948b8e4ddb94fa7067d2b1facd5ac89f8de5148602d33fce43c05b6514a2d38f26615110d1ea14252a12250372544d364073c6e1b7dca2e4f9ca77e29dbe69b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd761f2fbe93d7b04703fb13b8d7f5d1c42d0ea60299fd3bb14f0ce87d558d450e96409879f52baafe867b3e886abea253f8d0dfd3295068f0d164830ea5898e817425ad1780660512d1d96f4c007536621627a98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he61ce62ac3405995687b35c1a300dad8b5dc457d019b7106e4bbf25b792828900b292d653dbfe3f1dd3fa563f0bdbc75e910ddc7acb8a747e8d9517cffcfa99a13f847df5a3eda34c40648360509ccb056942b42d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ab893351235e13c7b9dabe662dba75a53197f45273e50105b5922cd4f4cb98c6ccc27e998ae7811a9b9a0b03b13e656a3ed32bf7e0574dd6ff2473ea3cd4f9743a4069eaadea696c3ef0af65aed3fa58be550e84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb933dcbe385a77582dcfc79af80ae5935af88ec89291ea4f4c4bca05393a9849795d6282becc25ba88225ed2a47bc696ae0d7c5eb350b0e008f8cb8ed7f250e433f3adce7e78a75590186c3e39f50ddced93345f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10e3fb2566e2604b68fb66a24e68d829f2e376d09e0999d99a29d66bd2c7574dac23f3f5de81d252c85c4cfda30b1c37410f6a02bda62870224137f1a8137909dd391c342634836625c6e73e36d8e24377d89ef51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9490d67eb28f560cb696193dd816edf2d711d934f67e07b8e963c8c8d2fd364498516a3acf3530624ec424d9487754e0a2238b1e01c22d9b7c3a904fc216f1bff2c27d3128ab35df00386afaaa70b88aa86bb3977;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaa4f36d61b33ceb3494a74b916cfbacdb1775a2e1ff206a9885b2318d422be932844a37e576350f5417d8cd36ba60c590cfc358a37326a8b7b36785bc82d78e9efedda92c4b1833264dbb1179f2e390ad7db22b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2912763588bc253d44900a3f58ac3ead8ff4acd856fa8d4cb519e58184c27dc2eb0f4b3bbd6fdafa97164d096e57a6406fb32ed35251343abe8c1d052ea37e8334d1be962966ca50120c08e1cbc054f09e21aa2dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbfd763776b19b6e6bbda51cde67d30ca918a6bf3546cba6c1eabfe2dd24ff6e8f3a41c7a25faaef8fff1354eeb5c583d3cb588a94fe65883fc2cade61fc54e4272152ed0b128449bff8070cf90ccb7771de820c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79400ef2834ca4d7caa37b955cdaae4ff640769fc67d7656ae90fd42eee2b91e781675f85bab958c390b26fb2eb6bf90e9c4010d102b8dbe3b635902e15497c00bc5fa78faeb84898bdaffef594d87d16a61bd3c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55ff9addf41d6e0b1c153dc2b92fb13e0b14d44bb9f30ceba73b9d7e628d6f41b116c8e45f9f2dd2a9d7fe8d78873ee003071f28ac44bcb0cc3cac00724f0d9e5245e8f6bbb52edb33f32814e190b5c41ebb9fdb3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16d4ae62dd920874ce9c3eecf0a193d2c76469bdc2919cf7b0a17e2b513829a52fecca81f1690b9abc63ab7a5bac4d2aa940a3acf460723aa1c02a61129f5814c1f24835c7087eea51b1a9311a7e63dc09f914b01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca8050c30236344242a324a3e67448bdbf0452fb563361bc66f7908788228ea9d8313f08120a9a0f663228e78a7d7318a7991901a9bf90822f2d87ada79282232078e4e05b4173083ebbc6b2f8d9771616cb1a09c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5d5b74bb14e81e9b32ccbeb922baa754842e6ef1f212eb716280b6246dae5e533f7b34b643f397f509437658519a890da0c5d2a2d4698d90886abaec57ad5761d0d4322ea78f8b462b4f0dbafc0320f3c404ed50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h588b371f5f3ddfeff409b3ce47b97a2a752414df3c8e7724c1b91aa587018c76c4809f3479e4533ac66f365902a20454767cea6b7e7d54e195398702c2aa4490494af16808344adea59507b6d0adb16eeedef1496;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf165416e0e6099971977d32adc1173ea2a039f04a5d95f275a9410d5f392013895ac291902468c92da98343b478cece44101e04a159f29fa819e9423c9f40b4027c634bfee4eda648d31f2bb0f0c6480b764221f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd07a5587b4bbd4abb047ddb18c6613027858f16fb0e066acced62eb4563f56ce6d2283c49f7dfb7fedf13a81c4c1819d7aa57794c3df737ca64bcbc4da5735fc4b36815605d440efe0b0c05f571597cce5765f6ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1160b3146a76c19ab5714bbb39175886f6cc9ff0c696efce283fb4f09eaad9bdb43d9b1a2fcc3e02cad4cc4fec14e60c6e5e5336b20159e2cc5589cbacca5a4aa441be5771cf17463341594bb33d28e3619b9a34b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2430e96862b379d35ffe67756de76a2e562148b5d587b398bafd27f803d9c95de4748b1852becbafec68ee3111bbc49a6bca40eb472bf14f8c033731ab64afa39d7a507dd0355ca03ca72443dc62c85cb77137fa2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1657ae15996284b35528af68c37f85872f57d7c5db8c8ce0fc242c94c6a8c181c9019f4eea5175ff3af98dd41b77c2f861152c7c03d920e55ffa05f8eedd2fce740fe4916676596eb7ca4679908a519e4789fb43e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5f7cb8463329e5ff2565eb2daef945848f89a82090be826688ec209ba57085ff449b91f42d0ccdbf8d354e78e509077502776771553a30d40160c7bde216790b07ffda77450a640486c8d4eae9f155fd5b741e49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf70ac351e50c5e4733cebd9e85d1ba5c61c4655a0bf0a6c9bd1fe43c1b2a27c48bf57003fb411004616e3d91ddf5f12d56b3b94b7ba0b1e84ad6d24a7af6e4e6b0e4067ba5ca448cac206499988a7cc7533a05257;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf42ef2579b80608da45f5d4a1a51994a88d54d86751df9d766d4e036c5975054d7e615f980fd92e859ee3ce22b395bbbf3fa2a0b1c031871ae4447dc335e52967ac0fa3904bca167cffd15e8dcd3543e0fcb8ca90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1aaa1ca15a34d8d717a7c6f0f8faad80162917cfdda04937b694ae914e92ba86c1c6fe2466834cd36a4bcd504b8c288b1a48c315dd7337cd4083414c24b4c6a0257d32e2048a9c97b9a29762e6e61a53c4dbb6c3e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3134b15c528e671242d07c88e25e0cb8cf3d8090f6327d530b24ae15f1d7e6bf3f8a6af94d41ce13cbd4fc9fac3736ea1d294ae9483ff5fee55141d962f68109ff1e0bb75497c0eab833759c3c2b06352623d70a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22c19d0def1496433d2d0f420b2590e80a4e316b29c7e0c18cb5f5427088f31e7e75c914216b8edc240eec0db2bbc3e86303acd93bfa475cc8892334c8747a400fbc5225953e5b9897f048bb0d093676416047dfd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf196b67c11b33e965455ea82ad5da00594818d6f3ce8e00908d3031d8b8074bc4aa6e3fed8bbb0f414388b1359c2182568095c7f3b8a5fd081cdc61111ae0500f6a900579366b63a577e2f95ed90008f527960af1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37f590148f3398970b2ea510f8f01e17d75474393c438a8f9b9965160b014c0759a56d5459bed0e1ea3943fdb337cfd243f58c09393c93539259021d12415b4dfe59128a00e9843cb67e076e34d99f822b712a76d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he571b51334ded58ddcbd70e07361bff8e5ca944b8a427e1becd55ba1529ee2c23e1722e8426ed4b41c7c0c739b1b7acf374ec7ebedcbc9ad0c06acb6e540f272e133498a0009364a63145f7dcfbe2e1a97214ec5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31769a526a8a00562ca660c5e1962409db6d18fa27bbe0245296140fadbca7f63b6f325d3d877c61c4ed4dff2d5e07c1bb07b25cc42aee46961ee33816ea1d3fc93fae545bfc0d617ef73a2571c7d8df46c06862b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30408fb5718d5024d6eba096fb40f63da2f00bea1d9a4a26a9a90d534e65d35562ded1b2a5594c774668f1bfdbaef5ecfb1c2f1383e256343a1ec3dac00d5fb3b430a3a79e4c79723b1993ccd73e2c4b6925042ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f9b96606403a00a79c8fbdd8fc51701631bd2f35dd8bfd1c2751bcaf09e005d415c6e019f292fcd8ad9e341dc9fb060e4d415aecc79e86b05b24841c388aec6a9375740e777f6e5a05493425c9fac7c1b7b7a3ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed021f85a8377b762697d1a5aabbb7e655499e31bd0542dab99bd7f60fb9f3197f74deef573c30be8ffbd0815443b55be7356e780398456b83eb7bc162772baa405bbb5ea548982609c166f1e685fb87bb1142bab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdff95b5c7ed6b4041a03a514b1cab24a867cced8a37e381ab4245095b21862e2ace4b78e99b87c7362e161174c656bd17ed8450fe822057b71f1989b01c45005a6023a621e8a874232f9fb542f3d3dab03a6561ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b89dd9a400adfe42ec45392c23119a8136deec38fcde80f25721b38d33671e4a9b212292a96bbd5d851184abf4da236009c6c825d7703fcadc3ea032198b414896dff8f191d8369975f533f6b696db30d925609e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9531cb1c7c0bd9e74c8c61a68e9178535d0478871ce395fa74f1264374f150dc4c6ea71fdfc02219975f1cba2d79c7cabd3a220d136f2841037662dabcd995ecf9606e6746a217befc0850720d9095efad4319be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a5a6bdd27af81bcb3db1da1c630bccd55fca366c6203914e0d358e8e529f473d36dc2a6e73741981ed392aea70f4b5c83bb14d17f7f986570005ae96f9d8470369b385ddb7cd8bf51cb7f2888ecb99672781cb99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f56991b168c66c9ee051fcfa2c09d50a43c9bcbc3dc1599a336a63965d9a54ee1bcfb108a5b002201f0ac6ca323eb7cc97bfae949407c4a59b45abc959727570f203139e5ef211674a1682383f1a1cd215c58b69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb155a8dfe0c44d2e2261fcd21073bfa0932e8a7ee28891129eab45b337603cac4a4792f741a58e6564188e7a0eb72bd204f4c59948f3ef945e049197d6c340522d6d301f9c89bf6f37a47231a5cbb4aceafabb2f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4ee7111b1a93851fb5e6ae01786120b4c247ff9e6394c9288bef0aa1814d7c012f1bb453437471e61df3535af8fcea93ed8dd71df1fe28a033ffb642816b47f75db39d4b0a147f64325f9c0ac047a0e47dbec6ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2581d14ec4de22c861d957f21c2e0b22ea61fcad57dbaf2b313be760afa4b66db9dc27f3252f866ea66bd527cc4405fbb8098f4320c9e13752ff587e609fb7c8f83b37b6e83d2e7f6c85503968d63f9564bc43b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc93c824ecfe2ed363a1e94ad0c3a72eb574ea017794e26ad239f5d520bcf7d1bc02e291e77dd85d8b45b766b7b3fd0d0433fc34806809e1302f8970e630fb0a1766b0a8a9be587465fd7e8d908ce5a9ba193b192;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78da70e367384aa75b92488164c3ee594f21e5cdc683ac0524fdfa93d86bfe5b008536f94c7747414b34ad823cb7f150adc3ca28577c9e99bbd7f8512d36d870ffd29cae30db770f2ed2683dcca4f8e06f590e0a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c56557f72ebe8ea3a67cea07605e258a4f48d35dc9ecba61269b2be6aea8ce771fde4de471627e2d787cffc70ab7feea7b8fe98e601d7e1675fbda060e1cec0241664f7234c83addc3f1f69c92a347154f57c69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8a15bd007563963056da9da21930814c9de8db68c2e29830f4e9cfd606fc430226d0d6717dc9383bf0947dbb1fb1d41a235850fc6e9bb1ee3059db666c23146a35a7f7e9bf7d32f8a3743a1238a55baba51109b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d8e722d64bf258599294df5906ebd9d9de39a5a6e74dc51e6844de53845d2bc10037224256bbadca51c546eee7a041702b99b11d4069600506fd421ebdc86ee7224bec51c789fbaf469e28c4fc5b929ad3e444c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebcce117cbc2963c029a5092fd27c30dacb5f44f2e34515533e5a32e73c193c8720bbc5a07dc840ad12f5e656e8ee36357993bd3596a4e4a06f80bab99bc46c393062c4d69a1bbcde914f7c9a0b603a6e32a162ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h320fb40a2bfee1d010297e5110864d8e7cb5958b6acc1cd1c608aacb870dd49c4ff9e3e1500b61787964cd802aeb89bdb067828ac5cd5fd0db790a1546b400c662e6f14500f0610fd09978c048707a3fe4ad6ff45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6612f1e9e7c14705bdbe202d1c488b0cceb3aba9bb348e8cd037dee3616aa3c83645024b9b69c1e7cea1d397731fd45327173a6c35e3079fe06f90991e245b561eb030c657b97e739847bf2dd2e669c5a5fceb9bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b08c6c33581c26eca5a49031bf3a6b01aafd94b9be4c855df4e88a919b35665d570d90f5ad5c5e0bbc0205a15de884b43ce321e714cf6b9f01206c50b173fa1f50bdfeacad140ef4a390c242eb661314c3104a05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he42991479dadcc66ee12c36b823c69664e9daf10c7c0ca6a2d65a57e8b54ba1f55a1de08e32306f02a0ac5ad29b4a76efbee16029a82126590892fbf4b1a901d31ef5d2d4451099e1aabdea886bd2164240a64567;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7923a006ac53a29dd4b9bbc466950abfe226145788c396c03e2d3af726226b94e7f853dfe95cf4d02834dfc7384657c32e9d9ba75b78b4e119fb15547615037a16ae7aee3ca1716a5e17385de6f2a14961206438;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadb2508e78c328dfcaeb5779b93a4b8b5a7dd62ee54d625c46876c4ef27358e7e40a6781a43fdff3cb197baee85e7922d7b46a8ed5795c67b663c630fd95e76c64b403ae31bd42979c02db7459a5f930fbe5a3690;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d69df08ad3c7f54b97dedf03e5cf1fe9b58092e65eb111bbd266768651fcbad429beb3c248c12daa7845830d22945337c8af3df67d4b7e055c789971f5b0d0febf187f6d65aa4112765477991777a215ee145d49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24f184d8cbe97a01cb8e9be6dd4eff8155794b3937337439e6603943c7bea828989e5086bd59a2f722a9a1f117e1a2f16128fcd195d865a66e92c38031b64d3c314001cb9fe4aa59946630fa89ec94b05383f51e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e39619c8a58d862bcbb483d1902f1360ed887b9585d766d7cfcec815e22337658139390d12c364c4058fff7527b969bfaa8c754a2fbdad92140c04cb07ca7f0f4d7adb96ade8f6ccdac4c93d85b00d6f286015d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b0f31a396ffea30aad1408ab9abf8a7ec3665e1a699b945dea747b09c9e722de82e02bd66605678ea9c855fd7c74013f6e25c1cfb1ccd0f37d16f1e80e728d394e11c4b1cec5511ec3934e6619727ffd79c4274a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e5cfc533f1eaf203e5077cdee0c1b62253913285118c877aff467694419290fc23358184b0e640241aa75902bfee38498702d03101dbbbfe49832e1c3231b14e593507e4097512343b1fe938c181fbb0081a56e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36fe78ef70226017091f7fb2079aa8d56a99f5bfcfb0820fddd04328f03545d8d12a45dc0786e2ce9c0f457e7c27d0147b70d4946d54c9d2e67b890adaa77e492858dfcfc7d3ca2905d2195fac632faea877e1bb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fcd18319aaaa908ee9d4a2020fe32d95dc197f77ac7edbce0187a342abe395b8ff1b7ebe2e94e99a0f84a796a6dfcff83cd773f7fad7479f7d5b47c44c1c80204b9f37b94acfde59f708c02cede35b839711e183;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c16e10eda4b4405846f2f6248706bbaa84d8dc1aa906dcadd1e045a85cde454efbdbbb34f9256da787a04c6c22f0ace8cc8d4f5cd5e0cef97862b7d2094f7de6a00abcb8030ffb123538e70a9d915c5b87b7013c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd07d3ebbfce57cf2798c23050a80624a0a409f1af1ac30ce7078192c67d59913d3edc0af3a59b69f8828bd599de47e2f82e51286de608be67ed61f13dd875e8547e76b02e3f98b7f0122d7b62a2ee77bec013e3ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf42cb1f7e465d81990438c8e9d7bee23219f1163bd5026ab982effc9bedf6c2ba434254d9b14ca097881eab90b3e6680638ff6762dd7789a14a43a676d49930df552cd2c5e5e819b1b87695428b90c32a04a7dfdd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e3beebaac3fe5798367dc2c35346bdef883886ee9dcf94a49d3dd85545d8f8b3dfee38b7aa4492d8e4fa952f9af160a51ad084368ee361857cf641add4452906eadbcd77db2a6e97fd771f990559bce11837eb0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf656bc5fa0f8509ada25471e27c8e42eb805a8f2678bfcaddd25d9d15e259116180442088735aa94ad6a03864837586ba5b354179e1fe4cbe63686b18f97fd0196987fec0398a6a4605455d0687330100a4008f18;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50c4aa5409289a07483c582318113225d42ca1d041f90695e831f5b50869b3efe450f06f3cdd0d46fb53ce8f18a47adc824bb4b04491b1b9ddfe7e9df39db95d6adda195b603c68308f30e87dc07f6e65cf8ab14b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29536076d56917d005cbd6abd98aba98f858fbfcf545140f16d57f15d15d6751fffd2973a783af404599cdfdc06e7ecd0537e86e34897f68247d4b227518d80124b5cdce1a4a1ab72f1f426b5baddcfb3c2e8b1e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h720ffd2948322ccadba495049fdec62860c05d40c5f1e006d108658e3389eeba29e7683084c311a0c1a9666b5da1c8f501ad250df0e46eda53ddf062ca4221f445fd7436c605dbc8bf702cf1f2af5eb36fdea30e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cd75859297c92d6ffa4bf7ea4f0dc21329af39442bca3d9ecfe9e8cccea6bf5221d08ecc2ffd74bebe90bf609194c686e80a59007d1acad9a3c475dc58d49c07aaa3aa111bf00da1275d7ade972bbc8ac9f05ddd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fcb74d8e73ccd5dcf1a6243a06c33c1a88e4e0331cbd319a850f449c88377daeca82f90f7e8332e035dc3082f43c6539b5154ad511959abc432a9bdca808d58b385fcfe863348f43cb4567a994ffb5f5346a3666;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2404d89c57bb792815722bfa0a8eb9ae162d8bba4bc3ce7d8c72edb4c120536a1a8bb908d72a6ab649b17d3609928dc3a368cd3906422bddd8986c16b023f777857b0672907caaa620a7a7b69832d20775391c4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6383126f02fed3d4971d99dd6fd7ae5a734172334abc088821e1306d1eab28155ebbc55c6c906b229e55de217f6c3680675e0842d963c6d2d205ddf79486a16cb2e8293797cf23812ae6739f33c0993e64a4cef2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb73d48d96ce70196165eeaa3b367b2a03b2571c3607709de197ddf7865a84b94ad9d4d8cb01a51a47d27e1f2c6c49a124e5222cfd69730d44ee00fdcfc46ca0f118d784e8952329244b5b1fa234e57e78d529c58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2756c7cbbc1a7e3986c3928510ca7b9eb5df90fbaddd245826a9b595446800cb332c9787eda1b9f106276f4a6a675c0dcb0ba6b536d30fe789109a5320f47f60405106345a4a19446249d4d689e28edf4c3f8a509;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf6ab7e789b1cad3896e4e3fb5f40583b049518eaf2bf2f8ac48cac0d6be5938813100ab92fc899be66038ecf9aa4dd25a099bac731ebb781bf79afce410941789dacfe688bb616e929540e30668fd6b1cc0ca654;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c5007f41fea282467b08e39587e69ae1b60b48d32407f84555f90804bd68969921430d937733edee5f774c88b7fc7f46462c31aeb9edfd03ff9803d52e9d5df2dc7af292e0d43a50c0835ae1bc0000fcad784007;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54eefc77047f73a3e2d97364aa478c1f8b6e959220a23afb22045e8b63cae8c2dab1d58ea477860da0530928a8d389b9a80a7ea53168dd240b9a069cb9145d6639e6b579204aac7f64bc49752c48c06f1f56b4722;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcea117484fd4eb126f59607672e88ee1adace698fa8fc195fb4272942f87d944d8fa493f0f2afcc66866cf1aec87f66ae75203cb5c55ad71f615b0898fc3572055d1c887a9417cb259f4df93ecb515e4f8febd881;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb08e8e4bee22a3b3d7aa85162493e9c1dada7e8c1177e07d902bb0f4d53d9b4e12eca695c89b3ddf157932884de9400211b7fe73efd88bfb5920380a8936bd3bb6472068e148f9f89eca98ed5bf9077bbcec6d4c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99679c44577daf7f7dac9cd49f4f4db7b7531928b0d1b204474caf51616fac2b6898a4ad72f68dc6446b5a5da6c3710270865bc0d82c75cea85bf327fc2b269cb2a8beae12ef3c933832e54748ca6749c5b028fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a117ee2e43bdde8a6e3095baea1f7d99a20fe9a42f32afe4d604890ffe68c075f7f5ed5b8f9677d7da1c005e8c8f5bf22187d28af14c57b339ac94aaf7554b2e03e5b0940f0f0b22a7a865af67f47232da6d8a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10d37df08539ffadd190f67c96f52b3793965e9c4791ae182791103db56ed067c0fa65b55c97cae8134677df3f40c457ba99f0cb449c7b17715e10d88e1f7fef11bbd043ca13cf70151b9fea9d54ddbab947d62b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab14fa18d36d4ad3855f4349d4e4d9660c640a035f36865e94f74932dd6263d4264cc7c45313ea9027cfb1fc37b71e650c30c747cf65d535168d68fdec10df96bd045848eeda84df69cbe923d46c7a83f72f98b03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcee2d3b74a6710bbcfcf2b9421c4555d11b8bb349d5bd4bc33b44a6a5681eb893cc994da9d68b55ca109cedea5f802727870f691816b0345ec469647c4a684ddf455b0b6d86db00e837d0eaa90ae625fed08b8b93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8aa349dabccef0469bab7c9c29933a70ff3f608e1c1a1b9d89f19f1da9498ff866f7d3d13950ed099f210fe779892b034d1e9a83bdb3514808da229efd4799c38517d9295a6feea6649d15e4acdaa9f6dcd3b35fc;
        #1
        $finish();
    end
endmodule
