module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    compressor2_1_128_16 compressor2_1_128_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_128_16(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    rowadder2_1_23 rowadder2_1inst(
        .src0({comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [45:0] stage1_0;
   wire [63:0] stage1_1;
   wire [38:0] stage1_2;
   wire [48:0] stage1_3;
   wire [59:0] stage1_4;
   wire [56:0] stage1_5;
   wire [47:0] stage1_6;
   wire [64:0] stage1_7;
   wire [55:0] stage1_8;
   wire [57:0] stage1_9;
   wire [53:0] stage1_10;
   wire [51:0] stage1_11;
   wire [56:0] stage1_12;
   wire [71:0] stage1_13;
   wire [70:0] stage1_14;
   wire [37:0] stage1_15;
   wire [35:0] stage1_16;
   wire [20:0] stage1_17;
   wire [14:0] stage2_0;
   wire [13:0] stage2_1;
   wire [19:0] stage2_2;
   wire [19:0] stage2_3;
   wire [27:0] stage2_4;
   wire [27:0] stage2_5;
   wire [16:0] stage2_6;
   wire [30:0] stage2_7;
   wire [28:0] stage2_8;
   wire [20:0] stage2_9;
   wire [17:0] stage2_10;
   wire [37:0] stage2_11;
   wire [28:0] stage2_12;
   wire [18:0] stage2_13;
   wire [34:0] stage2_14;
   wire [26:0] stage2_15;
   wire [19:0] stage2_16;
   wire [19:0] stage2_17;
   wire [6:0] stage2_18;
   wire [1:0] stage2_19;
   wire [14:0] stage3_0;
   wire [8:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [8:0] stage3_4;
   wire [9:0] stage3_5;
   wire [10:0] stage3_6;
   wire [8:0] stage3_7;
   wire [13:0] stage3_8;
   wire [12:0] stage3_9;
   wire [7:0] stage3_10;
   wire [16:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [15:0] stage3_14;
   wire [10:0] stage3_15;
   wire [19:0] stage3_16;
   wire [6:0] stage3_17;
   wire [5:0] stage3_18;
   wire [5:0] stage3_19;
   wire [0:0] stage3_20;
   wire [5:0] stage4_0;
   wire [9:0] stage4_1;
   wire [2:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [4:0] stage4_5;
   wire [3:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [5:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [5:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [2:0] stage5_2;
   wire [6:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [0:0] stage5_6;
   wire [4:0] stage5_7;
   wire [1:0] stage5_8;
   wire [6:0] stage5_9;
   wire [0:0] stage5_10;
   wire [4:0] stage5_11;
   wire [1:0] stage5_12;
   wire [6:0] stage5_13;
   wire [0:0] stage5_14;
   wire [4:0] stage5_15;
   wire [5:0] stage5_16;
   wire [5:0] stage5_17;
   wire [2:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [0:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc606_5 gpc18 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc606_5 gpc19 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc606_5 gpc20 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20]}
   );
   gpc606_5 gpc21 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage1_5[4],stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21]}
   );
   gpc606_5 gpc22 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[5],stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[6],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[7],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[8],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[9],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[10],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[11],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[12],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[13],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[14],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[15],stage1_4[32],stage1_3[32],stage1_2[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[16],stage1_4[33],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[17],stage1_4[34],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[18],stage1_4[35],stage1_3[35],stage1_2[35]}
   );
   gpc615_5 gpc36 (
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage0_3[91]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[19],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc615_5 gpc37 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[30]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[5],stage1_5[20],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[31]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[6],stage1_5[21],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[32]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[7],stage1_5[22],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[33]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[8],stage1_5[23],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[34]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[9],stage1_5[24],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage0_4[35]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[10],stage1_5[25],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[6],stage1_6[11],stage1_5[26],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[7],stage1_6[12],stage1_5[27],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[8],stage1_6[13],stage1_5[28],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[9],stage1_6[14],stage1_5[29],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[10],stage1_6[15],stage1_5[30],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[11],stage1_6[16],stage1_5[31],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[12],stage1_6[17],stage1_5[32],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[13],stage1_6[18],stage1_5[33],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[14],stage1_6[19],stage1_5[34],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[15],stage1_6[20],stage1_5[35],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[16],stage1_6[21],stage1_5[36],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[17],stage1_6[22],stage1_5[37],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[18],stage1_6[23],stage1_5[38],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[19],stage1_6[24],stage1_5[39],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[20],stage1_6[25],stage1_5[40],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[21],stage1_6[26],stage1_5[41]}
   );
   gpc606_5 gpc59 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[22],stage1_6[27],stage1_5[42]}
   );
   gpc606_5 gpc60 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[23],stage1_6[28],stage1_5[43]}
   );
   gpc606_5 gpc61 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[24],stage1_6[29],stage1_5[44]}
   );
   gpc606_5 gpc62 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[25],stage1_6[30],stage1_5[45]}
   );
   gpc606_5 gpc63 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[26],stage1_6[31],stage1_5[46]}
   );
   gpc606_5 gpc64 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[27],stage1_6[32],stage1_5[47]}
   );
   gpc606_5 gpc65 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[28],stage1_6[33],stage1_5[48]}
   );
   gpc606_5 gpc66 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[29],stage1_6[34],stage1_5[49]}
   );
   gpc606_5 gpc67 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[30],stage1_6[35],stage1_5[50]}
   );
   gpc606_5 gpc68 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[31],stage1_6[36],stage1_5[51]}
   );
   gpc606_5 gpc69 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[32],stage1_6[37],stage1_5[52]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[90]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[33],stage1_6[38],stage1_5[53]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[91]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[34],stage1_6[39],stage1_5[54]}
   );
   gpc615_5 gpc72 (
      {stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_6[92]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[35],stage1_6[40],stage1_5[55]}
   );
   gpc615_5 gpc73 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_6[93]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[36],stage1_6[41],stage1_5[56]}
   );
   gpc606_5 gpc74 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[16],stage1_8[31],stage1_7[37],stage1_6[42]}
   );
   gpc606_5 gpc75 (
      {stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[17],stage1_8[32],stage1_7[38],stage1_6[43]}
   );
   gpc606_5 gpc76 (
      {stage0_6[106], stage0_6[107], stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[18],stage1_8[33],stage1_7[39],stage1_6[44]}
   );
   gpc606_5 gpc77 (
      {stage0_6[112], stage0_6[113], stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[19],stage1_8[34],stage1_7[40],stage1_6[45]}
   );
   gpc615_5 gpc78 (
      {stage0_6[118], stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122]},
      {stage0_7[96]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[20],stage1_8[35],stage1_7[41],stage1_6[46]}
   );
   gpc615_5 gpc79 (
      {stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127]},
      {stage0_7[97]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[21],stage1_8[36],stage1_7[42],stage1_6[47]}
   );
   gpc615_5 gpc80 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[36]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[6],stage1_9[22],stage1_8[37],stage1_7[43]}
   );
   gpc615_5 gpc81 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[7],stage1_9[23],stage1_8[38],stage1_7[44]}
   );
   gpc606_5 gpc82 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[8],stage1_9[24],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[9],stage1_9[25],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[10],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[11],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[12],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[13],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[14],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[15],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[16],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[17],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[18],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[19],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[20],stage1_9[36],stage1_8[51]}
   );
   gpc615_5 gpc95 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_9[12]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[21],stage1_9[37],stage1_8[52]}
   );
   gpc615_5 gpc96 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_9[13]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[22],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc97 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[15],stage1_11[17],stage1_10[23],stage1_9[39]}
   );
   gpc606_5 gpc98 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[16],stage1_11[18],stage1_10[24],stage1_9[40]}
   );
   gpc606_5 gpc99 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[17],stage1_11[19],stage1_10[25],stage1_9[41]}
   );
   gpc606_5 gpc100 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[18],stage1_11[20],stage1_10[26],stage1_9[42]}
   );
   gpc606_5 gpc101 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[19],stage1_11[21],stage1_10[27],stage1_9[43]}
   );
   gpc606_5 gpc102 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[20],stage1_11[22],stage1_10[28],stage1_9[44]}
   );
   gpc606_5 gpc103 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[21],stage1_11[23],stage1_10[29],stage1_9[45]}
   );
   gpc606_5 gpc104 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[22],stage1_11[24],stage1_10[30],stage1_9[46]}
   );
   gpc606_5 gpc105 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[23],stage1_11[25],stage1_10[31],stage1_9[47]}
   );
   gpc606_5 gpc106 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[24],stage1_11[26],stage1_10[32],stage1_9[48]}
   );
   gpc606_5 gpc107 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[25],stage1_11[27],stage1_10[33],stage1_9[49]}
   );
   gpc606_5 gpc108 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[26],stage1_11[28],stage1_10[34],stage1_9[50]}
   );
   gpc606_5 gpc109 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[27],stage1_11[29],stage1_10[35],stage1_9[51]}
   );
   gpc606_5 gpc110 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[28],stage1_11[30],stage1_10[36],stage1_9[52]}
   );
   gpc606_5 gpc111 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[29],stage1_11[31],stage1_10[37],stage1_9[53]}
   );
   gpc606_5 gpc112 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[30],stage1_11[32],stage1_10[38],stage1_9[54]}
   );
   gpc606_5 gpc113 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[31],stage1_11[33],stage1_10[39],stage1_9[55]}
   );
   gpc606_5 gpc114 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[32],stage1_11[34],stage1_10[40],stage1_9[56]}
   );
   gpc606_5 gpc115 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[33],stage1_11[35],stage1_10[41],stage1_9[57]}
   );
   gpc606_5 gpc116 (
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[19],stage1_12[34],stage1_11[36],stage1_10[42]}
   );
   gpc606_5 gpc117 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[20],stage1_12[35],stage1_11[37],stage1_10[43]}
   );
   gpc615_5 gpc118 (
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106]},
      {stage0_11[114]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[21],stage1_12[36],stage1_11[38],stage1_10[44]}
   );
   gpc615_5 gpc119 (
      {stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111]},
      {stage0_11[115]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[22],stage1_12[37],stage1_11[39],stage1_10[45]}
   );
   gpc615_5 gpc120 (
      {stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116]},
      {stage0_11[116]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[23],stage1_12[38],stage1_11[40],stage1_10[46]}
   );
   gpc615_5 gpc121 (
      {stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121]},
      {stage0_11[117]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[24],stage1_12[39],stage1_11[41],stage1_10[47]}
   );
   gpc606_5 gpc122 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[6],stage1_13[25],stage1_12[40]}
   );
   gpc606_5 gpc123 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[7],stage1_13[26],stage1_12[41]}
   );
   gpc606_5 gpc124 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[8],stage1_13[27],stage1_12[42]}
   );
   gpc606_5 gpc125 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[9],stage1_13[28],stage1_12[43]}
   );
   gpc606_5 gpc126 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[4],stage1_14[10],stage1_13[29],stage1_12[44]}
   );
   gpc606_5 gpc127 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[5],stage1_14[11],stage1_13[30],stage1_12[45]}
   );
   gpc606_5 gpc128 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[6],stage1_14[12],stage1_13[31],stage1_12[46]}
   );
   gpc606_5 gpc129 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[7],stage1_14[13],stage1_13[32],stage1_12[47]}
   );
   gpc606_5 gpc130 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[8],stage1_14[14],stage1_13[33],stage1_12[48]}
   );
   gpc606_5 gpc131 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[9],stage1_14[15],stage1_13[34],stage1_12[49]}
   );
   gpc606_5 gpc132 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[10],stage1_14[16],stage1_13[35],stage1_12[50]}
   );
   gpc606_5 gpc133 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[11],stage1_14[17],stage1_13[36],stage1_12[51]}
   );
   gpc606_5 gpc134 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[12],stage1_14[18],stage1_13[37],stage1_12[52]}
   );
   gpc606_5 gpc135 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[13],stage1_14[19],stage1_13[38],stage1_12[53]}
   );
   gpc606_5 gpc136 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[14],stage1_14[20],stage1_13[39],stage1_12[54]}
   );
   gpc606_5 gpc137 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[15],stage1_15[15],stage1_14[21],stage1_13[40]}
   );
   gpc606_5 gpc138 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[16],stage1_15[16],stage1_14[22],stage1_13[41]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[17],stage1_15[17],stage1_14[23],stage1_13[42]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[18],stage1_15[18],stage1_14[24],stage1_13[43]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[19],stage1_15[19],stage1_14[25],stage1_13[44]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[20],stage1_15[20],stage1_14[26],stage1_13[45]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[21],stage1_15[21],stage1_14[27],stage1_13[46]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[22],stage1_15[22],stage1_14[28],stage1_13[47]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[23],stage1_15[23],stage1_14[29],stage1_13[48]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[24],stage1_15[24],stage1_14[30],stage1_13[49]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[25],stage1_15[25],stage1_14[31],stage1_13[50]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[26],stage1_15[26],stage1_14[32],stage1_13[51]}
   );
   gpc615_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76]},
      {stage0_14[90]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[27],stage1_15[27],stage1_14[33],stage1_13[52]}
   );
   gpc615_5 gpc150 (
      {stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_14[91]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[28],stage1_15[28],stage1_14[34],stage1_13[53]}
   );
   gpc615_5 gpc151 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86]},
      {stage0_14[92]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[29],stage1_15[29],stage1_14[35],stage1_13[54]}
   );
   gpc615_5 gpc152 (
      {stage0_13[87], stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91]},
      {stage0_14[93]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[30],stage1_15[30],stage1_14[36],stage1_13[55]}
   );
   gpc615_5 gpc153 (
      {stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95], stage0_13[96]},
      {stage0_14[94]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[31],stage1_15[31],stage1_14[37],stage1_13[56]}
   );
   gpc615_5 gpc154 (
      {stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_14[95]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[32],stage1_15[32],stage1_14[38],stage1_13[57]}
   );
   gpc615_5 gpc155 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106]},
      {stage0_14[96]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[33],stage1_15[33],stage1_14[39],stage1_13[58]}
   );
   gpc615_5 gpc156 (
      {stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_14[97]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[34],stage1_15[34],stage1_14[40],stage1_13[59]}
   );
   gpc615_5 gpc157 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116]},
      {stage0_14[98]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[35],stage1_15[35],stage1_14[41],stage1_13[60]}
   );
   gpc1_1 gpc158 (
      {stage0_0[99]},
      {stage1_0[17]}
   );
   gpc1_1 gpc159 (
      {stage0_0[100]},
      {stage1_0[18]}
   );
   gpc1_1 gpc160 (
      {stage0_0[101]},
      {stage1_0[19]}
   );
   gpc1_1 gpc161 (
      {stage0_0[102]},
      {stage1_0[20]}
   );
   gpc1_1 gpc162 (
      {stage0_0[103]},
      {stage1_0[21]}
   );
   gpc1_1 gpc163 (
      {stage0_0[104]},
      {stage1_0[22]}
   );
   gpc1_1 gpc164 (
      {stage0_0[105]},
      {stage1_0[23]}
   );
   gpc1_1 gpc165 (
      {stage0_0[106]},
      {stage1_0[24]}
   );
   gpc1_1 gpc166 (
      {stage0_0[107]},
      {stage1_0[25]}
   );
   gpc1_1 gpc167 (
      {stage0_0[108]},
      {stage1_0[26]}
   );
   gpc1_1 gpc168 (
      {stage0_0[109]},
      {stage1_0[27]}
   );
   gpc1_1 gpc169 (
      {stage0_0[110]},
      {stage1_0[28]}
   );
   gpc1_1 gpc170 (
      {stage0_0[111]},
      {stage1_0[29]}
   );
   gpc1_1 gpc171 (
      {stage0_0[112]},
      {stage1_0[30]}
   );
   gpc1_1 gpc172 (
      {stage0_0[113]},
      {stage1_0[31]}
   );
   gpc1_1 gpc173 (
      {stage0_0[114]},
      {stage1_0[32]}
   );
   gpc1_1 gpc174 (
      {stage0_0[115]},
      {stage1_0[33]}
   );
   gpc1_1 gpc175 (
      {stage0_0[116]},
      {stage1_0[34]}
   );
   gpc1_1 gpc176 (
      {stage0_0[117]},
      {stage1_0[35]}
   );
   gpc1_1 gpc177 (
      {stage0_0[118]},
      {stage1_0[36]}
   );
   gpc1_1 gpc178 (
      {stage0_0[119]},
      {stage1_0[37]}
   );
   gpc1_1 gpc179 (
      {stage0_0[120]},
      {stage1_0[38]}
   );
   gpc1_1 gpc180 (
      {stage0_0[121]},
      {stage1_0[39]}
   );
   gpc1_1 gpc181 (
      {stage0_0[122]},
      {stage1_0[40]}
   );
   gpc1_1 gpc182 (
      {stage0_0[123]},
      {stage1_0[41]}
   );
   gpc1_1 gpc183 (
      {stage0_0[124]},
      {stage1_0[42]}
   );
   gpc1_1 gpc184 (
      {stage0_0[125]},
      {stage1_0[43]}
   );
   gpc1_1 gpc185 (
      {stage0_0[126]},
      {stage1_0[44]}
   );
   gpc1_1 gpc186 (
      {stage0_0[127]},
      {stage1_0[45]}
   );
   gpc1_1 gpc187 (
      {stage0_1[96]},
      {stage1_1[32]}
   );
   gpc1_1 gpc188 (
      {stage0_1[97]},
      {stage1_1[33]}
   );
   gpc1_1 gpc189 (
      {stage0_1[98]},
      {stage1_1[34]}
   );
   gpc1_1 gpc190 (
      {stage0_1[99]},
      {stage1_1[35]}
   );
   gpc1_1 gpc191 (
      {stage0_1[100]},
      {stage1_1[36]}
   );
   gpc1_1 gpc192 (
      {stage0_1[101]},
      {stage1_1[37]}
   );
   gpc1_1 gpc193 (
      {stage0_1[102]},
      {stage1_1[38]}
   );
   gpc1_1 gpc194 (
      {stage0_1[103]},
      {stage1_1[39]}
   );
   gpc1_1 gpc195 (
      {stage0_1[104]},
      {stage1_1[40]}
   );
   gpc1_1 gpc196 (
      {stage0_1[105]},
      {stage1_1[41]}
   );
   gpc1_1 gpc197 (
      {stage0_1[106]},
      {stage1_1[42]}
   );
   gpc1_1 gpc198 (
      {stage0_1[107]},
      {stage1_1[43]}
   );
   gpc1_1 gpc199 (
      {stage0_1[108]},
      {stage1_1[44]}
   );
   gpc1_1 gpc200 (
      {stage0_1[109]},
      {stage1_1[45]}
   );
   gpc1_1 gpc201 (
      {stage0_1[110]},
      {stage1_1[46]}
   );
   gpc1_1 gpc202 (
      {stage0_1[111]},
      {stage1_1[47]}
   );
   gpc1_1 gpc203 (
      {stage0_1[112]},
      {stage1_1[48]}
   );
   gpc1_1 gpc204 (
      {stage0_1[113]},
      {stage1_1[49]}
   );
   gpc1_1 gpc205 (
      {stage0_1[114]},
      {stage1_1[50]}
   );
   gpc1_1 gpc206 (
      {stage0_1[115]},
      {stage1_1[51]}
   );
   gpc1_1 gpc207 (
      {stage0_1[116]},
      {stage1_1[52]}
   );
   gpc1_1 gpc208 (
      {stage0_1[117]},
      {stage1_1[53]}
   );
   gpc1_1 gpc209 (
      {stage0_1[118]},
      {stage1_1[54]}
   );
   gpc1_1 gpc210 (
      {stage0_1[119]},
      {stage1_1[55]}
   );
   gpc1_1 gpc211 (
      {stage0_1[120]},
      {stage1_1[56]}
   );
   gpc1_1 gpc212 (
      {stage0_1[121]},
      {stage1_1[57]}
   );
   gpc1_1 gpc213 (
      {stage0_1[122]},
      {stage1_1[58]}
   );
   gpc1_1 gpc214 (
      {stage0_1[123]},
      {stage1_1[59]}
   );
   gpc1_1 gpc215 (
      {stage0_1[124]},
      {stage1_1[60]}
   );
   gpc1_1 gpc216 (
      {stage0_1[125]},
      {stage1_1[61]}
   );
   gpc1_1 gpc217 (
      {stage0_1[126]},
      {stage1_1[62]}
   );
   gpc1_1 gpc218 (
      {stage0_1[127]},
      {stage1_1[63]}
   );
   gpc1_1 gpc219 (
      {stage0_2[126]},
      {stage1_2[37]}
   );
   gpc1_1 gpc220 (
      {stage0_2[127]},
      {stage1_2[38]}
   );
   gpc1_1 gpc221 (
      {stage0_3[122]},
      {stage1_3[43]}
   );
   gpc1_1 gpc222 (
      {stage0_3[123]},
      {stage1_3[44]}
   );
   gpc1_1 gpc223 (
      {stage0_3[124]},
      {stage1_3[45]}
   );
   gpc1_1 gpc224 (
      {stage0_3[125]},
      {stage1_3[46]}
   );
   gpc1_1 gpc225 (
      {stage0_3[126]},
      {stage1_3[47]}
   );
   gpc1_1 gpc226 (
      {stage0_3[127]},
      {stage1_3[48]}
   );
   gpc1_1 gpc227 (
      {stage0_4[126]},
      {stage1_4[58]}
   );
   gpc1_1 gpc228 (
      {stage0_4[127]},
      {stage1_4[59]}
   );
   gpc1_1 gpc229 (
      {stage0_7[108]},
      {stage1_7[45]}
   );
   gpc1_1 gpc230 (
      {stage0_7[109]},
      {stage1_7[46]}
   );
   gpc1_1 gpc231 (
      {stage0_7[110]},
      {stage1_7[47]}
   );
   gpc1_1 gpc232 (
      {stage0_7[111]},
      {stage1_7[48]}
   );
   gpc1_1 gpc233 (
      {stage0_7[112]},
      {stage1_7[49]}
   );
   gpc1_1 gpc234 (
      {stage0_7[113]},
      {stage1_7[50]}
   );
   gpc1_1 gpc235 (
      {stage0_7[114]},
      {stage1_7[51]}
   );
   gpc1_1 gpc236 (
      {stage0_7[115]},
      {stage1_7[52]}
   );
   gpc1_1 gpc237 (
      {stage0_7[116]},
      {stage1_7[53]}
   );
   gpc1_1 gpc238 (
      {stage0_7[117]},
      {stage1_7[54]}
   );
   gpc1_1 gpc239 (
      {stage0_7[118]},
      {stage1_7[55]}
   );
   gpc1_1 gpc240 (
      {stage0_7[119]},
      {stage1_7[56]}
   );
   gpc1_1 gpc241 (
      {stage0_7[120]},
      {stage1_7[57]}
   );
   gpc1_1 gpc242 (
      {stage0_7[121]},
      {stage1_7[58]}
   );
   gpc1_1 gpc243 (
      {stage0_7[122]},
      {stage1_7[59]}
   );
   gpc1_1 gpc244 (
      {stage0_7[123]},
      {stage1_7[60]}
   );
   gpc1_1 gpc245 (
      {stage0_7[124]},
      {stage1_7[61]}
   );
   gpc1_1 gpc246 (
      {stage0_7[125]},
      {stage1_7[62]}
   );
   gpc1_1 gpc247 (
      {stage0_7[126]},
      {stage1_7[63]}
   );
   gpc1_1 gpc248 (
      {stage0_7[127]},
      {stage1_7[64]}
   );
   gpc1_1 gpc249 (
      {stage0_8[126]},
      {stage1_8[54]}
   );
   gpc1_1 gpc250 (
      {stage0_8[127]},
      {stage1_8[55]}
   );
   gpc1_1 gpc251 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc252 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc253 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc254 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc255 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc256 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc257 (
      {stage0_11[118]},
      {stage1_11[42]}
   );
   gpc1_1 gpc258 (
      {stage0_11[119]},
      {stage1_11[43]}
   );
   gpc1_1 gpc259 (
      {stage0_11[120]},
      {stage1_11[44]}
   );
   gpc1_1 gpc260 (
      {stage0_11[121]},
      {stage1_11[45]}
   );
   gpc1_1 gpc261 (
      {stage0_11[122]},
      {stage1_11[46]}
   );
   gpc1_1 gpc262 (
      {stage0_11[123]},
      {stage1_11[47]}
   );
   gpc1_1 gpc263 (
      {stage0_11[124]},
      {stage1_11[48]}
   );
   gpc1_1 gpc264 (
      {stage0_11[125]},
      {stage1_11[49]}
   );
   gpc1_1 gpc265 (
      {stage0_11[126]},
      {stage1_11[50]}
   );
   gpc1_1 gpc266 (
      {stage0_11[127]},
      {stage1_11[51]}
   );
   gpc1_1 gpc267 (
      {stage0_12[126]},
      {stage1_12[55]}
   );
   gpc1_1 gpc268 (
      {stage0_12[127]},
      {stage1_12[56]}
   );
   gpc1_1 gpc269 (
      {stage0_13[117]},
      {stage1_13[61]}
   );
   gpc1_1 gpc270 (
      {stage0_13[118]},
      {stage1_13[62]}
   );
   gpc1_1 gpc271 (
      {stage0_13[119]},
      {stage1_13[63]}
   );
   gpc1_1 gpc272 (
      {stage0_13[120]},
      {stage1_13[64]}
   );
   gpc1_1 gpc273 (
      {stage0_13[121]},
      {stage1_13[65]}
   );
   gpc1_1 gpc274 (
      {stage0_13[122]},
      {stage1_13[66]}
   );
   gpc1_1 gpc275 (
      {stage0_13[123]},
      {stage1_13[67]}
   );
   gpc1_1 gpc276 (
      {stage0_13[124]},
      {stage1_13[68]}
   );
   gpc1_1 gpc277 (
      {stage0_13[125]},
      {stage1_13[69]}
   );
   gpc1_1 gpc278 (
      {stage0_13[126]},
      {stage1_13[70]}
   );
   gpc1_1 gpc279 (
      {stage0_13[127]},
      {stage1_13[71]}
   );
   gpc1_1 gpc280 (
      {stage0_14[99]},
      {stage1_14[42]}
   );
   gpc1_1 gpc281 (
      {stage0_14[100]},
      {stage1_14[43]}
   );
   gpc1_1 gpc282 (
      {stage0_14[101]},
      {stage1_14[44]}
   );
   gpc1_1 gpc283 (
      {stage0_14[102]},
      {stage1_14[45]}
   );
   gpc1_1 gpc284 (
      {stage0_14[103]},
      {stage1_14[46]}
   );
   gpc1_1 gpc285 (
      {stage0_14[104]},
      {stage1_14[47]}
   );
   gpc1_1 gpc286 (
      {stage0_14[105]},
      {stage1_14[48]}
   );
   gpc1_1 gpc287 (
      {stage0_14[106]},
      {stage1_14[49]}
   );
   gpc1_1 gpc288 (
      {stage0_14[107]},
      {stage1_14[50]}
   );
   gpc1_1 gpc289 (
      {stage0_14[108]},
      {stage1_14[51]}
   );
   gpc1_1 gpc290 (
      {stage0_14[109]},
      {stage1_14[52]}
   );
   gpc1_1 gpc291 (
      {stage0_14[110]},
      {stage1_14[53]}
   );
   gpc1_1 gpc292 (
      {stage0_14[111]},
      {stage1_14[54]}
   );
   gpc1_1 gpc293 (
      {stage0_14[112]},
      {stage1_14[55]}
   );
   gpc1_1 gpc294 (
      {stage0_14[113]},
      {stage1_14[56]}
   );
   gpc1_1 gpc295 (
      {stage0_14[114]},
      {stage1_14[57]}
   );
   gpc1_1 gpc296 (
      {stage0_14[115]},
      {stage1_14[58]}
   );
   gpc1_1 gpc297 (
      {stage0_14[116]},
      {stage1_14[59]}
   );
   gpc1_1 gpc298 (
      {stage0_14[117]},
      {stage1_14[60]}
   );
   gpc1_1 gpc299 (
      {stage0_14[118]},
      {stage1_14[61]}
   );
   gpc1_1 gpc300 (
      {stage0_14[119]},
      {stage1_14[62]}
   );
   gpc1_1 gpc301 (
      {stage0_14[120]},
      {stage1_14[63]}
   );
   gpc1_1 gpc302 (
      {stage0_14[121]},
      {stage1_14[64]}
   );
   gpc1_1 gpc303 (
      {stage0_14[122]},
      {stage1_14[65]}
   );
   gpc1_1 gpc304 (
      {stage0_14[123]},
      {stage1_14[66]}
   );
   gpc1_1 gpc305 (
      {stage0_14[124]},
      {stage1_14[67]}
   );
   gpc1_1 gpc306 (
      {stage0_14[125]},
      {stage1_14[68]}
   );
   gpc1_1 gpc307 (
      {stage0_14[126]},
      {stage1_14[69]}
   );
   gpc1_1 gpc308 (
      {stage0_14[127]},
      {stage1_14[70]}
   );
   gpc1_1 gpc309 (
      {stage0_15[126]},
      {stage1_15[36]}
   );
   gpc1_1 gpc310 (
      {stage0_15[127]},
      {stage1_15[37]}
   );
   gpc1163_5 gpc311 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc312 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc313 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc314 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc315 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc316 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc317 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc319 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc320 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc321 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1406_5 gpc322 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[0]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc615_5 gpc323 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[26]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc615_5 gpc324 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[27]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc325 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage2_6[0],stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc326 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[7]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[4],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc327 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[8]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[5],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc328 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[9]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc329 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[10]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc330 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[11]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc606_5 gpc331 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[5],stage2_6[6],stage2_5[9],stage2_4[20]}
   );
   gpc606_5 gpc332 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[6],stage2_6[7],stage2_5[10],stage2_4[21]}
   );
   gpc606_5 gpc333 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[7],stage2_6[8],stage2_5[11],stage2_4[22]}
   );
   gpc606_5 gpc334 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[8],stage2_6[9],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc335 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[9],stage2_6[10],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc336 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[10],stage2_6[11],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc337 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[11],stage2_6[12],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc338 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[12],stage2_6[13],stage2_5[16],stage2_4[27]}
   );
   gpc207_4 gpc339 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[8],stage2_7[13],stage2_6[14],stage2_5[17]}
   );
   gpc606_5 gpc340 (
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[9],stage2_7[14],stage2_6[15],stage2_5[18]}
   );
   gpc606_5 gpc341 (
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[10],stage2_7[15],stage2_6[16],stage2_5[19]}
   );
   gpc615_5 gpc342 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[2],stage2_8[11],stage2_7[16]}
   );
   gpc615_5 gpc343 (
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[3],stage2_8[12],stage2_7[17]}
   );
   gpc615_5 gpc344 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[4],stage2_8[13],stage2_7[18]}
   );
   gpc615_5 gpc345 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[5],stage2_8[14],stage2_7[19]}
   );
   gpc615_5 gpc346 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[6],stage2_8[15],stage2_7[20]}
   );
   gpc615_5 gpc347 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[7],stage2_8[16],stage2_7[21]}
   );
   gpc615_5 gpc348 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[8],stage2_8[17],stage2_7[22]}
   );
   gpc615_5 gpc349 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[9],stage2_8[18],stage2_7[23]}
   );
   gpc615_5 gpc350 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[10],stage2_8[19],stage2_7[24]}
   );
   gpc606_5 gpc351 (
      {stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[9],stage2_10[9],stage2_9[11],stage2_8[20]}
   );
   gpc606_5 gpc352 (
      {stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[10],stage2_10[10],stage2_9[12],stage2_8[21]}
   );
   gpc606_5 gpc353 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[11],stage2_10[11],stage2_9[13],stage2_8[22]}
   );
   gpc606_5 gpc354 (
      {stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[12],stage2_10[12],stage2_9[14],stage2_8[23]}
   );
   gpc606_5 gpc355 (
      {stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[13],stage2_10[13],stage2_9[15],stage2_8[24]}
   );
   gpc606_5 gpc356 (
      {stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[14],stage2_10[14],stage2_9[16],stage2_8[25]}
   );
   gpc615_5 gpc357 (
      {stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_9[54]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[15],stage2_10[15],stage2_9[17],stage2_8[26]}
   );
   gpc615_5 gpc358 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_9[55]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[16],stage2_10[16],stage2_9[18],stage2_8[27]}
   );
   gpc606_5 gpc359 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[8],stage2_11[17],stage2_10[17]}
   );
   gpc615_5 gpc360 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[9],stage2_11[18]}
   );
   gpc615_5 gpc361 (
      {stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[10],stage2_11[19]}
   );
   gpc615_5 gpc362 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[11],stage2_11[20]}
   );
   gpc615_5 gpc363 (
      {stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[12],stage2_11[21]}
   );
   gpc615_5 gpc364 (
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_12[10]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[13],stage2_11[22]}
   );
   gpc615_5 gpc365 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_12[11]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[14],stage2_11[23]}
   );
   gpc615_5 gpc366 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[12]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[7],stage2_12[15],stage2_11[24]}
   );
   gpc615_5 gpc367 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[13]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[8],stage2_12[16],stage2_11[25]}
   );
   gpc207_4 gpc368 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19], stage1_12[20]},
      {stage1_14[0], stage1_14[1]},
      {stage2_15[8],stage2_14[9],stage2_13[9],stage2_12[17]}
   );
   gpc606_5 gpc369 (
      {stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25], stage1_12[26]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[0],stage2_15[9],stage2_14[10],stage2_13[10],stage2_12[18]}
   );
   gpc606_5 gpc370 (
      {stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[1],stage2_15[10],stage2_14[11],stage2_13[11],stage2_12[19]}
   );
   gpc606_5 gpc371 (
      {stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[2],stage2_15[11],stage2_14[12],stage2_13[12],stage2_12[20]}
   );
   gpc606_5 gpc372 (
      {stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[3],stage2_15[12],stage2_14[13],stage2_13[13],stage2_12[21]}
   );
   gpc606_5 gpc373 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[4],stage2_15[13],stage2_14[14],stage2_13[14],stage2_12[22]}
   );
   gpc606_5 gpc374 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[15],stage2_13[15]}
   );
   gpc606_5 gpc375 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[16],stage2_13[16]}
   );
   gpc606_5 gpc376 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[17],stage2_13[17]}
   );
   gpc606_5 gpc377 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[18],stage2_13[18]}
   );
   gpc606_5 gpc378 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[19]}
   );
   gpc606_5 gpc379 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[20]}
   );
   gpc606_5 gpc380 (
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[21]}
   );
   gpc615_5 gpc381 (
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_15[24]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[22]}
   );
   gpc615_5 gpc382 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[25]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[23]}
   );
   gpc615_5 gpc383 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30]},
      {stage1_16[30]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23]}
   );
   gpc615_5 gpc384 (
      {stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[31]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24]}
   );
   gpc1_1 gpc385 (
      {stage1_0[42]},
      {stage2_0[11]}
   );
   gpc1_1 gpc386 (
      {stage1_0[43]},
      {stage2_0[12]}
   );
   gpc1_1 gpc387 (
      {stage1_0[44]},
      {stage2_0[13]}
   );
   gpc1_1 gpc388 (
      {stage1_0[45]},
      {stage2_0[14]}
   );
   gpc1_1 gpc389 (
      {stage1_2[34]},
      {stage2_2[15]}
   );
   gpc1_1 gpc390 (
      {stage1_2[35]},
      {stage2_2[16]}
   );
   gpc1_1 gpc391 (
      {stage1_2[36]},
      {stage2_2[17]}
   );
   gpc1_1 gpc392 (
      {stage1_2[37]},
      {stage2_2[18]}
   );
   gpc1_1 gpc393 (
      {stage1_2[38]},
      {stage2_2[19]}
   );
   gpc1_1 gpc394 (
      {stage1_5[49]},
      {stage2_5[20]}
   );
   gpc1_1 gpc395 (
      {stage1_5[50]},
      {stage2_5[21]}
   );
   gpc1_1 gpc396 (
      {stage1_5[51]},
      {stage2_5[22]}
   );
   gpc1_1 gpc397 (
      {stage1_5[52]},
      {stage2_5[23]}
   );
   gpc1_1 gpc398 (
      {stage1_5[53]},
      {stage2_5[24]}
   );
   gpc1_1 gpc399 (
      {stage1_5[54]},
      {stage2_5[25]}
   );
   gpc1_1 gpc400 (
      {stage1_5[55]},
      {stage2_5[26]}
   );
   gpc1_1 gpc401 (
      {stage1_5[56]},
      {stage2_5[27]}
   );
   gpc1_1 gpc402 (
      {stage1_7[59]},
      {stage2_7[25]}
   );
   gpc1_1 gpc403 (
      {stage1_7[60]},
      {stage2_7[26]}
   );
   gpc1_1 gpc404 (
      {stage1_7[61]},
      {stage2_7[27]}
   );
   gpc1_1 gpc405 (
      {stage1_7[62]},
      {stage2_7[28]}
   );
   gpc1_1 gpc406 (
      {stage1_7[63]},
      {stage2_7[29]}
   );
   gpc1_1 gpc407 (
      {stage1_7[64]},
      {stage2_7[30]}
   );
   gpc1_1 gpc408 (
      {stage1_8[55]},
      {stage2_8[28]}
   );
   gpc1_1 gpc409 (
      {stage1_9[56]},
      {stage2_9[19]}
   );
   gpc1_1 gpc410 (
      {stage1_9[57]},
      {stage2_9[20]}
   );
   gpc1_1 gpc411 (
      {stage1_11[40]},
      {stage2_11[26]}
   );
   gpc1_1 gpc412 (
      {stage1_11[41]},
      {stage2_11[27]}
   );
   gpc1_1 gpc413 (
      {stage1_11[42]},
      {stage2_11[28]}
   );
   gpc1_1 gpc414 (
      {stage1_11[43]},
      {stage2_11[29]}
   );
   gpc1_1 gpc415 (
      {stage1_11[44]},
      {stage2_11[30]}
   );
   gpc1_1 gpc416 (
      {stage1_11[45]},
      {stage2_11[31]}
   );
   gpc1_1 gpc417 (
      {stage1_11[46]},
      {stage2_11[32]}
   );
   gpc1_1 gpc418 (
      {stage1_11[47]},
      {stage2_11[33]}
   );
   gpc1_1 gpc419 (
      {stage1_11[48]},
      {stage2_11[34]}
   );
   gpc1_1 gpc420 (
      {stage1_11[49]},
      {stage2_11[35]}
   );
   gpc1_1 gpc421 (
      {stage1_11[50]},
      {stage2_11[36]}
   );
   gpc1_1 gpc422 (
      {stage1_11[51]},
      {stage2_11[37]}
   );
   gpc1_1 gpc423 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc424 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc425 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc426 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc427 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc428 (
      {stage1_12[56]},
      {stage2_12[28]}
   );
   gpc1_1 gpc429 (
      {stage1_14[60]},
      {stage2_14[24]}
   );
   gpc1_1 gpc430 (
      {stage1_14[61]},
      {stage2_14[25]}
   );
   gpc1_1 gpc431 (
      {stage1_14[62]},
      {stage2_14[26]}
   );
   gpc1_1 gpc432 (
      {stage1_14[63]},
      {stage2_14[27]}
   );
   gpc1_1 gpc433 (
      {stage1_14[64]},
      {stage2_14[28]}
   );
   gpc1_1 gpc434 (
      {stage1_14[65]},
      {stage2_14[29]}
   );
   gpc1_1 gpc435 (
      {stage1_14[66]},
      {stage2_14[30]}
   );
   gpc1_1 gpc436 (
      {stage1_14[67]},
      {stage2_14[31]}
   );
   gpc1_1 gpc437 (
      {stage1_14[68]},
      {stage2_14[32]}
   );
   gpc1_1 gpc438 (
      {stage1_14[69]},
      {stage2_14[33]}
   );
   gpc1_1 gpc439 (
      {stage1_14[70]},
      {stage2_14[34]}
   );
   gpc1_1 gpc440 (
      {stage1_15[36]},
      {stage2_15[25]}
   );
   gpc1_1 gpc441 (
      {stage1_15[37]},
      {stage2_15[26]}
   );
   gpc1_1 gpc442 (
      {stage1_16[32]},
      {stage2_16[16]}
   );
   gpc1_1 gpc443 (
      {stage1_16[33]},
      {stage2_16[17]}
   );
   gpc1_1 gpc444 (
      {stage1_16[34]},
      {stage2_16[18]}
   );
   gpc1_1 gpc445 (
      {stage1_16[35]},
      {stage2_16[19]}
   );
   gpc1_1 gpc446 (
      {stage1_17[12]},
      {stage2_17[11]}
   );
   gpc1_1 gpc447 (
      {stage1_17[13]},
      {stage2_17[12]}
   );
   gpc1_1 gpc448 (
      {stage1_17[14]},
      {stage2_17[13]}
   );
   gpc1_1 gpc449 (
      {stage1_17[15]},
      {stage2_17[14]}
   );
   gpc1_1 gpc450 (
      {stage1_17[16]},
      {stage2_17[15]}
   );
   gpc1_1 gpc451 (
      {stage1_17[17]},
      {stage2_17[16]}
   );
   gpc1_1 gpc452 (
      {stage1_17[18]},
      {stage2_17[17]}
   );
   gpc1_1 gpc453 (
      {stage1_17[19]},
      {stage2_17[18]}
   );
   gpc1_1 gpc454 (
      {stage1_17[20]},
      {stage2_17[19]}
   );
   gpc606_5 gpc455 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc456 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc615_5 gpc457 (
      {stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc458 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc1163_5 gpc459 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[4]}
   );
   gpc606_5 gpc460 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[4],stage3_5[5]}
   );
   gpc615_5 gpc461 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_6[2]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc615_5 gpc462 (
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_6[3]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc615_5 gpc463 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_6[4]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc615_5 gpc464 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27]},
      {stage2_6[5]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[4],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc465 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[5],stage3_7[7],stage3_6[9]}
   );
   gpc615_5 gpc466 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_7[30]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[6],stage3_7[8],stage3_6[10]}
   );
   gpc606_5 gpc467 (
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[2],stage3_9[7],stage3_8[7]}
   );
   gpc606_5 gpc468 (
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[3],stage3_9[8],stage3_8[8]}
   );
   gpc1163_5 gpc469 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[2],stage3_10[4],stage3_9[9]}
   );
   gpc606_5 gpc470 (
      {stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage3_13[1],stage3_12[3],stage3_11[3],stage3_10[5],stage3_9[10]}
   );
   gpc606_5 gpc471 (
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage3_13[2],stage3_12[4],stage3_11[4],stage3_10[6],stage3_9[11]}
   );
   gpc606_5 gpc472 (
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage3_13[3],stage3_12[5],stage3_11[5],stage3_10[7],stage3_9[12]}
   );
   gpc615_5 gpc473 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_12[1]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[6],stage3_11[6]}
   );
   gpc615_5 gpc474 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[7],stage3_11[7]}
   );
   gpc606_5 gpc475 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[8]}
   );
   gpc606_5 gpc476 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[9]}
   );
   gpc606_5 gpc477 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[10]}
   );
   gpc606_5 gpc478 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[11]}
   );
   gpc606_5 gpc479 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[6],stage3_14[6],stage3_13[10]}
   );
   gpc1163_5 gpc480 (
      {stage2_14[24], stage2_14[25], stage2_14[26]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc481 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[1]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[0],stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[8]}
   );
   gpc615_5 gpc482 (
      {stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_16[2]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[1],stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[9]}
   );
   gpc615_5 gpc483 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26]},
      {stage2_16[3]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[2],stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[10]}
   );
   gpc606_5 gpc484 (
      {stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[3],stage3_18[4],stage3_17[5],stage3_16[9]}
   );
   gpc1_1 gpc485 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc486 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc487 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc488 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc489 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc490 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc491 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc492 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc493 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc494 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc495 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc496 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc497 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc498 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc499 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc500 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc501 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc502 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc503 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc504 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc505 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc506 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc507 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc508 (
      {stage2_2[10]},
      {stage3_2[3]}
   );
   gpc1_1 gpc509 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc510 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc511 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc512 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc513 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc514 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc515 (
      {stage2_2[17]},
      {stage3_2[10]}
   );
   gpc1_1 gpc516 (
      {stage2_2[18]},
      {stage3_2[11]}
   );
   gpc1_1 gpc517 (
      {stage2_2[19]},
      {stage3_2[12]}
   );
   gpc1_1 gpc518 (
      {stage2_3[14]},
      {stage3_3[5]}
   );
   gpc1_1 gpc519 (
      {stage2_3[15]},
      {stage3_3[6]}
   );
   gpc1_1 gpc520 (
      {stage2_3[16]},
      {stage3_3[7]}
   );
   gpc1_1 gpc521 (
      {stage2_3[17]},
      {stage3_3[8]}
   );
   gpc1_1 gpc522 (
      {stage2_3[18]},
      {stage3_3[9]}
   );
   gpc1_1 gpc523 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc524 (
      {stage2_4[24]},
      {stage3_4[5]}
   );
   gpc1_1 gpc525 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc526 (
      {stage2_4[26]},
      {stage3_4[7]}
   );
   gpc1_1 gpc527 (
      {stage2_4[27]},
      {stage3_4[8]}
   );
   gpc1_1 gpc528 (
      {stage2_8[24]},
      {stage3_8[9]}
   );
   gpc1_1 gpc529 (
      {stage2_8[25]},
      {stage3_8[10]}
   );
   gpc1_1 gpc530 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc531 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc532 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc533 (
      {stage2_11[29]},
      {stage3_11[8]}
   );
   gpc1_1 gpc534 (
      {stage2_11[30]},
      {stage3_11[9]}
   );
   gpc1_1 gpc535 (
      {stage2_11[31]},
      {stage3_11[10]}
   );
   gpc1_1 gpc536 (
      {stage2_11[32]},
      {stage3_11[11]}
   );
   gpc1_1 gpc537 (
      {stage2_11[33]},
      {stage3_11[12]}
   );
   gpc1_1 gpc538 (
      {stage2_11[34]},
      {stage3_11[13]}
   );
   gpc1_1 gpc539 (
      {stage2_11[35]},
      {stage3_11[14]}
   );
   gpc1_1 gpc540 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc541 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc542 (
      {stage2_12[27]},
      {stage3_12[12]}
   );
   gpc1_1 gpc543 (
      {stage2_12[28]},
      {stage3_12[13]}
   );
   gpc1_1 gpc544 (
      {stage2_13[18]},
      {stage3_13[11]}
   );
   gpc1_1 gpc545 (
      {stage2_14[27]},
      {stage3_14[8]}
   );
   gpc1_1 gpc546 (
      {stage2_14[28]},
      {stage3_14[9]}
   );
   gpc1_1 gpc547 (
      {stage2_14[29]},
      {stage3_14[10]}
   );
   gpc1_1 gpc548 (
      {stage2_14[30]},
      {stage3_14[11]}
   );
   gpc1_1 gpc549 (
      {stage2_14[31]},
      {stage3_14[12]}
   );
   gpc1_1 gpc550 (
      {stage2_14[32]},
      {stage3_14[13]}
   );
   gpc1_1 gpc551 (
      {stage2_14[33]},
      {stage3_14[14]}
   );
   gpc1_1 gpc552 (
      {stage2_14[34]},
      {stage3_14[15]}
   );
   gpc1_1 gpc553 (
      {stage2_16[10]},
      {stage3_16[10]}
   );
   gpc1_1 gpc554 (
      {stage2_16[11]},
      {stage3_16[11]}
   );
   gpc1_1 gpc555 (
      {stage2_16[12]},
      {stage3_16[12]}
   );
   gpc1_1 gpc556 (
      {stage2_16[13]},
      {stage3_16[13]}
   );
   gpc1_1 gpc557 (
      {stage2_16[14]},
      {stage3_16[14]}
   );
   gpc1_1 gpc558 (
      {stage2_16[15]},
      {stage3_16[15]}
   );
   gpc1_1 gpc559 (
      {stage2_16[16]},
      {stage3_16[16]}
   );
   gpc1_1 gpc560 (
      {stage2_16[17]},
      {stage3_16[17]}
   );
   gpc1_1 gpc561 (
      {stage2_16[18]},
      {stage3_16[18]}
   );
   gpc1_1 gpc562 (
      {stage2_16[19]},
      {stage3_16[19]}
   );
   gpc1_1 gpc563 (
      {stage2_17[19]},
      {stage3_17[6]}
   );
   gpc1_1 gpc564 (
      {stage2_18[6]},
      {stage3_18[5]}
   );
   gpc1_1 gpc565 (
      {stage2_19[0]},
      {stage3_19[4]}
   );
   gpc1_1 gpc566 (
      {stage2_19[1]},
      {stage3_19[5]}
   );
   gpc606_5 gpc567 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc568 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10]},
      {stage3_1[0]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1163_5 gpc569 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc570 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc615_5 gpc571 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc572 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[2],stage4_7[3],stage4_6[3]}
   );
   gpc606_5 gpc573 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[2],stage4_9[3]}
   );
   gpc615_5 gpc574 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[3],stage4_9[4]}
   );
   gpc606_5 gpc575 (
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[4]}
   );
   gpc615_5 gpc576 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16]},
      {stage3_12[6]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc577 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc578 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[5]}
   );
   gpc615_5 gpc579 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[4]}
   );
   gpc615_5 gpc580 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[7]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[5]}
   );
   gpc606_5 gpc581 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4]}
   );
   gpc606_5 gpc582 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[3],stage4_17[4]}
   );
   gpc1_1 gpc583 (
      {stage3_0[11]},
      {stage4_0[2]}
   );
   gpc1_1 gpc584 (
      {stage3_0[12]},
      {stage4_0[3]}
   );
   gpc1_1 gpc585 (
      {stage3_0[13]},
      {stage4_0[4]}
   );
   gpc1_1 gpc586 (
      {stage3_0[14]},
      {stage4_0[5]}
   );
   gpc1_1 gpc587 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc588 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc589 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc590 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc591 (
      {stage3_1[5]},
      {stage4_1[6]}
   );
   gpc1_1 gpc592 (
      {stage3_1[6]},
      {stage4_1[7]}
   );
   gpc1_1 gpc593 (
      {stage3_1[7]},
      {stage4_1[8]}
   );
   gpc1_1 gpc594 (
      {stage3_1[8]},
      {stage4_1[9]}
   );
   gpc1_1 gpc595 (
      {stage3_2[12]},
      {stage4_2[2]}
   );
   gpc1_1 gpc596 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc597 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc598 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc599 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc600 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc601 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc602 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc603 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc604 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc605 (
      {stage3_4[7]},
      {stage4_4[4]}
   );
   gpc1_1 gpc606 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc607 (
      {stage3_5[7]},
      {stage4_5[2]}
   );
   gpc1_1 gpc608 (
      {stage3_5[8]},
      {stage4_5[3]}
   );
   gpc1_1 gpc609 (
      {stage3_5[9]},
      {stage4_5[4]}
   );
   gpc1_1 gpc610 (
      {stage3_7[8]},
      {stage4_7[4]}
   );
   gpc1_1 gpc611 (
      {stage3_8[12]},
      {stage4_8[3]}
   );
   gpc1_1 gpc612 (
      {stage3_8[13]},
      {stage4_8[4]}
   );
   gpc1_1 gpc613 (
      {stage3_9[11]},
      {stage4_9[5]}
   );
   gpc1_1 gpc614 (
      {stage3_9[12]},
      {stage4_9[6]}
   );
   gpc1_1 gpc615 (
      {stage3_10[7]},
      {stage4_10[5]}
   );
   gpc1_1 gpc616 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc617 (
      {stage3_15[8]},
      {stage4_15[5]}
   );
   gpc1_1 gpc618 (
      {stage3_15[9]},
      {stage4_15[6]}
   );
   gpc1_1 gpc619 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc620 (
      {stage3_16[18]},
      {stage4_16[5]}
   );
   gpc1_1 gpc621 (
      {stage3_16[19]},
      {stage4_16[6]}
   );
   gpc1_1 gpc622 (
      {stage3_17[6]},
      {stage4_17[5]}
   );
   gpc1_1 gpc623 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc2135_5 gpc624 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1415_5 gpc625 (
      {stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6], stage4_1[7]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1415_5 gpc626 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc627 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[1]}
   );
   gpc606_5 gpc628 (
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc135_4 gpc629 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1]}
   );
   gpc1343_5 gpc630 (
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0], stage4_19[1], 1'b0, 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1_1 gpc631 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc632 (
      {stage4_1[8]},
      {stage5_1[2]}
   );
   gpc1_1 gpc633 (
      {stage4_1[9]},
      {stage5_1[3]}
   );
   gpc1_1 gpc634 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc635 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc636 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc637 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc638 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc639 (
      {stage4_3[10]},
      {stage5_3[6]}
   );
   gpc1_1 gpc640 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc641 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc642 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc643 (
      {stage4_5[4]},
      {stage5_5[5]}
   );
   gpc1_1 gpc644 (
      {stage4_7[1]},
      {stage5_7[1]}
   );
   gpc1_1 gpc645 (
      {stage4_7[2]},
      {stage5_7[2]}
   );
   gpc1_1 gpc646 (
      {stage4_7[3]},
      {stage5_7[3]}
   );
   gpc1_1 gpc647 (
      {stage4_7[4]},
      {stage5_7[4]}
   );
   gpc1_1 gpc648 (
      {stage4_9[1]},
      {stage5_9[1]}
   );
   gpc1_1 gpc649 (
      {stage4_9[2]},
      {stage5_9[2]}
   );
   gpc1_1 gpc650 (
      {stage4_9[3]},
      {stage5_9[3]}
   );
   gpc1_1 gpc651 (
      {stage4_9[4]},
      {stage5_9[4]}
   );
   gpc1_1 gpc652 (
      {stage4_9[5]},
      {stage5_9[5]}
   );
   gpc1_1 gpc653 (
      {stage4_9[6]},
      {stage5_9[6]}
   );
   gpc1_1 gpc654 (
      {stage4_11[0]},
      {stage5_11[1]}
   );
   gpc1_1 gpc655 (
      {stage4_11[1]},
      {stage5_11[2]}
   );
   gpc1_1 gpc656 (
      {stage4_11[2]},
      {stage5_11[3]}
   );
   gpc1_1 gpc657 (
      {stage4_11[3]},
      {stage5_11[4]}
   );
   gpc1_1 gpc658 (
      {stage4_13[0]},
      {stage5_13[1]}
   );
   gpc1_1 gpc659 (
      {stage4_13[1]},
      {stage5_13[2]}
   );
   gpc1_1 gpc660 (
      {stage4_13[2]},
      {stage5_13[3]}
   );
   gpc1_1 gpc661 (
      {stage4_13[3]},
      {stage5_13[4]}
   );
   gpc1_1 gpc662 (
      {stage4_13[4]},
      {stage5_13[5]}
   );
   gpc1_1 gpc663 (
      {stage4_13[5]},
      {stage5_13[6]}
   );
   gpc1_1 gpc664 (
      {stage4_15[5]},
      {stage5_15[2]}
   );
   gpc1_1 gpc665 (
      {stage4_15[6]},
      {stage5_15[3]}
   );
   gpc1_1 gpc666 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc667 (
      {stage4_16[3]},
      {stage5_16[2]}
   );
   gpc1_1 gpc668 (
      {stage4_16[4]},
      {stage5_16[3]}
   );
   gpc1_1 gpc669 (
      {stage4_16[5]},
      {stage5_16[4]}
   );
   gpc1_1 gpc670 (
      {stage4_16[6]},
      {stage5_16[5]}
   );
   gpc1_1 gpc671 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc672 (
      {stage4_17[2]},
      {stage5_17[2]}
   );
   gpc1_1 gpc673 (
      {stage4_17[3]},
      {stage5_17[3]}
   );
   gpc1_1 gpc674 (
      {stage4_17[4]},
      {stage5_17[4]}
   );
   gpc1_1 gpc675 (
      {stage4_17[5]},
      {stage5_17[5]}
   );
   gpc1_1 gpc676 (
      {stage4_18[3]},
      {stage5_18[2]}
   );
   gpc2223_5 gpc677 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1]},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc678 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc679 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1]}
   );
   gpc615_5 gpc680 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1]}
   );
   gpc615_5 gpc681 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc682 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2], 1'b0},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc1_1 gpc683 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc684 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc685 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc686 (
      {stage5_2[2]},
      {stage6_2[1]}
   );
   gpc1_1 gpc687 (
      {stage5_6[0]},
      {stage6_6[1]}
   );
   gpc1_1 gpc688 (
      {stage5_8[1]},
      {stage6_8[1]}
   );
   gpc1_1 gpc689 (
      {stage5_9[6]},
      {stage6_9[1]}
   );
   gpc1_1 gpc690 (
      {stage5_10[0]},
      {stage6_10[1]}
   );
   gpc1_1 gpc691 (
      {stage5_12[1]},
      {stage6_12[1]}
   );
   gpc1_1 gpc692 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc693 (
      {stage5_14[0]},
      {stage6_14[1]}
   );
   gpc1_1 gpc694 (
      {stage5_20[0]},
      {stage6_20[1]}
   );
   gpc1_1 gpc695 (
      {stage5_21[0]},
      {stage6_21[0]}
   );
   gpc1_1 gpc696 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
endmodule
module rowadder2_1_23(input [22:0] src0, input [22:0] src1, output [23:0] dst0);
    wire [22:0] gene;
    wire [22:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[22:20]}),
        .S({1'h0, prop[22:20]})
    );
    assign dst0 = {carryout[22], out[22:0]};
endmodule


module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor2_1_128_16 compressor2_1_128_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h949fbf79ea7f5e71d1e960bbb99bb0749613bf1e2ebd5ba8ae6edb7a6945d48b65766e4e4a6b6d7a81e7afb98b74ce7862999e780f3f5bbf541c3b100947743447ee72a17c0217b9cee20d85362819359dcd5b0652aca41586ff851d0be6143b29497394a92b2888e58129abe16b6aafac9d5d963943c941329bb4edbbc19e3e557d51dbcde4e5dfcf7cd20a8d94919669349645e07f6fe716d9af742603d426c03bcbd34b517ca8f98aaf6850f40cd4115f407a097f4f39c2e84d7f06b7535386ea67098af8c1e1f7828bd3989c22eeb093ebc784826763d8b2027a40abd42e4f8145e672def26da8749cc8880edca5f0a025e35b96b0e09c6178b3ced994db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5ecc14923e572a95345790621b7704022cfd4427561eca21528b0d4be977453aefcebf4ea85630230fb25ad6ac6478b0af5a19011dfc2fa080ca981557f6080181765bb72dfc63e30f6a59aae43c69dfee699395534741de54e1002921eb948ef93bf2c576d5868adbec78469fca62647c95cc8ff470e48ec9e7300780273b887ed8ee78784292cab9a69152acf491487c40420a715202bee098ae4fdb610ed54bf1471ba1a7c5e9b325213fd21dfac91163183db97389a63fc9eeacd62a1f48a09e3ed0d12bcc7e1efc54b54d0148261d14e79a14788df827b37c1b9977c8f9bb6501a9faef1bc5f6a9c7f74ed6cbbeb3bdadfbd73eba0e003d82b0571fef2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4f01c22d535ffaf5aad7b9196cd9361d97fa1e98395f0811856fe51f944ecc96231672240e84489cc2cd6e63fd0bd4dd045e3df760bcaaae73b70fe21056ea39f3fc8075e4d7511ae6d5352a94be54fe79006401831e7525ec9581e0c77c00f86a1fccc9c085695091051bdaf1a1c163e1db91d87284077dbc6b62c8d7ade8d83159113573ac3dc26a3f8d226cf5749139515c609b1e2f67aa8edb45c1198dc4993199b3b9364622d488d78f4ff33f9bc25304d4c3f970029c08f45ff6b8c291a3eb423e25ccb6f1b49f62a7f8de0d429bc295bfe2950f5f724266f88639e3ba99e72ba8c903776ad919e1b7f643f5684e45915c65c892fa7ea27a52e2d5b508;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd48320f4061a6449d0562eefb7352d903e25ed15d347b84eeee15cdfcdc64ebb6f281f245ee917da58691312a44b5f336bdb5ef0e98a7226dc290f15b9772ee67534226a4d833e61a27dca819b8ce6d45c47e6142e1fa009a5812067f9fdd867e946979109ccd906b48c18d6efdb9f4c3cc60b0949d58f6aefe3d7b14db20fde39c72dca5edafb69fba2f170941947cd6f00dd0c2be28bd871979470ff1b1747432511eb827402c1f5ac8398d731876084246cd786891bb12198ae9b4713d20f5914a5257f56e43917fe2b081ff4046fbb651e844d1884a43f54c0ba121f816c0227933fd2e59f916f6c2d6fe50f1cf91548168b937ec3d633e5b5fee2aaa20a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8a20a2da062a0469cb7bf2b3bd96ec6b339bd1d96bbe5374b5ddfa65991a21b7f07c562fb31a9c030880b6f3450f37f5e3bafe0b5232cb4558afb5d3157d1ca6f7df02f9f243f9a9cc4ea547d4bb5e1bd352a4b06bd65b2c8a961b11d32af1878ba03ff0ebeca2347e71b23f66d2922c01236aee15abd0b169c91d3de1310c742d6ece78e67b23567a09c0bba20e82f7a54f656eb9ada8895a9354d0613b73fa08962a2cd14f203f1f330d6512c84590d0d43c649d4ce066ddc142986971023bfb0d2f8c43ff20c1e98700902f07a2451d46f30dbebf0eac1ce07fa2cad86ae363e0b1cde5120917c0c742048bf9c78b07ef92ea7b578577de613ee5b0c9a18f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4ba4d35903c3114f78b47c5a1496e06f927af7efcc01424ce5d5664ed95b640c8c0fef94f9197f0c6f8102eb5613421a2df644bce8883ce7f6320e0615f6f265adae637ea64820d7440866bad76fbcedc7333f2df13960269d787c79d04628cda64d72e9a48adc159d1d8413a483eee332e51ea59e11e9114197588b86d9a50a197a9ed4d32ae855d19f34a532ac91b2a73b1f9179d7d361e807363c15136e86c3ff0215df49fb7cd77ed5a25c7ebde45c2a2db6c1efd9b3e8a52ec57121f3dc5d20cdbd4511a2341c2f92155ad003ec6764977167739a3c8b85daf2c5feed96a4683e4ff646f6fc0688220e49724c6b91528598b8c000598a76040170b7de8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6c85783f2b4f7814591fee04da570a2140aaa76cb547885d352e2d04585ed2dec8986a49eda80ae7d69129b6d975532c85659544b808c84d151e15001481b5fd8e29d5fe6f5820f3803bd1479a2a95783035303f60a9a0a5641be416e15aa2eab1b349c633d80c5977478fb830cee4a02231106a3504f98a7bd50948eb165eb54325ba776b149241d96bccced127a437ff6676e7eb1072240573de5d04b642b5416f59c787127fcadce1b6a8e9f57aaa1b5bd87a2c1f9521438bb3f5fad6916001c1294a28802f7aacee4363c241e7cb54542fefc893ae46b511e855dc8278241d3daf0dc9aece2a9f99e16bf6b4a6af602b2078dd3af2a0523ccd298e18c167;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h395945a2f1a4f5a45bb124697c875e38ef69e414670e743c680e966d8cacd97a42a6170bcd4bdc79d543b5709d42b638164bd1858091db4b0e240df0d8957fc84b97f0e1dd4f883ce0b7216754195fc9ead736157a7fa9e96a0657753b9d5227c023f040af69b2cbc8508721b82d04bfc176f7be6cc07e08269dfb1d722eba596048294a3c35e8d6737f38e2971ab7c862dbb52213a599b920c41c3b5fd7bbf7b00d2759e992cbfd7a8121fca1b29aeb912c3b4bd9f3fa32416b7a379db0198641066061f3706da2bea757bf29f68762892b7b848c4023b57383decd3bd13dcd943b413c7f094398ff3248a2c07cb073cbd258aa35739dd62ddfce7d21b531d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h909f5abfcdfb7c1f5a712a4bc449069a48ea5f59ce82d75a36ca686d0c91ccd926df599b5bda8ba396a4a8633d05990a04586eaee4048735d5830f586ea0c1eaadf8f8451f78e5ee75b6e03bf02bf396b65ec14020aa519f9ccb7b2bc429448becd3c62c112d95c6cf179f096964b1bc821970ff8bf2a158e444c2e6515717b2dd4faba66c41a8b9dca9445fb29b006d7054a330df42a00504cb7ed784a688132603a32e12541320b36b4037436eae72568cd384b3c887e7d6214e9aa837c3baedcef20f6ab7bd9714cafedd976438c71e502a0ba2eb937a4f4cd2f6147f158567ed48cd40269d1580fb91e7801a3d084b1f02249c4af6dc521d1c360088d02a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd59cb805230737c0beae3fd29ba3f299c577c494040e210be827cb22325cae4f2bc5c35ffae6af9ad1c12702e61fcbd689de690672e3653471e2cc7213a81f08a98f97c7238c95be08f796b825347df2e2cdf5276f9194bb03c06f15d837752c798b56e7416ac79e5fd9968261560eceec77f6122bab4572d49b9c2f5443dc808e79bf3b632269e77eabf242b6c1dd26fbe9576588894dbb41e0af236497cfe042a39450a852d42ac6d097dae5e1f262238078c6d76d535f3c0f6cd1dac9999a78a789386b589c195fd63fda1ad0351955c07041537064a5822e4e0732b05f5f2cbd4c8470e394c62b574b0134fce415a46b77bf0acbbdd75bafa4f6c09a50c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2d98337752731eb9c2c94da7cfa938438bf4655d6aa00462af8af010e568b97c4240d1da4d20c0d84f993a9c2eeefcffdf62bb42af7c6ad67bbde69ab9bb22c40f6c5921b132b06bb6c32814a776e2d71b637607124e7613552e60b3aea6c42ff3d66bd0779370868ca3ea13b6abe33ef089ed2f5172d600164270f952e10775dc6e3bf63e543e21c38da6966d9110f9f583355b3f6d9ebc24e30f55514ae20eb5b83dd262f267abaad31523d36f6afc45cf0ec711565b21d14b17e745bb9b6c6d55f35df46baec431ec75bb7ffe997028ac1d43beadbd1ad11f77b4657cc8785e94f548cb9e00c854f51a30fb0781a53d354dd4a8542eaa41f7e8360922aee5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb650038c48adac261fca2413fb6b0843e445e15bd768cc7f28f26f09fc89dafab85daaf70603da557a1159047c8633d7d2be6e8d2c7c1034112aee02adb187762246acb11c6cb0e650b2a6a2148b66adee5c542e5b75f2dff905f47ab64ac0093c293a849691419ca995398018674c48cdaa22a654f7e6360339d851f9b97c12f967ac63e25af397cb461247853eaa60c24c75fe49706d2cdd7280c4c3bddceab5b78aaa585c914ac485b28e433ba3b94f138aa9b1a62b1a2fd8a5e0d1eaadfde1b8ba0375d67a37980dad76d9e71845a29640bdc278f3cd544974442d9948b31f1c5a17451c0a1356b37569ba7e4f2a9d548f60f82559bbcf60edf2657341d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3208b31f2172aa957422bf44d95c320cf84f859524ceb65cd52789b5d22b9ed3cde78ec56fd1e4f42489d0b45f65bf738713814396202c630b88276bc564636289aaa54195ef0ba23fb2aa34609bd064c4ac97a9f425f15ba03f56977f4a134388b233e8bba57b244ace2dbea386b192977b4f20effa0c9b12998be33460fad7fcccecb2cd1ce3f8055ef5edaa724e7b261745b4fda568251e89da633a5232ae9479a0e5c0160e030440a80ec56118dcdb815d2a62fc87483b3c4beb4c38d3b515e5b0360365dffad08f3a5d7bb95f65ae5cb091dffb5b57637e17ff0a2019289750aba9cbc21c8726948f80af05d182e8f15ca111ca97348031ab25b517dabb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcdeee29b4701e675184c5ec61f39cfbb955abe1924f88aaaecc0c6250ba513dc0650492f24a8c764f1c01c1f53e426e7e36d5f7b12ceca1b7b97d5562cd8225178c31cabe6efa78276a2defa059d2d1ad146079264b7fa3bae509ef3c24e3f41331e237322f0c08ff0416682d2f0656549ea7a2c72860c39fecd12d269cd9325f2ef1644c03c5b0b919fff0687f45a02f3e82a324c76cb27495cf3d33804e785c5ccdc24fdcb065ef4ad938f9445d543827f3787efdb7f9f749331902ad4b67e340613749095eeb73960a53cd153f691c8b74b400102270a91a51aafd04aac2707312f9bf8d6bf7ff5a90cd329aade9d6ea0d5e7527d8ba713d22a3402ba293e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h133965497077496bb781b1ba07ff298233be9561f6a11a7f3734e0659547f2bb4c0d578a969c76af5734fbffdf2ac2a30c3e45fbcb7dff3a13be442bf41a72f4e4d12d2abe2cd8db49b6998232e03754b79d003d036586cfffe939d93b8d22994d370c80e4c388b8bcdd8c7e99f6cdd589c5f46be98ca02ce8c19015e11b82bd6bce8537b67d86a3fe9709c9af45fb460cbca1d5efbc37cc3860ae77551cee8040331fb6a2db582b73613330ef2c51e4af46c4ca1f9e6e7e478aa9a1785495c90518b1ac993af2dba9c8a7afe6f344a0fee8bc57e0b400344c4a78c950c5e8cc851362c8124b3459747325fdd578c8c88d62cce73b9b7ee883f2ecafe3a3b790;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he47eb8c2950027df80e58f9a82612f29dd085fc0a57defabf257824f4994d6fb01844a2ee41103a618f65352760167fe3895d2a02e94690fd5c1b9aa79e81f077ca9932042ad05a965b5096afe61c579c56ffd10aae64931f9d14c2cbf4f91a0ef433ef024142edede085b232b3b42137b467e3cee9eea068bb406e46ea5d83af0a5b0a768c9d1cc39aa6926e34f8e4f0428be44550db94c5e19bc54281cec0a4f39958a9efbb437d9f20ac9ac3f3cc0405a440dfa4288075b354174be41983b38c30b7e5de2ef78883767941c0920153b578682b93bdba3e37986bd4767128eccb21818e04e4c8b66797623c59cd0ae26ee40cd49457a78df34115b1e2931d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2864ed7eef26e2aa224524a9f3104192b86f805a6011948093b34a5bb525d97fe7b6d43bfbbbc1fae179af8c777858095d450cbc60e64eab787045a6090e0bfcfdfe75a1e9c8a7a2a537c3e3d6a8ed0f51bb23227cd3273872abc18ecdfcfd42ae90ad44a6970e0b9d9e531f48ce099b61ab9c32651e22ddb47d10a60bed790158ac8a60c187291ba60f24d1fcabe23857d2c3e774d19c93d5d5714674f3200417e3a369634c7d7d339aa585708fe1132c7fb2fce27415ab3c8a5967eee1c7757ee65c39fc3980b4122609d153ed2469c142c1f897bb73c92779b1c4ca4cb0ab7cd84b82a2ab9a362635e4d0d435c60f3c5bf6570c86b1da71da0d0bc9ad3ca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea0b657219730098090b567209ef635ff7e60c570aff6a86051d0d430be2ea8c27c9b92bfc9ba4ff36ddbd6a981fffff779804da56bda2f558454b32ce1524cf8c27769ca8c930701dd62a805f1c1007fc59854ecc6f60afc4ba22508f642b1c98126752c7d060a1e28dd3bedd741a72dd6213b05dfe6352173a8522bfa7734f67ca4b561d7a65fdb8a3cddbf71ef4f3dabb869f2c0beacbff0ad0aa6917751c42715d7e7f680711c4ef0e44834c8ba03950f7066a4735b13bbc4dad92580ec4671b3f5b27181e80b8a63923a1c294dc4d8a122567047e0591db77879e1c0869fe2be30b0934b18ff3eae44f6be18a908de80e38212d3e7b17c12aab0831ac5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h51112ffce63d2aba8d19c9a155aab5f742352cec7e9dbf0499fee633cb6251afa0304efefbdaa824ecc80c013c118c65c191960fef21b097e72db8fcffc5b90cd3e5d07f0c60251ec435438232d0a1037064063b8da3f203169de940049db7c45094cb3350c1e671ced0a309c5f4d93ed46e812229054730f6ca86220a8d0934c42ff649467cf2df8ce5ae1802ae0eb02a6cb55ccccab516c9c6e7866ab2d88d76b30fa2165618d896c1533c3e17268c598bdcb2ae5a6fb8b3b0947265cee0fdd1e46abafe87cdf376980f315cdcb03e391793b479cca12aab7eddfe450b4df7cce10b8689bfe40f9039dec95dda506fea9717713d79948bbfa89cc3dd1013e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf665b3f794d47e70bf9abebb109ef10949f82d60d01062d0367f9828c4050889327228b470140836ccc669d0de6fdd3316251e48fee76ca4afae72fbc15281fe4a1cf999addf10ee2e8380ca8a58e04aa7684d01de878d29e11da5750b83799a744fbf037f20146223581d27494af1a0b5ce62a8da97bd746161d05f016ce7bb780a69b4e4daacb293904f4ca4a91a26c33e0d758949fbaa49a8acf735c3298b57028129cabd79cffad1bdec42e178c51c179943923c720fc0841bbec30f05ce2373763dc5ea92162b8253d7f2b8d4a57dc2928364393654d88062cc54c4f10a8b42c3f7677637897ab19d9855bda48cb4c46260526a9093deccbb7bffb0829e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf66ad6c723e06a5dc02517c72e17ae48f79a6a4e617a3768b1c3134b2544b71548c6bcc3bf4f617798add52f4177b066160c126b1b493cd1f5272b55882d7e2473f2e2181fa3112eb273dd1ea86c044828c3962d6a844f11518c878c517d477f8698104ea5fb202e70f34f0d626e20f07e1439cdb69433bfc15fa8d3d2049c3b1a2891713fc5e6b1b46dbcfc7705561d867027207635f8736e0c5df9ebe13bf86172212123b2f3c87bb90e8cbb35fd5e42cfcceb4b2023a7c3db8847aa2b57310fd4425869d9993f2d335023801985b55c0d19272c987666edfc0d78cfbadf840cd7114a5268cebc5cff5c9256458e9877d06b03cc043b072910ce23b359ab3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha658ff49146a17917e2da60134c362f1246027b827b70a326e49abc2bab081955cac645e06420cace5eebc4da3a23c953ab876640efa763cbd47206c3c0399bbff2a739319845166dec3e3549c3bd149b4c95a5f64ef16c56520349fc1fb9d58c13232e92b2eab32fe6e5cc276585d76ddbd5a4cfb53b539b033dcf353b484d8f60be8e925812c0cd05eb4576d2753aaeef4f2a4cf4ea16258376113eadb31c956c7c9749cd985efae31e627757a70ab103ba8c7241e661268f520dd8995413fd385a1deb8416147ec7742efa79a5086ab293fb9183abdc8c04529e72c9cdd04b928e44e0150f6594e1df5322d33705ae5ed49a6aba41ce6d56d40e81c570431;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h74e69ddb5ff141398b67ac69e5aa191a0b5dfdd88c9b429ebfa7849649bb5cc0ebe660181561b96c2492d203e103bbafa8386948f04418e23f7fb1b38d5b7cdff05d6681e8a7c9a151407636d83173413f10a0f42b09f001e9a04fea11d2589fb0ab53bc76fedc730b2e46bf5af52a1cf07ff8ec12b27d6fca16efcbffd634eb3884e0f2f0078ccb08c4cbf2661b9c3c7be45e06ad4a473b47d032d6d2b99b52e3b0cdf8285b099ab7fd44328e676ab4de7917375939710510c5b21c7c6445a5e881da4e8d77b0269c192a2f553d81fc6a3e9f7e7fc99070b932f0a3b0984d6b1b5c5d3d871a64dbef2e95680a59f0a079f6b0b91a822bdda1ad5df4f9812d09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6959d22dd79df33273b4126e22f9e8b17e59591926da0bf4edf8677cde418cd35cc273cecfe6dbee95815d5db938af3d147364a2e5a636d2c4bcdc7bdc7caee57a17d6d656199f84873b866ed99ce138d69fe1f81e0c80b1ff7f046fadeea769f21ec2e0f066ad341438dcce1224017275695e1d108c9c537e9d1c341ac06797371b7030cc1593936f07f533fc167573975f8aa25b6a48fd9efd8542184c098686c60667dcf1793c80dc4a08b3cfc674c37c497941aefc4d3715e99d2abb84b4708b23903ae45aedc5e2a7360965b690651c3d64126f6197738dccefa6f58329a73420f2aaef5889bee2d73431b294c36fc73812ab45b93070d6b43d2e9ac4a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1dad5cd96176efadefb4b9ece0e82b8ed2c3d1d87520e828a8c2d91f23a6588d6e94084b7dba5291e4eab551f738e36648313920829cf37bf1d416412a1e3e471a574b27b1dcfb75863e5f2797cd75940f1495584d501193c155700af81bad98fc5080ee3ef54f577e26d8cb3c753848bad8ca7fd2f9cb39df96cd35204e52f0f59e82056235f4249f2ed2d2a51198a0f01b9f6ba02a3d6c4dd6bc260be4e89e05656bc446c917e66b43ea8651b9e7d848819b2111a0803e84c52e60f5ca057e719a96292a4433b794bae59a5c4cc3bd2a5409f66c8e1e057bdae929b9bb37ec03600e51d6291956880893701f01d6074259d9ab775605da3bc72155ec45b340;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4d2c0765f30a4fe4e809f8f991cdbd6c12db737fa405b9583a06058a1d18772a453e957af4313f299dddd8b475aa0e64e4e252947fdcdaa3a2463a965058d901a24fe80c7702e0cc980110609c684f81c65cd57c698e909c48848aef2d02fd15987d4bd1403cb67a9a152cb57d0ae7073287b61416aeb2cad3e5ff04499b33260582f6051ce9be375185f1716f39a12f8c36230ffe88ae6b5ae9b707adc84f94df2f973be865dd788bb5b38738694e8ac2c7cb6d67e8bde79822e3d13413c89f18e10d854b532c56c6caf9a26d04619c4f1eca9eaa927bf55da5a80a5c51ecef4c82c74b722accb32129bd875b4a0b6e03c2456498eb4c790867f6b41f36b8fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h52ba8b2a117b38d1979f43923239ec57471624f62dfba19d3fb67c78b427dc42c7416fc9694a9c5c3654580bdd703072ae5d5eba95f8fa9caf8788485bf46642ca9c1ec567493bd5937ad60654025af916c41878190e248334793ef8174637efa94fc7f1da0e5f2211d2f73fad196011ebcfab72ff5c0a2ee72fbd18b9909030ef2a2b708afcf016dbb70912a518be93dff65b68e8a1dd40691aeb025efb28164481d0a39d116ebd5c237019873c1562ec252547067409615e6595c3137d739fdac1ade3bbcd205aa736cf67279c1eaad7d42d5233713322847f71c280a97fdcf1a473d49830f5a529c64c6eea627ebe322fdcf208f26bf625158c555168e805;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1a698694a27de286b59e12293fb4a7230caf9a431f631c9701ddee111fabc9480d772b328119799aa9e3c7232c23c4ece2c11d7699f383faac5f21aff992505c31c1e248cfc0e3c2e11347df048c447e7ffef8556e76e9f7790a74ef17cb0a0c6a5e7b70bcf06e5a91ec5229d61297acec66f4376daec9f9aadc7046d54c45cffd7669ac4fc5f9cc1f5c046133c00a009f64561f82181e85098bb72e4192e8d07f808e9fc9364c144cd529a1d6d7571ad954e0260b31f6ce8e7c3bfde1997d6ea1b41a73024911c1228576d224ffeda90b055ffbf6e2631aab1216fd70c11e141a9b8fde9c3d5ec08cfb6891808c85e980cac3b9d761bad974350255ff81ec7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6ea79294a0a5690b63196d4aaca8ef7c5e15f33f7d6b4536487d6f891e5f37e30979794bc428c8cbf7beac99a8c286ec27945a6c22d86076d6d602259102e0e6a918d2b230246838b627d5712a1008201bc7e6d49dbc4e25dc5759e8ece0995a2c377eb79f4728ec271d4e8b02eb3041a8f70bf3842a37ead4f7fde749a754ad81c1dafcaa50e029bb7058a1003d9584041e7062c96f2af0b8a7d242e5797bf414efc3a0286816f3535c57f16638aa67589395f57d42adf19ebf4936a874005d3973e7c708f0d008383e9211d5215d9fa1aaa699c395c775ef4bc618c3076e5cb655285289d2985b45ee5b5f16610ce508579441879b9b68ff4ee07ddfc411d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3a0f9024f68617ff7421305e9639e6f3d28ff71da44f65a43f4921032fe3149dca3f63288e50e2d3de57c59620a93f02f9dd2311b61cf5b3b58133885f4db293df95589b8bc4a23cd3b44892633d51365a5fb4e352b873046cb3823e0d4d407500154c5cb2d68033eb8750d38fb221305affa798db56faed7699e5516bea27f66a82db82ba5d1205fa994fa33852c641a18d1cc2d30ff106dc73e32148fdeea7a983550967056f6e1ea7aa5e9aed4db35e603f12f42b9aefe4b68ff58dee6bc122887a147fa96dbeb82757c9b6175c257b59219640dce08ea22861d5aedd61c57024ef270e3329b6ea144d3b2ee82983c45a33e673f9eedbca4d2ed8565e5f50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcffffad365e8dfadd292fac30f50cae589a38747b5d5f4c4ce12b071f4c285eb2d9c2c7ab3ff103ec9d53cc8de2586b0212cc5f88e15ed87621b42aeac22325f7ae1ba9af8bc77bad99d6bc95484646d3c4eb86323f139e1d57426fc07f04f1c7daa24ccc4f561aa82a81685180c58b8787214871f0e50ac55dacc42a1aeceac2765016cdec1a715d6bb4f83210d28966fa8217e00bdd6aac82ec89b8eb364f9173acb824ce03d57ba8f717e4bdca18e1f28fbf3a148f5484bb237c377cbda48d85622392009cd42554b096755d46a1ee79e4f89b3c07c22e8b60c735c396f7baf7f8ec04f3f5a32e133d3e18ffb40c38a854863844296492f004dfdbd88432e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha66280a54b120cf537ac7153689ddd0a4c7dd6fb02cec06c32162fbb09770d26947c78b1f76ac9aeb6c76d2dbb1b4adf0c2d1dcd61bc6657ba31a975fb7e5ad4bd0b2e123cca124891bd7b519d10889a87d739980449081a1d9c82852d44a977321d8decc040dfb13a88076d3be4dff5e664918fb0d13cedb7f591d15f96392ae198cee31b4171954531fc92904e46f5059f967fe67efb5cc5681faae73ff716da854c9d6b78d62036c166e72067a93a08c03217888685385acfc0c1eb092da54b439546dc5af722833602124d7312ecb56c6bf321cfa5273dec84fd976820587863459f9c024a4459afcf5c7885032786e23e7f590e7599498b549d5051a579;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h82d58ccb71a19588e592f12cba8364093d2d30bf4f126e644208c315fba18aeddc9d424bc5d5a56db0ba292424d1bd271d031d3a0968257a6c606f59502a10952d14547a07da5914604281a6046326e9136dd000d140881af31b9f745dc024c2d439dc2ce018288cc84ef2dbb9dcb8934b7f83f66611215ee7212ccc0a1710654d99fdd27cf49884494ba9520b5621d4f9ee8236b487d1297b89b1b81ee9941f5b9b1a6ed6cca6509b6725e3cd83cfbf3188dcc242c98718153ec2f396b203a534242c1772fb59eb33de7f20bcdcf731bb14adaf36f8f17281c62601c50305075f1eb52b5cd2af42bb8f66a7c29e09a9e4aebc2792173e90d2416996dee402dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h671325427300a5ac45e5c7734cc49b07550edb5c8be46f57801ba44d29e0e8fd46da099f7ed169ebd769ea9d35478ff4b65c3c744aed5ad76c30a2a9e7df2ca2044b87a26b43c3ccb8b369627c20ff08ef077ab304d942050ca29cc7949e1e54766b894ab63d30a292dc9a6b13c5efa873152953b9e28efea5611dbcfeda4d633c9ba61c78cdcc0052884239678b3f485d4422dbd39926eba9092220b0098aaf6d0f23f194abc0fabaa0dc9ccc3375201155fa696ba8d64bb8a04a4f38f40417f5a06b4922e5a1df1bd73f184d8e459d3974762d676e2946ba8e6280294b126c80585a61a2593bd585010e2d51c2fa2d147fbde9936bec735b0ec2e8823071f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9fb8bef35b05b842c2e18f1317ecbf2956fe2678ab69505aa62e5cb2c76d7414e05271ff85f04b9612ea35c7bd1f0704838007024ecb90d38635b4d5373708fa4f57f4cdfb646ad4558866aa10b26b6c30879de730493bb1c4539895174c16bf1fc056ea6e114d6272a12e6023d397ed416b2af4c0198653c5a00301cdd9aecc21c535dd70cd9ae2529d4b9f5474037141a11180667e5ec71f3b42ba9cb2fd851ed5d1d7cb847e4c01f4ff006d0c5138d11b864e97b12f2a84dada5d65a8ad839383ffe3fb66351445edb95cd5702f24890aab639b96c017aa2fe3396935d800388f5110c78a6b7eacb01b3399d41201fba837d929d27649a530f38a0d5b9934;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h200afdd286295c72a5259477793b24a5f10d706e57bd577571bb2c0fb0a2c32063fec87b0a8f704cd2b298eabdd79942b70ece9d566857ad50129cab3001c5435dd281a1d103adc3cf82e6daeb212f28c200aaee94c1114b2cf5836d127a3593f8f1cd0b198348f6b848938f1b989f042b96a0345b703412b929291d58e4e2454cb2058cfc9f1f1b8da7d2a881a955e7d199327030cb4833f055102e884c5908c00fe04e9fd24f8001170f714eeec32457b92388b9f9f8cad6be1465fd24541dcf3adb55f14e2e3a890e3166fd950c7831b894acdf9d910b7736a82ab27db2fd1f47bb9c3931bb06653366c285491694c633ce8ec6c3907038492bbec98a3ecc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he82db72c7c4002022020845b62d3b7c24f15a32605c0603d03a3797b2a74bee94f7320c508bc78127c17cf3c8e5f65c54f77f99b002423cb073186e3d396539e8334fd04a3b792c94f15018a5db758adef9b1c71fa7a425af10de057d5606b776f27ce9c876a511e5fd4c0421b3c131b79ee0aecd5d0de18473dff5b5dfabd25344b006a8f1e07d95126f7706bd15b9497714db6286d6762dd98122ceda5f69ceff911e647c30bcc5b0a14a8816fbbd0aebfab23372b1e8897d4b7a584cae7dddf9c48c35d383a18cba340769db4232addcbfc117cad0ce63d9f8d5b1250319ca9c16e70ac94d8c4a5d69018feb6ce6faa568ed2140875f6112dea67dd9f2c56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha12327e92521ac6b35ae3ad66934d6ff418615f5f9641cd66cadb1d217bdfc13f2ab36cc1349dda14c57d6810b8a2c9f58a1c99fc482b929cee327128646f859cf323741d9ef6712becee2ed971ba42ecb381aa12199881feb4d3e50138444fc39c194a9a07aaff62ed00ca1112c3e0f18ba9404d2b42f2bd99e3d601d1358034309ea4996b9c11771e7523543d7dd0759ed80d9a558862ceb8f9c933d43200ca110e4a3f1d486bdbd3ec2a7e5e7eac140eef776816526d38b94bc07d7c13fd9233e33886ab1301a5626bb9387218ced8ef945db313a818d831f0f0dfe233c7f54dc1c00c4336f5212b3459ce8dab5c32edfed2303fefdcebc85573e4b7e49f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7035e7b2f60d724106796742f2482397c8a8c4b47ed36874b96ea7d05885e0607e59f1501cc54c4a3ca9d37af9a3a3f6a7a8a67197549709366a2f72b0cedd47ba4a8bacba12b4cec8bb79474cd0e3c57f8d4ce23dbeed9c7261dc932a174119cc9e910f4701dff5cf72e5c20faa13435a317f24b42e7b183566b76584cb23c46c6e520254493d1f175f05bfbec6e911d71177993dc641cf1ad13960227c271e3bd04a3ec72ffb761b3320550cee29f79a94a156b92103d8e2aac0a384b4c9bea6663d08cb37f53e73762ccd0b6731ef2b166cfbffdea8bf75c2c9acd1251ac807ac30356f482279f33d424420e442782c26f4943682b0078616549f1d447613;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfd6b09f41f6ded0d82b06074d14f3616f7e825e3bd6deae7150cc59a686c7a58a4645ec0e75e0e9e2944b26d58bb18ceea1d9280bb9d2525f4eab8d67c52609b7c56d9a948b46e0163090e3110e85a5531a5874f4fb71f4ba5bd29af45b23d80bf9a722e748c09e0ffbd17a0ed76d50c7b664f11267bb73575898bffed432ee1fc9527b806a36aacdb5916e1cbbeda4c7ec03c37efc14d3a03555864a1438b8047f93190f535515c7a496bce71ebd7c0635a7b5c71b4b209b8a8a6afc52d77ff15b7ebcb02a38db953bae13992e762dbb966e8157d777ae924cbcb118f7da985582f236e6920ec87980d45ab4cc9b0ec9692dd57c49fb0992e724a8cc1febe43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7382320eadda1f8b7409a1b818d04ac09a3690b1c10bc66a99efc65219ae7bf6bcd1ec4f95abc5ee42259cb78521f7b702f6b386cbd85d11b60fb8944932b356639509a6df44301bdf0db34bf77622a7e9a4f483f9f192cb494e9adcae974645d6ad3a79657970fd3bb5898cf8775d26fad26b2675b50fe34abec18568438224f95a6ccc13a322206a57c487461a3e695915a88685012606c732b6f11a87e9be65882f6911921468fc1ad15c74acc30a13d85e202ddb1c625f4aa49f6db56c5ed4ceec020c0dce2c00aaef8f2c9f15172214998a4c39b874bdb0d9d858e00a183dcc23b8871c0c1251e25f8e6678504c171e05f220e080913a9f6fb34b391e47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h370841b50f2519f4851d5245e80f86eee4aadfb762f9f86fd237d96799ebe37a3bdd6ea9a56d688c57b9832854a915eedca2e5fcc62f58775b1507f763ed8a3fa2b66c8b5b1f31351fbc2c0a68cb05e8ce19c4b104651feb19156138e53a80be61616e2558f47e0ac10f0700b85a1c27d3388666565faec4bd9b1fc5b8efec2d5e5117e7a845188a830b95c17a00ebc0468d18674b9023128659fdc028779d66ff55260c5a587738539d3dce741d923f035e06dc306e8c0f075a038c93c09c10ac55a33aefcc7d787e1cc84acbeb6f5eced3173a08d1aa148bf3572086fbe8a4f5be3ccc98b14dbdd03383cc28f4a590f83fa3284bb2f158160f583de11808bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'had97b4aac42b11d2b0d1fd8cf76a57cb6b9a6cf5f47740b13a72f98e0f7279ad57bc6849b3abb6d0764f20a8a3319498160c0104d2385e0da57e6215d847f0e6372fe4655931d4a14aee77a851fbc91fb5946afc84bd589001e1c423fbe3db0f327049cbcba5237f7ce141769ae1478cb3066f579c137b2d45c363c2d84ece98a589bde88c756b6f4ad016a093e5445131b4bcb49f5fee2beeff70210b3a3960925c8df96158517c2620b8accbe66e69b9dda65f047d0e3f4cc4cbbc2b44076abaeed1c65eee9358e9bbdd52b1535ea5da64e31912ca484350180ae09a279d20167666ed20752e7e5464c1d5ac2189cef2fa6e803a80f1759ebcd7ac37897c66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2acf4266cfa817f4bd185b6d45934517c9503e554a5abd06906d8c06a915384fc0b09852420d866e95732d426f696de00cac61d6c7b3b768646b276dbd64735d021ac5cfe147b0a4261c13df6ccc3a0f59c75fd50741b5b4b0be974a27324257e5418fe73c090325c6d9618cd711d80188104afeba030d4cbb3e86d566ab950fcbd8f57a7766b021683f26e0e49e0a6aa05707f3134407a159d4488659e5c56d3c943de4a3df4db7c0393d10d566a677fd526f8e1c24ea0ab0ef9b80475d8199e0f7ecb1704ee7e99069931e0984ce74121f2e0d865031bce33f406ea4374eebf50092a9c3d7adde6e39d9f81cd7ff33da8f122e0116520c6f039cdbefc2573b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h281b3ac13f68787a97f3ad6cb4ff729b8002ee9d8bb2ac497f0d83b60aaf8c461edc1d2b3a7e53bebdfa2097893401d6ee907603634fe1a3f978060790f7d94865a1789da6e71fef11897f6abbc8894f96de5e96e68291db8ce336c518bd484bf714cd3f86619460163969d009c632b10206f5b2127b19e10aa6e1e7f5a303abcb261d3c1ddbca9cffd62f8a5dbab1fb95c1d2014b7238fadb0ac28e31d54e2eb134ee3563b7f24dbc38e9b640605468d83c4be6d9ca84aec63608827e179675dc5f974f1a79ab950a2cac70a4dd7691db80fc26dba42c96d388f797488f4b7fe30ad441d2804febc8531e3ea11a8abeef848e6ef0800d82a3ecf5008854fecc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hce572fc2c625cc667dff20b663cae3faf862409d70b5c90c28b382b694148cea65f9d11dc097ea1a75a32366650751d8f76f81e602954d533b2c060f37d79eede248bd963c08b4b98c44d221711e5b6cdba2d2be68f59af372eb5d3d946d20a4008ab1341d6924d7762d469425d9b075af013e118b56ea76bef7e0397794b732a284fbe5f787865a74fe8e9b4fc89c58069d1c7d7d5dad029629a6b51f5b9021cddf89b3f6727fb463bdbed82a662762c0b5ef1da8281aff15ba10ada6417b0fc99021083137a01117d6e9eebd0cf74b7736402555577d93f613fbc0915601f5a38867a8e3fb3c0496c5d99554f4333beb2b5d2ebb20b9e97b822424a7ab06c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9e83e1e24ce1dcd40cb39dbf1b36e57279a41221769f70f3dbed79d0ad6f733c38aed9e9c2be389ae1fa49fe724ebe904fdd7259d8aa76ae4b880de1349a6581feef1a24bf39c34fc7e665133e667c60430d164d6d89460eb42c1a999796ffa68b29e0086a8912d3ceda741be78af40cadc79ad874a3f5331d26fc4653e944bdaecda445bdc5e63bf09f06389fb91fdf582f106cf8d4af7f8fadcea3d4fc5b962a9e22b32e889407c5ca9174d9e21a200881727e0f8978691c01aa02758b57dbbc33f9e07e5283bbf9f4812827c17a90b730690b6646300d1c229237790e70b389d7ea98d1cc170024722d4faea3cc5beb64132a19eb15efb8a5c88fa9578c36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h206ce2ee4fb8686bd616d8505564938b4f444b308e8ff92feeaa50c9531e2ea6aaf542aa8e70d03fddce8b0dc5d931f04c60efb8c0d85a41e5a7b40aaa146ce4b95c84cdeadc5e544fc60f846fd3cd9733644380cf7e7249b7f94a39b29ae8ecc7232ab66aecc846f068f5f42151a362abc1fe04110ffcfa3ecb79ec437bcca9f7e8b7001c2883fd9f6f7eea4e7ceac534fe2c486498b0c1b890d596227c0ef2872e5db78ac432a02350ab56403de4f58e3771ab3b7a59bf91ec978231282bb9569f868d66d62b8ce30687cc9d64bfcccdbf0d07a4e4a59c03aaf3976ac955eaafbe5aa1da6a08281319afa51449ab97af84895d10569bd24602216353db7662;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8912e164c35a324b8cdb0deac9f32bf3285d149b19ae73408691389f903d4f32d28c1c5c04efc6c4e41654f9665ad50ca6fe6c7818e9246dae9e74fd5f4a48151636c407f477e2f385f97f76732de72d942a399f53796e7abf818322b9438a1945705c042b61ccc66eaca33b0fcaeec20a2150e2540be7910acf41dfce28076595e65842693a2f76eaa2fe3bba754d095a1466a30ff350004c612b41f149c923fc7ec7c0e89b10c196f57b3b771781ff8e67da78c59c7804d0dcbf6494f2baa603250093ada40c0115eb828084b7e4735a4ac39766d969deaeda5ebab454d9975cebeb4f7e83fd45bd257dd06171c0026f3a9d1c0cf98768c2f38eadf1ea408d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1ffa6bdfc27cbf8f6e4bbbf3405978d5ed49a625a911001431ba89a973e0a06604f2143e0716fb23e2c48d081b4e7ebbed44de651ff6ab5c8584e115b42ff0bcc93c8e9e6b7b48d31928bc3e9cc192d5177e646ad71be7413a255200fdb8338bb81e5d471e3a34f35dc4650a6fbe8832d1582cec7802e8ae6e374e3446ecba8e47ad39ce0d20717fee85322a9f17b9f4722298fe1182af61e189ec116780e906d8853479a28e7ca6b8bf93c07aeeadf96d4f2377d258cb0f2fa3e5de4f2a28b21fce4a1172c31ebb3ddc1b593d7f2baa3d6a6e4342a741cf1a115f22ff2ddd2ad9c11007036ec55827de8eac3c4fca8ac5939a7702cdadda2cba821d359869ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc7a0d7bd8262edf6c904bcdc1c29bf2a3dcc8fe670f83e82828b3b1e6ab9b1f324fc3cbfa4ae5d010731694da6156ab9de0df5d5c1505db2915da25abf501b7cf2740f00381bffafc83ec7f17773a5b107ebb70f52d1113dda46044689f452015852b40d9a6bc84bad34a4f31a737df1dfa9bec5994904e1114fbbe295c9b63e12bdfe5b35585ef1f7edef0f3eb2a9bbd1598b8530b518021dc7b46c5f7e4d52d9f61423995dd6dd9271ecc1b36161353777b3823dfd1d81b04fd300ae301aa0ed01440235d3cd2d2c830d3aaaf8886bc266f6ae6e9ae94aaf07a219ef8755a01c6c314f6ea0920ac4e3bea1078dc410f97ac3b8587997a001f5fb1ba7dfca8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2cacf116dc043063a1c3335d3aa27ec36b1c6c733d573ef8348e81225e030877e0bd76a6ab9424f1258019085e3c4ed4b67d02c97a7c5f910b8912974ac038f6f3a9ffdccf2daad49ac2e5ed20c044d4bf3a0747cdd26080985f10b1f64697b5b8ab6af5eb59715803f71dfac5ac9ca2490a466fab725d81e41bb5895c4fc0581256af31203e063a5b6a82d20c9e0e49c51a713dc4c6ceb6ea374032475c5fd6ad0d33fd675dd50e1295b4947cce04843dd387ee9bace4811ea8eb6e94e6ffb85db1535540afb194bba4110482a1da352ccb209ce187995487b0b5d6b830bdadd30550ee40bbaec86047911f77d0e9afdac215a3097dacce94c6fba3e4cc549b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd5e670899d804436b3d9e151d70a690f0c7cb399d4dfd32013d801f6b1ae3450218252adbd603b960b4ad530d45cf07f03057a63cd60b65a15f7044fdb6bac802f9c53da337d6d0eb7e34dc147be3818d6c3382cdaacb072a4b4dcc26d4bb51a7c102c4555fe5fb434b32c5d0be82a022209ffc1f141ba9c83d9bfcfc61d9aa46962904cdf08d63874364357831790201370d7918bdb599b643d1a470ec04e1eddd82a02f00a20e44e910cfe2b4a9321514b03109d109cc502ff88292661bb21c21e51dac8c2ab1ce22a4514381852a6b29e7f82406615e03546377eb88bbad1df1775693e67aeb14a1d46d0ba9caf5f197a8c46ed29cfabc1d3d517287afb04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf40a046586ee0c074ae16e56a57e5153e190dd8a471839d05fd40c640e53a8f0d9eb227bccd907eb91f744d93b25a684dde5e98dc8e9b1b13defa4e5807428a3d93e83365a05c5742fe78d7a018402d776762fbdb909bd39f463707eba1e8850c5305379f847dfd988583bb305f084e6bdb5851900c07fbbdf255309210a23d3155aceb1d971cfb45cee8cf2f8183633fb44e0711846891517fc8db7e175f36aa6c9e07d671db9cab1abdb151ceb0ede207bed32bc2af232546bd6f214334311879cb57cd08f6b01ab3e4459919cdd450b009962ee6ad5269f463ff58d01face7c2c4b8005a9feb62f859f7ada627cde1232982a641931d4c9d2c15c14dbf971;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5b7209e54d67a3ae73daff5374cedfd035c265891ba30930fb8aa3cb86b03c934a265d2c4325a81b4689b8a90364332b206420dbb53e63d219ce9ef594d6f2fe4fb76b1a27c3fa635ba0ba26ac8a9d28104252d98fe68e52f2fb175502fef1168af3e0660107627ecef37f4d02ab88306f7535e0991a1e2e8b4d3f6b7e620e3c25f9c112d3ad5957ffdee45ee70a9219b172faa0b9ad3d0fcbb00d09f3cfff3f2a4bb53cefc5c771ab6231cbd24539f30ca77770e37dfe74fd1f2e6b06adf74377698ec0514bc700f0a663120955743d7e574208d02608219a0602d178e38f98b946899d950148059a54e5929c4df16cce9b92948c157651c8e6ee7e2c9cad87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7b251b98cafdde543d523da960ab044ef8df5ace2f6bda104dfddafd30afe2fc42a36d78c5756c1706efa8a2182662181f687f70183b52bbe72a8987ee75c7d16caa40785a8baead201faa8d38cf80c6508eb0df2850b3abfbe938ab005fa9a6ba2ef2e9fbe0f216adba2311ad35b1e32ddaa0a09e96dc986c7ad827258fc3b6449b448787e4a55cd2c10b2b17adae5579ae64292deb3ec757ae1b961205e60b6d60e4283e6beeb72e91a03189c80678988e90daaf1818c40f55ac5131c159bd446c3d249e93e70f71aed7a06b70a907d90201639af8d4df2544004266f5951f0fcd4b5d6dba6882a4fda9ba06e6a6e6f2a4dc043af9f39687c1c933666cfe60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h588d922688703ca7812a4c6bb453b159c837462b158820e6bd542f4099100c075657de6758c8f74a01843b53d90a17de877ccc693436385f1b043cdec7c9efcaf98bf3c3da1a209466138f50f47cc3199dd65af487353a19f95f764892714a0e0dc4c1ae6cec8193b9ff04314c3fb0040a2645d9ab3bc480542817a33f2b95901908bf881853eee9e1f1062b5c5babdf3fea1fcd15e45eeda046816a29370083ed7ac018cb58c8b433cd0ba18d2be00ae9f47d60abc7daacbfb5d0bd1481660e68cc2f720087a46efbd317f08b9167e223a24a347f22123fd28e0ace1c7d6a817dbe159a2ea2e342cd03b5db23fde616505e2e17dcdb1bd3885f576f24373e43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb383532a8b46ce0160a0fde0d2f190814767de8ba947631df794e74c760ed056e8e7235749eb79eaa216f0876ba82006ae0e8261677c4957ba94171cf035042b3edb6710a50d7b658561e519af82a3525403245b3be8c735664c744221bc0b3e127a2f7e22f8e882ad59b4e89401773fdf599e29951b5be8c16435dea9f450c7efc879cb347570029cc5edba9f6f63891ed7ea252ee12863e2763f5f4145fb8c54c2d37a91314bf396b513c8a4070e9ed28e26faf92d0e15adaf1e45792aa3977a8ee1cd84476d0ac911b6e92d2cfa31763217dcc4a719525c576b1058b8a8c6118311fa16bffff07d3ae8cc69e94444b488bf0678bf2dbb7e362ea50069d069;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6266f423cefd89ff02b94b1dfb878b07b786ed4bfa5ea542e144ec4dc500fe95de9c0d4d4f5639e447f94daa72bd2a516352e63bd18701e6be0c02d1c8e0709015b54c7031a4ff09e3dc968f228843629292dbdb3171e5780719de2d418504d270c430679826f6edee2d36f50984b6779b2af27810434bddf81b14e71d926dbe5ed3883ac4df65f835fb41f24a22361a9e604cad0143b973164a6df8b522e7a0932837538ebe831dfbf95103b2cb25820933d4bd46416007a331357af8dc0b5ab83ebd74934eaf270f65be1b6dc7b5f510de8e3962e8f8e2a86902638fc93bd9d79a3ba8ed8b98f4357b339dcde201d711fcd71074beb0f3d897a2cbf80dc42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h81acf1a9f713d03d5da4befc08184d5dc42760997981e38a4a3e4e689e34f28c08c405ed6ef0623ea4fa471fdcc978cd9d1b7642870867e1e73be76ea2245609f401c44618aeeae07123ba0312af32335e711d8fc2ecce3f55f6f56167a758ab01849f51237e5c99cd032fe53810c95591c07bde231bc4634b5c984ba930b025219eef2238235cfb1398091a47680afcf070cdaefdef5d20a6722b53794dc84a368be35ecfe987259e5b9f2ad2002942c66099837e62423fb0cba8287bd5aef76847c62330cdce019198193f5802a64a632e327fd5153b68cf35e8fd0d6cf4d28918c54557703c3f21cf412233bdb3af7bb1288ec54f44ab7e4c98a1edc93106;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hec4bc2154ed09990ec4c19c57a14a7d073157449c930165a91321dda0ef9c62adcaee2a98120eb06e450e33aabefc808b15651a2424973ae7449d0fb13b40a994d2da7b71fef48f48fcc8884bb3a214d50d68fc4e0a420576c59b82344697d6bef1f80bcdc986c1fe31aedec74cf29b8013b3fcda4d0129e7cc828076bc49226eb679514b73baaa8ebb9dbe07692f955ac592a4fda691b6df160656d1876b877cc353ac92d1836c264417d3cc47b33513d83c34c4c29fbb48111c0aba2054065d623f4dda7912cb88ca5d8c04fcc5d6f60dd86a0b5c7c33fca51e5ce77d2919909ed07a82d96fae647cf2ad9e0f88750444704d0c30f7f59e3d6fef181e190ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb68302072194e59c3d07aced7b492570b90060f4727cd6285d7e7da48c05c56e86ca65c1ab55732642b9ffb2c388aabc3e6888b4a21405835c32dd26eb73637a72d81cf3ae828835fa92442cce4f6eca781e18aeea285edddace02b199b8ab9a8f00c21978a7c87b49c1fc2616395c387bb035ea5dff709c819fc433650a1fa4d6d98058737d59cd554d82fff975c13f9b15b411cefbad7a5f768f12f2e5df1582bbfdef9eec56fc1c8bddf81fb6310e601561cdc8ad12d217907846c31f2714fcb85a538c19a55665fc860befaaa82c81bfdbb0374767a9254bf8e8c48a4b653d3ebe9809929ff562cc024be3c81d69c7590baff9fad067e70cecb65a17cb2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1de48282b7b17510da6bb680328a332ae87714bd8817e34a2427214a32a8c124533b8620efdcdded5e709acfa2cb9b63b8795984a37dde27052f55369c3983b845eb7ce2f121ee4caa9b16872b69a8ad0e6dfb1ae96dc919208b695dfcad58607fc38ebf2347521f402331f71189523821136d8da18674cdddbdb5d78231d0d46845c8d9306fbd524044e8b53a2b20f0de5968b00af9ce3805f8c23abb69be832cee508b01406a7e4074f1a4375c99b0a51d895f47b4ab2fbd73bcdf7f94c74397f85aa17d7f9e4f556ccfaaa11292ad13d219631e76a73ed325ddaabdc4c7fc59b454330d642fbcc3993be6f356354bfe267b641e80a6a0729b3b5cb806232;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h600e19385249aa09505342cbe2a6623fb0a9edf3f46858103ccdd14d5acfa47942eeddf3006584e05e4106415f72bfed77c7acd22af05bf1035f6acfc9cbffd22a74833203795ea85820a40111a2b4be267d6d27438bfd61b3c737eb4ca8c1ad807f7439b0348b3873d9be3858e3fcc6aaeb87e2d23d0d3b17412ffbd75a5b518bf62009dc7ba7bd172879930259bc905eb31180c09932db486e7d6c1931c86faae8580f58769e0900001694b18fd2d6e705462951f8a867fc4b4b0b6c0c2c569bdb512c884d4c41bc677056267586a376f80821270055d69801501382a0c6e3178d2f98e7a865b3f1de4d6b5a8611b55dc9b3438076028ebcd6cb3d34872fca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4725a867b1df9c5da78eec73486287ec71c1a5a20e5deb120c59b97ea4dc21569c086438c1a173df1dc9fb7673fe210a8bec0f677e2bc24540c018f2398bd10f912c87905a87481060c02769c2cfd9bea711052cecf8a3251c7f6dbce248a02c7ca705fee727c5656efe6aee8d87e95d7c49c4d6ae34cddd409ca7420daf3801253a157ecf4ca48cc6ec5889918f1d2912d753051609043873c5aa9409c4df9701ba8da64620758aa4bbd66f7b385d9839f6973d481e0cf485fd6036b65c9e508d24fe643a5263dab8d5674734abf7d8408b371c41d19b684a542375c73a1c4e5b16378bd611c803e5639129b3c9773b7fe3e21284d6f9a9f07e19ff68cc28d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hba0db4d0e7435b6256b7f12b9352ffacc06d8b4a377ba5abc5a293e6ff9e1cc83997032e5d7b901f9ef167b06e5f8185f932153dee19769fd0b8982dd7881469a3710333630097f2def489bcdf26110350f84ed3721e8204c8b033f995396905f3dbd52ad28b26a9f1d3954057cf84a7a68955a6e1057e81e475ab78f3538fcf6ac311aefa6cae881f23a85c6e27c0e0e3be5d22523dca9adb6953b9589b7310e30ab2e99e7cdc79bf6c7c763abcc3c99a3a0ff1fc0f0fdb4815c06f686f19cd6245155e9f1c4bd46d447e1a80543be0a3603e7cc08efe60c68b68e2f273d77503d0a632a9ddd78af3cc2fe5a6c3fb962bfaf38230fe752d32fc4ddeaa94b4e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h92335a59a2976768ec714b559be4d6881929b90f572c70586ca34aa4c231f30bd42a842e4d4ccacaaeb711e700369fc03f53db2cf6f5050a4fbaabd1fc3e8e6a4e2e7de4c909c7a35e81c82dbf3451eded4a7239a9e03c6fc102f2f9456bf69300d03276c8542b7a1237c85dee1c7faa3eee50a12de3094e2a99e03e88c486a0e94db809efb0358aaebc32e35a45a43b006e5e592ef5d06f3d87213b089283051093c3ee805e77cf09119240b48313f9ccf7484c0155166f4574041576bb98fad6b55d6b15b7d7abfcbd34080774c62df05cf8a7172e902cf2dfd2a498f672e0b51d98af991f49c006dc9191e3fc15900e0512ab87134d382c40c230d348dc23;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h72afc2f3eee252d36bc7e3180330744d60a992a0d590dd2c4fa75545c93e854dfd44daf52273635909d80a7b1e319588ac8f04aa8726298b215d502f7fea0e178ec942d97b893a567f046d1b54fb4b1625efaf1cfe3ebccd2b5ae34402a55caa6f4641c69f1e659507e540e24da523b82e280db1c60b55a80a891945b7f76f256ce70d4f98fb07e1aae96a5b1609c031f899278a6d5d6a48b4b27befefd782d4d4c7bc9c58989322d782f893bcab6c1bdf40cbb76020a9ac36c505cc5fe3cecd153bf6bd60de833c0c7237f21f3addc12a24cb55792803b2ab8db9192cbaad1ee8441bfc1c042c1cb2e34082ecb8cd9b3f882aa59eae733d6ef5916e94f22ff8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h99380891611cd0e5165e7928e472c5b5318ee328454709a35884ebf566344258aa9ab3a4081f395cb6a9369789395bdd920bd2b9204d19b819fe484ba115b4f84fd16d7f2dd60fab9ec2aa1a9ab008eaaef8f542acf938733144cdd35def9447150af7e1717788184361d226ca8f5991489030d53fb51d19834869789fdc0d1df22d8b86965b96bee180de0cf0defd418919591aabcfad4f44a2be3222f6c26d05c7094d2f29615f73bbfc5c210460a07df339b9ee901c539b1e6dbc1578a72dd8e14f8b0a6882e7ebd133daecfe09bc74c3d3907cf13cd065ef0c95e6aafed35cd74d6a004f8b72ae8f67f06d2d7520815796f20ab014f72cf401b35c2fe5a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hee2bd7faacebd27844669b2fbb21118b0a543e75be6ea451d3df34bb0407f03c93b0ae5f069d1a575d9b0b2ed88003814890e23cab1bee904848ea4b7b8d2b735ec7271f7c56feda9ee02a930efcee489b3ef4b6ce374536711c4db9931815a4267fbf17d906dacc2ef0c6a37ecd6c7fdcf8c08426cd541a65014e0fb06b148704f225666a102c41a0186d2169f91538795b97f67766c5588c089c25df9f7556467c4756ec91fbe8015dd36710211604b53f681d66ea4b7f775751024efff37e57795345804cafbb06dbc39a32f17f36ae393c63514e7ca17d5bbe016e2a58106833a8b96a688058094720bee69add0947e2ba1a70857e095995820b446f12e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h59bd8b4f6567de571564f3890f3b95129f8632a9d5a96fa99def4709e04c7dcd3455a2579addcf202be4070a0eafa94a3387552ba533afc37a9d0650ce972becbba75984788320eb8d6779658ca412c52484cffe9022c17f234122c35a087b5dc7c9c6a59ddd58940bdf4ce8550bf2fff18196e711462f6d503c9daed061a492f2771b7cda714024b496041961900eeb904eb00ab6d7e0e97c1643471fac12fffb5951a3e6df83505ba5979c0392ff7bf6b6dd5d78b0eee3291c86dfcbb5ba04942a5d4e9c76a02f3205f0743e56c1bbbbcf4e6a40663c745127bd79fcaa6a990a9051d86748317c0660f943f1b8fb3d38ee0e5589dabf433abc674f684bfe12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h79b3ea58b039c8796b7ef758d5757093148d286678cc81c16302da4d4bdd8bf91c1d2bde330bfca558543c0122ca175b9db9815e7c6bde8c26fc63205e4ab67f453f94cf53af65a535d4ffb4c2deac31dadf268b5c13c851e697a60ea04bf022f6f55e66b7180b8031e7663722ae2ea37b5c02a4a2560c978dd29b2f9acc5dabee4ab4d2ca707b9897654f18ffabb52a67058eef61b1415b5d7945d512a2f7b61777d7a0d4488ec5c63af85d3b073cdce71db10e45a056131cda89321a0fd1a4c74d7844f0338decb489d46b15345c3a6723f5aca18959c72f82928ad66fd686b6ae4913f047c693220c00decd084d98c173f3d0ae8ed278fce26753412c14ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha94c5b11f14fbdab498d5a69522edc745c5b249e6a169aa9f5906602df781233af70c4afd94bff8011287a498866d986187fce0790a6172d61068cb4f64054896e5a98f6f9fe543329582f1e2ac75ae7fab475cc8503cb43e1c6e0052c37291105226a420d66ce3c2db9201451825126c4547ae7e65f808d1461a923098b6f26c0966db051b050f5cf901d483bca49af3550866a9e4d6a7380f6e55569fd7ad9f9d93647cc4b71fa369223dd0380e60686b68df73aa8ae9f384941ebbd1baacbb62c7dc0194a1181fdbdbfe341b94999bb78949fffef461815a2d50c8ef0aa21acb3651a61065cf1b9bd1510dbf0a6b2186f33fa43fe23a24e3aaecae0152f94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4db41614371612c9dbe6470177f4ad3f512c5d02f2d6b81b66ac0b02fc0edddcc42729247b6f45419f5edd7e46ddece9cc6d7da5d87e432f1bbbb3b6660423a68fa09c2aec103e23b954609ee9f0951d63301baa9de24ba81f51b564c178218516808cba12a9ed265f65dfe8e31ac0dce4e2bf3eaa5241fe20b5d70da03bdceb47207695ca8ec15888c0b3ca011e4a89a9d11524453626885534086d4ceeeb472660191ebea8caa780442e36b0a4a9c75b830ec8b8098f859d7c1b31e0de051d21f880a80488e96b21c9b067661c9ccb8446599a56f17a6d49d1e322b1effca51bfb3a9e7f3858e6fadc5f7228efb44693048cbb1232549c69bb465b5e38c8c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfa9625b4e306fce937be631bff16a402cd6e1b2be8260b2e4fffd623beaa9865f1d79b4d6d51067a60027346857a916bc321665ad216b36b99846bf4624a8601e04444c8048ff9c6ec4b823d28b427c99b52207569c1cf17d037ecbecdd02b31b225604be2e814630f0f2157a241431c7a4c962691a426de60cfa81943d5811f6daef359bcf3a0825270cb3939742f5da8687446d40871c0f747ee0e124b8ab75fc5c8c7cb049c3a76033e4ca8a9e3141047b0b8566b48a82303f782e2f699778efad5dfa00229b2609e9735cb0d8aef251354b95bdac64ef0485e9ffeee610713af33d4244b114323343cc29122f6ce3ceda3548f3ae554cefde4c58bd0e6e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6cf04151edfe158a291a272fc187d81e1fad91df6bd42838a6b2b05196b70439cb452dcb88d4a7f30b622cb7bdc8e9f5d3a03dba97a0ea644d6f3ab32b62e41300f127d01f9f27fd8f2e3508b40354191c7420f3ee500e6b0b88693a3eb9a78e68707c3ecf805e31d31d9c6f55fc8761d217f3587a98ef1fc0ae22dd21302895aeb40a0b1f2f4c296533f7e43f6c68e918ed76b10d5dac42f68d7cfa9207939a7ecc33b2ea688be13e9276e03aa73d30322327c8f085f18aef1f6b4d543de856de0c561f29aa2616a9a330da1d4967d03beed07a919c0931d9b785cd078404505cd4304df33fc84bbb0316aa1b32c6918c4a9ffcf06341a169919329e58d7a94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6fe165b102332465ce19dff76c4a0d43375de6396f65250771aa46776f9732384e306048e2878cd78e58181e826d1763383e563e92f586106f227c70539340ff481b3760d408976b011cbfd201e4660eef12289895a05305e2da0ee37e9c2be69d22d1e26418c7a0e131d5e2a05c48cba2796c649ec3e030c2f8fafbcef21a3a43e0aaa3d773e5f9171d6f49f081ae08a03464a63c8d2033b23e409200b33c1332d1225a3253d187cb34552cd38732d590f3ed6c77b698ab1e2c723d805092e6db05c1134d1216f7ab292e4cae301dce652a4416d4c89fa841dc1f18c3ec41a3a2e087a2765898f447de09294b0c37a8395848f63bb712d7e21f35fe50d7c136;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb37abae86c62d46a86d6510bc7ab4aff43715ff6b7e9551d563becda5f25ba6773e04a0e3b7282dc67fd219e7451ac564632e8d9001bdd63e7489bc1e85ea27bdb9dd5c77cf1483016057643b64da6b19d9e470a6262e1061c566cff8aa5d9b80a3942803cb808860fed920ebafee2160942504f3eb40306d329d15072a4cd12a2a0dc07ad7fb3a48cfecb9532e2c87c05220928af338f179dd5f02f237f5bafebf91c392c159ace85aff8b22fee82dfdd7f10f2f7fd0a5c406c77ef446187886d5dbc37d4f682efb8143e03f0f8a0da232f771deea67973f553244af4cc790d1a7dfc1084e4948370452604b31b3db2d51da2d839c085e02dfcba61b9d496bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he0adf01ae512edbc2c5df82b8ed9645989ee1eb94f8d5f3d83658adbf6461858d99f3ab1d9360c1a1118bff2e93bb48fd3b83b1728735d67413e985e9a6de4bb975d41a73baa91e37809964827ce1ade714ed0541bc92f6961791748bf44c2dc6c992f8f9ad23dae6a83559afe49c53b4a6e4111276990467439ddedc42d02d2f71c2c94ec5a4487fe70515c738491e22172433db36093bbb091afae5410921bc3279b9a99c38e66d1ec1bcfa4d879b9f73b4d495ea411ddd747fa5acbdfc2c132475ddfdd7f2e5d93d1977c311f4103b2e639973adcf3fac2fc0ea63365039114043a186d0c86ae6cbcddd9c499d546b002da8ab62f1546de6b407d36fc6bbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f41ba190f7ea03f01634ae9f8b1641c7505208eb78ff56e27e9d9fded9c8a0ef715616a79beafc100729ab5758c2d573341fd3d63c72f0d42c551b23800dccc34df4f1844b971eb27813af0c7dcc032027391c41e69d8ca40c93392c80ae4b8efe0a303f9a63990576c3b21b1ae92feb15519d643f332d8cbca15390a6ad9247a8676ea356b026cde35c814b58d83364477705a1a6e1a624cac5971ddf2e66fd57eb61d3f7daa5d1d864cb6f8f5ca2b19a1b49fe968392322a5d2a15547d4215496a2b8e53f6522faa681ddc8863b3c07432c441860ec7c8a28ef92dd3076f94e7745bf4096c43e6ef2a900b25f29d712c714a82fe768c9a96763b21a5ebf70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6a1938892ea471b0750b208fdaa0fc7d535c40a0611ab743984655eb618831ba4e44fc3d35178393deada0950da2e8c46e40570200be565dc1dcf059d05b5517e3d54a3a5c53dd3a0ce0f6a174af92441e79c88f2ee8941d43bda9f4652ee394268f4d139a29238cdc105458a9668808e0bd7f2d1932c7da98282b80ac365727878aa41fec003ad806f6c4e87c06256ac5408d52b834d04da9e927c7c9589182f2607e08a78ac9d7cd99f4ef86e133f5ca12b3bdb473b4572672bb0bd6de49fdf0df37288bc7f4013b95b1c2037de5fcc717b8cbb93b2f20b1f6d46c237f2a2f1712f24e1a21435af1028b9d1d5b3b73bacf9d0cd16140d5a591a0068d0afcf6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4941a967ab5c3aaaa7804776a076007ef48747d2d51c7fa19f6bbba83dc554ec8eb2432fd001e9e8ec98f2d53b6d23c7b8cd71b4a05391b76475a0f2b6fad19f40d2ec278b0bcfedeb38148595b981eb5f0467eaed4945c5b52a6ed05133846bb2a3ac2858d4a6307530d35c55673c568ebec6142a5d10567be92d185a6629fbb64f9dd985db42f417f17448376cde8f39d3a13899745121cc1884116aa63943959a8242f452bf0451f2d7a3a4f43383ebce86b92feaf006e01a1bea18817938db37abae4fd53370050c8d993a46921093c2fc3f3ed6a5196525fe185b7859fd94ce28215f72820c92ed89e8aed96e8f89a90ed860e15e6c776aa99381a0cf60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hba5faacff368570699150019f8462007d30d302a9dcb04be2bed17afe8dfe2bf3f9010f87ab27475702d5b05aa2ce6b10d3d23afa4b720a7eb17e75240c8fa1a9f0b4844fd21a7201f64220b89f4c95524c3d1c29190a52d8f9f694825f0d9108be960968792980d3b42fc0e972732227f1061630a8d0f12c4f1cd3e4a1d18cf5790ac4e90fbffe69285a28bd99e7b31ae65e0057c409b9ce18061cd3aa41207f33fbc0d7d0125769e482263358165c1ab4cd7cbc283b5ca6882bba6ff2abe1e3cc487bbadfbe3afc63f2b8e06316fb61681bfccc7ebd4749a355508cbe42ad17231d6bca5d5d79afbc028a26624390d0e4b2e68051de53a7f9652c5bb062a1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf6df9eb30b5dd28a327d0695753c911b3f79cb22b13ad5286fd71c4a389c3eeecd7e1669f226db60e3aba115b6997901d2bcfe6f7eb2eff19287a9aa8024fb953c15395832a895ca2e1294538795721c854d153ac59724f5a9a1c6693ff2170b4e5fe47950f10bad238cb3dcae3daf893df129f414fe2d9f064e7c250f5b2ac4ff440b9f3d58e9ae20d552af21effebbf79bc450bea1806193383c01e447cf8b8e530c8a33dedae6f07cd56cf9ec43b34ea96c8bb43f7a3ce639b730e99f903ebe89dcd5023733ae30b2cf5b4c1f0846cace0a3daaed19fe28e40c58042b0ebff57ef31ca1b28d6e9d95264f0aa4cdefca134da49caebf7d93474f17c83ea740;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2f2207525a6e20f66e0107a63b815aa4f26b4162022c153ebff42a1d6b436cb1078d7d2f85897b76c0ec19e34f98ae19e4663c7da1bb74ad22ad6de4eeb6e1eb1cbe5ac321f2e5ccba67c871065ca6a20c5b1d03939e8f4381142ff2c909b2f010d1a72e1f90f5ab3b995a58ec697dd39b49560417d8baa5ef13efbc03c0811107c1efe36313abbd91af20f15c26e434d6d8da6ee10eea3df016911f13fa98d4c02966c8aa18c090969ba3ca285408d5aeceba923cdb9f72e5ec8e23fe71dadd57b43ef36322cab14bca00f416f6ad6aa0f6ca6b01d7ef096d4a60abfb72e3bbeada2951266b08312cc91b3d7e216d3cbe77c7c08a5353e8173dde1a161ecdb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9fa44ab07d439e82d75494f1138416d02e860a5a8ee021b720ad8168a872092f52f3fca4fdd2ccd3770da9098acd0103b407b43a887d3f0bbb8eba8db371cc45e0cc449db2ba5057703605e95d7489655b81a19d82354dffb7b60ec0311bde5abe70f876101be8388077bf245175736c48a2a782367d4a11d81ce0c28f92b27f23331e3058ebf903122066af85524c83ca8fb1e6b0d1abfb268c474ae5db6df6c8305269b228d0212585d09ed37efb4fbc42778232734adf3104f879ef3ce1d1f9e193a046da899c75488cb7e4280c4d2d888314acf3834e64b8ed0daca03deebd162ed00624778c6150bbee6a990f3066480b61795a1f7f274add855a0edde8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h423d31f3f496dfab28d7ec4d6137336718873d8addbd66da8b7f18fca773c2f68e125711ba3072a20db865d95129456d88789383ba7398a4b82f9f5cf89381c9ec97a249a41a892eac1d6872046051fa9d18152f4ab81604f41526d6627d0257ff2049f851abc2b803134ef936e128c0f2ebb478c9b45966aebcaff491874240e9c586d905d502d73fae55e63bed3a8d7b5d731b13880247405ab5b9057e1339872dd2858d6400bac60273f80dff7b94f745065a29f9736efcc2a7ca193b18f1491af37d56b4f6a56179ffadb41ea9b8b41351869875e7a3924a503540935ab55ac451932663a37535f51b4c5cbbd95f9589b1c086cf9e3d96033e123def83d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc853ec06760c2d772fc6bbd95f1935592e4055e5c39a2c847ed2868d74975bb5697390e643510d13f433b5c1012aebc22669983abcee949867070577cf5b012a768b8b0a4dff9486ff8a2caf9c190040410a5021ef4570c906b4d757528f8e87fec12f0f345d953cfdfd0c18558d0390d54cb20733d58bf2cfa6ed352ba05bb7a107990178ee7a67a2aa20e8397933a6bfbeb752165eb14230b0c541564863bceb3a1e75d2a7272056525a651e9358b7dd885b48b6d7ebe718bb094dcfc635bccf2942a42154cba1edfae35734c4b162b943839dfcc6029f3ab8e229f310684d6ab628491b34cac8aa370a7dd34945f18fa0fc0193967f4a4eeb8f14943ea212;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd699353b6587cd0f378cbe3b9efd490ff40f568ab15aa663034da08ab4126e2081b68639d84bb9def511cdd8baabe402554ce6071623a52351780366dd1540874085bbe0955d6a1b916b713de8b2aac28b6b2be1d1d97018976dc88774129b037212bb9debc69e6f20d8f89c5a935fa5dfb945a37582bb5ed898915d5fb95bcf8a792edc36357b82712595bff4b91658cc0f0a865d0352cd57d5b46983f1fcdfbc199412fa4270cd1cc7fc58d385fb0c8624c3c060564e4c218be0ca6b382cd45a91cdbc6d36b1a326ac64e921d093e7d02261b827388eec164aab63207698744d4128553b275f312e7837a9d7037417d8d51e78f739d4e0330a802c4e1e5419;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h72b473a1195dacebe3f30deeb384a17611fa227d3762710434072f3fdc11a9854ed69a64436ccf4e1f6829746edb1067ae8a08bfe7df14eb4cb92457065ffe5e2f885ebb6c2746ec9610b864f6ab7cbd084e561f3fd48a8a89ecbf43ce8a5b04672b19f1b67f74afa84219b6362a16b11d565d918b69f8bc5a224803274bbd4b2cd4a8a7e3dc689c47e06fcc1e563cb06a0765ac2d0bbd8d2e9c6ff746698e953138b2090b1c9d678b32d53dba4a9f6358cb312cb99d73ea0917678ca93b9c634b344cf677d509e5a3f4cd12456edb5d60fc7c245564ee7f1f37a021f7e3a1a71b25099df224f5c3c21f8eddafd0456b27b8a6f7e333ceb9f4118e65f73ad1d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he60553c1d714d97b6a8c63812d511273b1ed67c4f3e9d27e276779b28c8a395331eea7e78c329beaa26d83737abaf0521e46e5312e2765e4bc737c1fc6aee0c8663a799c22a671b38c67101f61da024eedbc7fdc94603931e57a7b973ca264cef3fd066df2e6532aad34d31ed4954b8da700ffef6c9e67e7563dc8af1defbde82ffc6ed607b9c118d7a5b0f5d5808216d185d9af01d55345f1803399e64e4afdf667de041c9d2d5b2584c15f86f0ecf2820e250bac591088aad8e1daab7fc9575fa6e6ca508afe2f00b6e3e0385fd43ccf4f47b38cda50cb475b35b4f75e5419b0c925fe7063e288440193c97168b2d45729644848e33afb2ac17b9e15052a9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hefc81561f3ace568966e7e56d25abda5ae60c0ff137410e7df9105f98a5101ea2e5ed3a46b1383a8a315238feeb2b9ba2c122e73dee106965651e723d718c224f9c5f423e26ea5e4e6cd9abdfbdc9e108b8c4d4d479c736966a8076cbde1f607ecea51ba09df89e4a47f8e1ccb100715540f4bed2ba4592bad64113fa4b6c64c1c5d7074c5fcabe69a2dde36a90323c67d474de5c9ff1413dd7d5e478123a2a668a491b92ba220e2e57442b609221afb9c3f662bc241be228b9acdd90e6bf95b96e33bfdd809e1ef395c42e95082d916056071d381e99405cc7e21d964f847e56219d2634d774908647dc8095b69addc7457f449f956a5798d7cce8c2eedc167;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc457ee17b274eefce0ce566620ee2b35f6d1185f4cc12fd8e30b744b3e43e94a5758dde03f4604c2460df1bb6b0b2d4d98c1d73fc70308384d2ba0ecd99b1e514ca691a06094a08445e3b73904dea91d06da0a02c45b3db6f66e578f6d760e003f0dfc45a3b7ee13abf36234828a8351aedd14670c2568400ca6f046b089b2e03e080e637342c39176f2246cdb599f3e9dcb2ea6505a20a5a9acb05f57c63efea55e961527880938a75ff47d614f4d197a2603dd8d8c61cd42c968627073dfdcc5e4df646035a78469d285da2c7a974acf2feefa23a139b37ec017a84cb0a15e36a75ab04714d90935a0151d0e1703f1dcd09adb40ad51973029aefa6fd94722;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h40719f085c237d3709cb5a65e887cebee4e98c38fb513d40e48c149a110a024bdc01b4f44cb782330ffb1b4c13a105e41ae43b4bacde79055c6118b1f93c4c78c81e83e252ee3b1c2512b645b75abf83f027301cebd1a82143ab15faa92b1c99b0095f45c02eef2071d874bd6dd1c83c1fb2af63e3136e6f45fe40f6659e6793adbc5a24132074a1945947cfef113c86804248802b6e69d01b0a8e5e813f6b39355ee17803b3350ac2b118d9deb5be95136c7c795ae026227eff99b2d29fa5e448ff2561cf1513212f775853ae98ec5e324efcb6c6e5e7d823a2a4e15674e52fe437c03236191b2b2f23d2c31f045774bdd4234a7fb8e9179897914681d76b8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3075bcaf1dce3bd9f487c2f3180b48043ed53b781eccc230a41bbb63bc4b51c9d51da8611fa8dea5a92e491c94f245712534e09a5ed410b70abaddeb1230a6458a9ef34db8fa979191afebe6cec80075e2948e8d1d0120cee12edf4415080c16845fdc9a2fea9956828cb24417265f0f65b5ac90c6889b0d0d2e0111afdc121f0bacd2e1d32c6b3c3daffc726b39911c732c5a36bc6a724c731b6a50f3a029317edb771aaba12b9f996ee8702dccdfc2fd11a58f5baceaae6760213cb889b31dbd26f4635f3471295d26e39b0cfcc9fe835bfbf54426525427339238ca10cf0e1b931dd998bea67023861796d005261d358ca622672aa19400886d5001277441;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h383abd75666ee4639348c9a9c636c389781daa39b0f08fa2c40095c52fa95b4e088de82821f9781a8eb415a8808126d67401a45d910b93836e70fa81369ea5487089683b10a76c82a06070922941591c7b15ccb7ec76e464a55ad9ab48aea3b66bc0ac558dcfe8a52c5b752025864a5ddac7c3c6cd3cb9103cd345470f1b9102318036f750088c5a889a605acd32942c044e455e83e9e69c9ab3f7344d58d218d6942d470f58fb657fb329b09099bbf18305433ee50173cb991678468d65e881cc392ae54146216d429e9eee016b2ea40f62f2dd49058b02736f464b797981d435f91343f1d24c93f93e23291475869665035a76b9517c02db76bbd49184c8d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h84eadda09ed86b3f409dd1e078a52079b1c41055c0c24d6c4d404b2e6143c973bcce45683df5beb3d9d63d2257211924dbbcf073b3010711b2a72637d51f52d4e242a7257ef6686535f4166de2cb34df0f4194f8ca901a35c62358cf87fbb2a018afb00c9290c4e16b4738d4c88bfe1efe7752ade388783787608ab7761cc2754233400c7900751820a179fc6c612fea90e5e82a3f4a78aef709d11fb6660de7c78ceba0b53f54ec0c8213dfcf827882929319f2b4a0ffbdd1aaff0e43c8a6fbc6de3cfa77473e8ffc246370997c29ca9209e6e04cb6a605136763cca30c14c0590951225d51164ca32ce121e3149af9b363479ae3f685db5d59a83683447a36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8d70c85a233922dd43ab4f43266f5d20ce0f65f8ee0655934201a39a30c8930a4edea4897f5862e71f5984b226596a33ee05d2b5e1df1f8fff0bedf1c5c5f0847f0673c45b0a2b3e2f9e256f73c7a0e283991a9b01ae8095fa3c00024dd58640cd14c9ca28dcf1366ca83dfd84d8283805d1b4d973a083f4b6191cfef86ca15e46a47352c6f21418417e17ac7e531d7fb6640e537665d45503090c8d0bf659919ee1d70f6bd31e5b14213568f5492c1d5a4e0f4cffd0e451a11b8108609c889dc45d5edd8bdb5e803b033acfda57fa57d69ffeaaa2c1de48ca176c0182811b29d77e6b31f7c5efad1ecc0e7dce1aa31fde4a26f22b46487770b4d06f84fa14bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h639d6f51a100dcb84fb327017f5aa157bb42de04917d9c00fc337732913144182508ff183e6e5c5a6bb821de12f743a4a1dcc75a426f75cf569f13a0149ad68aaa544db2ee3f6630f8dea448b48d7b81530c53e620040184bf771d69b70a8209cd5bae0f74cd6b1c181bf83984b67d978f9d05263fb815a210ed1c35da0f1e4ce1d73525b5f22d55767e4ecffba4c0eb68a2b2fcf8f8f92441c7458eb265edf9846dd30ad96744d396919a1aeb4cd3ae3c7b657caf74ea273cfd8f851f77dc02e4ab3c924766a2152ba25c1c07c5433fe2bc8a49c5762a533faf2eed2d74f674550923c10da7b730a199b79b09a435947d13bb2eb17a512cebd0f2752fa80486;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha223367914bb3fb1ddab0ad604a63ae922e96e543d5169bb24434cd08298e09b098aefa764c334e50f1aa8f9643fc893d508797c408db9534e6c41ee385075c74835dcacf82ed1fc46a53708b61558dd721a8e243a8a2927d749d0aa3e31c3a37f8488b5b77f81fd1b70faebfeea9562a3570fcdc2c3e5f992f83f8d5df879dc72909d0937a17f5a58235dadf4380212332165fab48f06f5b22dc4d515f696b0f58b58ee245eab0f264aa30225283d9b457881ce9d5456f7c243256432a78946c4929a168859a1c261b9969adb673b8235f1aaedef6a77c464aa1aaf84fd853f0654631634b4ba025c20d3184758c779ac6b59603184b35a68634af3e7ecd165;
        #1
        $finish();
    end
endmodule
