module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e2fab392ea436685ba41c84c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5b8dd3f45d1d36f31522d076;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8253304a2c7f463c5e9ea9edf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2feca2dc71237ee6641c34d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f5a1187fcd84a9c629040bba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17e297e2c889db7ebc45c6c9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heefa01e226a22cbf53a6dcde5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heae02485d59f61c26929d6ca4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74c0090569a4b708631583f4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cf26f3b29a73baa47c8cc488;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5727ef53739d05a7bf0a68677;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf03f611c15a7b64bdf04a317;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3238356733460a4561483282e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbeb572b031819a00f2decdfa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14e4cf40bad80b0841da5e20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f2fd9c56427e59ccc19a8ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24dbd13143f518021a5989bbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd86e273d91a92b71a462e4d9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b5cc0ea8bbd84a6f1e21066f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17342b4eb1edeb133b48a3431;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac0e3253898ee87596adfe2fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3f06612ab05018b75152bee5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc12841a823b016d8e47e3a33b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb97f01e4b6cf424e0b7ec5af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36769dca9ab77733b1d941731;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0ae5443624f2c2d503c74fcb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e389fb83806debd27dc60da0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21a080e0e001b60b5cf161aca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h573d09f403eea61efef3e424f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcc22da23755d6802728a0625;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadce67ed572522d8c6c7350c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde963e13208962f915a04d972;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73cc3de4b3359c0f7884aaaa3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc150d3ba1b88120910cbb676;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1f0d67065da733447aa5550d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae54e102d20af3ac542900b7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39ad6d2214b54b12650403529;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb27373f3d19c8218273a59bba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc809c39bfe46301a315484e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h172701bc999b66dae0c7d2a84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89b593caa074f2e324a8adfe2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h427576cd84971d2ebdeeac790;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0780a771f96ecd8502d53733;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2df70b6be73c70f982f79c24c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9c5b0f9c76ba4bd5703d178d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7f640e8c8841fb847da49641;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72aa3328a152ba58d8fad3ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h915e92f960e5193a7e1c92a86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf27e17df6ce949d259c7b17f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3fe84a6c470f738350a67bcb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h633a2d52ce89a3d03b4de4bf0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa81255b253ae510af6eba5e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf296f7df6de4a4767c9f06c9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d06da6fb65f64108323e28ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf60b0cde405729264eeac889e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1ea742692870af340af1cae3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0d088c196c942341c6bc2d4c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78578eca4180f4a464c292414;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f52f7138ecaf8be4aa441510;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3fc20e006330cfd1db595873;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f0cd460ef09745af3585410;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43a21dfc9558f65d514564258;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf100f099285dd0bc191588e1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd18edc52b06959698a29d6a8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd46c04e95d1198711917090a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3f3833beacf7e663005732ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ca5fc0dda2ecef659b5796ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28e24c9e43ab32251f73ee53a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d47b4cf2749bd630213eeb80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34c07fa2adc8c0f76bf05ce46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f6b3d93100379f88f8837ee4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6115804c67be293225e464297;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcef3c61cae1ca045cde9803b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb3ab64a95d3c39641ed7440f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4cc271c5a41d555afba5844f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1839588a34f301dfd7616cf6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd8b1e2d135af1edb2b70fab9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h913880263b67cf8cd62ab418c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64c6a2ff8ca261f3d3c8a6250;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e2682831aeabb40c62ae47e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc34b2b99ac3a4ef53cb48a78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75d78d9501a3234b738a75180;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79a799f156fc07d6f19ee43dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e2539569cb2c4ff818b00759;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc459b1bbab76e3c7989667ffb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf41148ad983f03d10989f8c14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4351edb1c3b48c474baee0b02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46000c73041753b0bbab824a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdbe2077588e824d5f70bc7ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8beb9237381c9f3f5dbd92ac3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h170687c7dcba93559bb3cf39b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3f276a9318e788892ac4210f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h993c7c3c5b729161784f7dec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d0fc6fe3bb6965e8d1667e9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h429c0d5b1da752bb0c24a8f14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd24afae13176319ca4fb75bee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3102ad6bc667bf03f00745bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f4fbd079611e99af475574ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65dc43299997db3b28efd53ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4888db88f5b199a707f318dfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29c2f4f19df3ff82a07057de8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd85259c7f9b49a8f4f1fa5d76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf8443b59873cec73566ad940;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95ef645e6702efba6ad67ffaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb73bb8a442209d30f573a72aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83a699eb5f30814db20da19b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e38af1570533b020dbb8ea6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he612ee14c0288fe185f8d937f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7234ef24cb236da2bc647839c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd79ad654fa1300137f7148bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h234e796c4bb8583b45ad51801;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c6b369d8b110552fc9156a76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b850e9073e9b0358b7087d8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6598afd3a9da2feb2aac979b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74383651ab99eafc3e6520503;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0d1b4f3b03cb90f379e58b2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf85fee402aef569172b00b7fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef9918a8342b87c9cf21c259b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h793c29ac73467d7e3afd42743;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h460cfb55a9355b47ad23d5c7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4e96ca217500341837987feb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h305a1680957c607eaefd2c78f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59be06f28b4169db23730fd56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha334a2ee10e287167cc15854d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h672675098d5ec6b182248d157;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56ce2a0bc4e2afe67e6862858;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd5c50eaa07a0077a7845e230;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63d5dea8fe7da46ecd184b9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a1cf226621c28e6e13fc2e9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cbb3d7f1bce4b533a734ff82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9c15c69d1e74e05684096884;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b58e5bfc8841826bdd265db8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2a0783f31d4f660c35ebe150;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48b659ccf8c2a5690e56f87f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bfd58c55a34b1d38027a88f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13bc0a36ea52c4ef7a6aab8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8f9bbb8e4380e173e1baa886;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef85ad3c7eac3bb7a5c90c3d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h925a76f2052aae0d4324dd016;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h476c6c331a05bca56e040dc9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddfeb491c55056b308141baf4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bcfdd1f4330801155ee5393b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha16b9bfebc8bf5390ce1a3d5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43c8979e50464fae2ff3c1d5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c564db5d17b867e45197e2cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he91dd5724082fa45c1d176514;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h889bdf0ca74171ae03b80478e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2d3c51d19d353c01be8f6af3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88d8c57cebc52da1951349422;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha61cd6f4209c507184f9fce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c2829f667ef777f4bc5c9650;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3100b996002832401fed7f8b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef062bc738c1d3932d195b3b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb062bc5ac5f073d72c7da1ca8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd96dee100dfb8f8c1211608;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4898c80da945fc30a32397de4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h176225c48e534261cbcbc54f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fa6fba4794d611717afa5f26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59815b4e0688b51a798a54954;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h896db2f208b7937a90f458148;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf70dc15311e714266b4e7d5d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8962a30b37919e475b363be1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cccbe23e4742001c8289198a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5776bae3679e6ef242bda1c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e5d1b5d1a82dc539c5a3e768;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0fe5b9107f7f283d76559533;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83baaab1ad385b01d16683e07;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f9b3c2ad70dd3eb8eec78c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4425a0ea64a0b4d955af7fe90;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb63310e30b084cea01a3c0955;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d7bad3d056fb90ae83f7b15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e506a6197fe25643f4c36c68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3514aa0dba62f39229a6e074c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd36547af81789d89179ac0ef9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2a4edb1c9610bcdef57f2cd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1192897005923389ee8604fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb17040b3bb6a75541c99837f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9272211d5d17bd563ce00806;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d7baac5647ee84f0ae9214f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4031fbb3c7f5c8fdb1cfbb5d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7415fc5b4747b38ad8dfe785b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b02b1a26c7948ae2718575ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdcc452b3a5a83324d6270272;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d0fb3f23b48170e83fe5805c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h717e6ebccbe363b6c4d02da73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeba2c7c3988e30dbdb63faf7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ae28736c7b0f331873bd9d78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6aee4f32f64426f8e3c201a70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fe28e4affefa5f1c4ccc79ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e6194d34d10814b2aa1cd4df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8c6a9d2796b68751c187d291;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfae3d0ce181231bdec5360f97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc24ec13b03706fe81a7ecede1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee32f31c7c40451336f1f7601;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78c7edf65865ddb00b7017909;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69ce188df26ef619ecde9a68d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8af67e16d6ad16972872027d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h349d0357f935d9e116884edd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1392423909c60464da0cc7870;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5de598e48d28b9ac4fd7500d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa0924062c5e49c10e17122a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd296e51cc89938367c0b97ce5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce8aae3526da7703504216dc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haed47f3a7fcab34aa3ce676bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c5822e79f4d7ad3f17e56acf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h294572ffb7f3a93690b2a5987;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffe6b55678d7bc9489ef7f45b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9b6b205c07b160530d4f572d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h411f4d7b9d8615f641c8f3179;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e2d7cb1e78fcb2412ae5e50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd666aea1f244a91d78e728a9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29291ae0daa719f25f3dfbedc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8a382ba308e4f57268ca8fe4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h900f974cd2f242177f4687404;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53843f071a0ffc5bca52e1b90;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h817197e5f4c29314c0267b4cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbee747800a8093b9afea4715;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9627288f6acd9418cb73f79de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h756055d618dbb9ab5ea7529cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83a18fbcd7cdc8d85d5db420c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61db6044c6d5fa92f767fd73f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6218904511fef60a44f3e2855;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h519625634abd010ee758c6697;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb14219b558bc03042c82c6714;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc16f586e629cbb75eecd0a223;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h623321d6b260a8fcef2586db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0db7c51b40615d47622f68e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h711ad785bc3299c1aae746f2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58341762aebc13eafb39864ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h752f500f7dbd9a031ea3d8d8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc243b26f1cd44cea8c37845b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b74a7a666a431b7472403c33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2634740575ea1266b99f14ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he98445a27fd30d37b65289810;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he70e1ef55ceafacc4373e4163;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5472e749989ae97bfb512d7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5361be0b521e7c1721415f7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb89d04c7332f18b11a0f4e9c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce5ddd8cc2e0412d360c9cd15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6d88c71fdfaa0c4433d3f65b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7812d644eb722dc945431aca9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc331f5f3de3c859acbf33d702;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h885cd5cb90908243b49582770;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha30592cd5f803fb22b38732ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb14e9482aa9d75a55e19301d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29c1bc5449af36b12811d373a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha47d10ff5793a0ba909592c25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56b099596b54c393d03aa995c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4080672532b04e805c048becb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da35b3df07b7a4b33143a70b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfc4358696559501770217a18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87317e4252469221d5405a9a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a4734670a8578b1bae2f6d84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b016c0ea26f4ed5fc0b05cd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75681882f2d88a0c694f46c81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17506a1c7e866c93a4192ae84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa8d5bf8d5d31a208451ad2b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14f16e2d9bce24ec75bd699d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a3cc20321cd27c8b4f61a595;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17841490c28364e086e0fbbec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d1269ee39e5b2dcd7993e3e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d9034292ebaedb3cd8947c31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91b194cd7f14f58c9e676f559;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65c4840df23f5f615e29c8e68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90c60db81435887b203f7046c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h639868b5582c5e2eedf719549;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8aad032150a0dc464f6783c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heed6f32818dfb86827b5019ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb892f0635b430823428c80836;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha57ed80617ec092906257c551;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h728906305275306df289739a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf00442e004aeac258c0c08ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1eb7cf1d22f8f1755add9a15b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43b603703841260a664308cec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cadf2218287e2346377a52b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae78b52d6868b06c8be06cb64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ee7d0ffa18c09140c2aa0085;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde45240ea52eaa7bcf5a97097;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17f674ca3d72e02d20c675a30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc47abd82e8d70a9ee7eff0bdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec04b632c0ca17676af17d8a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1416e09a9c3461916f840f519;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82c66527950e38678b381b57a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbc2bfd7fabd3119d103215eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67becf053f3ed45d3f5638946;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9aa1af77c6e18ffa966659d66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33e2c59c0a7d43f6951fbae40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1013e7befa52e31c105592b63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33c9b3994300e3ad9d0d7630a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7a8681daa6a3e55d392439;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb35b41c6747680835a123e125;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fcec7ee9226af7d173199681;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0136db7900259b1786f99c06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h843324134589b5e40c9c5127c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf22afb594ffa783958490c2f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8abf521bbdc319033c593bfa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h681d203cb03b8610a8b194f02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h906a6662bd4e7c9aad6033e8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa4f4e1272e2d3b846d79b7ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae35c77479300c134d5d860f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae9207f9cb33ba133506d58d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc192dfafdd99eea2bcd1dabda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h410874006b5b15ca3fab44a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fc50bb0fe446fe7130f24bb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18ebcd632d92ddde9598f479e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1f54fe7a4e2f530462fc98e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d3a5e904a9e6407cb8aa2d2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf5275b6ef524a505e1d5cbf2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6a1bb8e7703a3196e3772abf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee730de1a6502554c029a1503;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d6e14afe28ab853452e867fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cb56e482f441d6e499417117;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a9eb6f4748f53f53142a1cc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30b0e76d825c752de34d3ad38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h111fc3758bfe10e7b2f5b6c8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19a189d3b21725adfa377a5c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c160cf5d387b478e07d6b113;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf02f9cb5e887e2446df2ebbca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb650db2f341d44c1caec3fdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb88642541848ce7756f839a33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba0b1e871875990d926af0907;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53dc36aa51ec03a28846f0f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ce4580a61d6b9a1c8c25b278;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f2dd268a0825c2117d2a7e61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18373262038603d2072db320;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76225c1891079bae341de4f60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d1af6062d51b67b26efec2c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fab17f9f6eb8da9960541ca8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h587e13e6c97d2dc8b03babeb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40368eee5e4719da4e4eb1a1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h669fd9b00609a38476e9721c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc96bc0a836c1d04d681182ad0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h440acaa6b2fcb1ea9611f8c43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ddeabe2f72f6a33e68e53df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8df59e2e5c1d1a483e18d409;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1ddf62d60e1546e7e27064b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ab4283791f9f27381d167dcb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b28649a7c3d7c8f8a48a53d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3a6f82725f55be7204eebf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9da56339a5de1479ceca4e937;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d485e8991c999b29cf4ae046;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf051269f7e0e05d0cd326d10d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h247e5cc3bf17ed5ab6fdeebef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63ea742005bebc29fd30035be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab8d22f7ccacb04a2d3012b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h929980863473a535ce7acba53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1c015573bb7f9aaf446fdf93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1917ada36337564625a6227a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8c414487208a235b035a7c65;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff44e090839a58befd223c5a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hade80d16c7869c99d9a0bacc5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2dd786d3436719c734c6511e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee08fe92283b9a12f4fdbb345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had74dca58b21ae30bcf25135d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39aed1a9bc0aaefdd807acc08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63d3da5f147f382a45ebc18e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35ac7cfcb9f25d20ed71224e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b260fa682d9e3b6aa103e1c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7ffc3f0e1609b7fd4f0c5cde;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0667ecafcff4bd052c3c4c7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5c7566ae17bc7de02e5e99c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h783bfce0243b40e1d8530560;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h219aef5e06f09db538f5d2396;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54f006440051eb85dfde96e5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34fe4aea2ca037a5f3093414d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h864f3229d6e485558871fb67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd52010e07d6eadb60bd25dd81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2c08a0f0060e4570ace4c290;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1d11e3a3c5545158d02b4e86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17324bc067404363d7118756d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24ce180fd715969d02c78420a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6b360a319788ffcf26b462cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6613d56b2247e704b350fd82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51cea2fccda9bd34bcf30305d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0fd0ffcb2832f7e30a41c273;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h464348d3a2e83c001694634bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha580c0f20bc23ffd862f2e23b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c81959c48e1c861f26b71aaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e1cd25e6c08bdb49e063dfff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62e59619a9df11855d42bca80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb534b4a573c74beb372e27892;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha041d7d11907eb12f072f0fc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3daf6b4d40f90a4bbfed6329e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h148bde56e050297a0900359a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4017f086ed12ecfcbd2d0d248;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45245a48c6f12224c4f866c16;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdae94ae799100625512653eea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdeaa0630f98907f5ca1acd3ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c2b6a1bdb9948ca010d97d63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9be55a7bff798abc5c7a63e26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h970b0f98c7343c4e181e08515;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h717e0ff1da7558eb55fc955a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2fc829e54fcc581d778c5300;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fa0c6244cc349f0f8fe7c401;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h371054071aa03ddb75f731403;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4bec4df05e9ce6d85ac5340c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha59e9caa42cf3effcfb89e7a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26c5bd94c2b7b1e4a835294cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h809463bf9a07c05323779957;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb54e405d82723d73ff47401b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49cf039e83cf9df1ce3374fc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ca0d5184053b622d06226ba9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h877b0566df5a48a7c897846ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ea70d96da00202754862e4dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7694a20f9d93ac23d811fb8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3de0ba1ea7a35eefe583c0efb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ef6e4cef9e8b56fe40265b96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28027f81b2bb673c06cb25182;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba3e8be51b0155e707a55e8ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h933b8273aab845be0c5e649cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha11b6ba574643dd62614818a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4fca24036ddd6e740f3162c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b39300912441d3e6f0e6a620;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce91557f8b3e9eb730b7ebf14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc16b4263158f24d67b4df50e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8f25ca2ddaa44e90ad6263ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h444125de94a37ac9c2a569e67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f71d2829fc58f9f38ab35da3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d639edca10d702e559d0df75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc69e0bc1eccb2f11ae3b0642;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f3b8c5204cb42d8bd469e5de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eaf217dad5dde91c3f755904;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8de7d82a2e4708bbe88bcf81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8a4547e1eeb706f67ee7e93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a7e299d52fc32fa477cff81b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd8bf1dca8c2eaaf0ce0b9cea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab60718ec4a22835d74f97bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83edbdd975ec27f4da53eaaab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9404a92ae318344e5f9faf747;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab545e64cb6d18108c2fb925;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3ba1eb7229f5f42fd0403e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h942a09ff6a40a30a72dd60084;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e62de6109041157c5b1f5fc3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h625288abad84e790a8adbe373;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a365843a7497913f4d6c0b49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha325b67f94f695deb2d139e10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd1b30368fde97008cdfe0c78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26a5bbfa4b2e2e332d3915f6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf89a77e10df2e902e9c960f71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9198fb34f7fa06fa93eec9178;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ea749353b1124933a0e3316a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54a40632978ab45f9391db85d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32df66be4d42770649a4a942e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f9cceda34ba303ccf3364d0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h633ad5f4e6452776358379615;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18125eab8351cd4fed081b190;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2c7aaf4a949ddac077060147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9f7ffb07190f1254537572a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c0b4b120a12976981a8af20c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heff7946b275e1ec845bdf8ebd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91ad1b409890f8286093dcf75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfa36409bad04ea9fbc57ffb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8b32e483bbf96c2d6d751d50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dc234a34852a2e7faa55a50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfd203c01c3bbafec46451b9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7f27e88ef16f28f9bca31cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5f6b60f2b8a8e605d6afd96d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd725653fee68cd5ddf28fa7f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h622386e3705e495648d23b932;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1f34ef75ac535be48219d15a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6eb50f3700a23e72952c349bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33cb1176082edf109b0bea9dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9661d49bed425bc9c93d28529;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85d9a1b8a5aa872d963622335;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3aec4d2f8582e719f92029492;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12228a52fce4a083492fc75bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h874a29b7446947b0e7272c607;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7fca00d8460072b7cbeb54f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1e5b51cf694a8eb85b4ca0dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6c2c7a9fe59e7a43a1f5cec2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dee81aa9e1ffb5ddf81f8bad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd28ab9ff2fffdcf74e3f27c98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc11ec30a7e35df75eeaa7417;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb47940df501eb92e1e33d7ca1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51e9179f5fc8acc161cabb944;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f316b0be1ce808b2d7cdcbb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b0940bc1cc54dced559490e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21e969343fa7d63b11cd0c5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62c4fbbb10b7c81c67b858365;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a7ff63c96e37c32f24f4c459;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fc98a7bce5b8d01ed60a6f33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h281e7e471612a8e6f8356a9c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7763b2667e5f76c3183f52416;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf62dcbd86aff7fba2ab05525;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5a72bfdc2a4d193fc7bef0c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9064a377af648b0044f735b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b88ff8861c2475a20edcba1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c6d37c0fce13c3e13474c833;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f2cd6edd13614b4fe6128485;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b7b26d610c806265093f0b8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2146a957ba71722e30c862735;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedc792b299027a74f512403a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50efc6e329eb16ab741ac29b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a9f427e788716e551ac53fb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ba84b97086275a6514dd6f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75f80b8ebed724bc60041e777;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aba5383a87114a107009304d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24cdf363bedd83754b4629a9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d25ce6c4ac02d6b470593b9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2edaa2bc20b6bcda914cdf1b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h718f729f8908ad772942b4e52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a14329ebbb2749f7df6c8671;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h906a87cbd457bd2a277fb3d49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7a69a6ef71c104ade548096e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50edba1e9ef7ae3868584cd31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9dbc589c12ff3aa08b120048;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0fef87bd59060f243969be46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ab724e9198a116d69ad40e49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5d11519b32251ae706bcdc38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74ab20863bdc0fa30d440557f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a4d431b34793ed6b7ec6da26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c5193f5b577cba1700a57397;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0e9f9484256a899977a0cc75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5db096a4e27a8acb425f38396;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4de55f9877adf1290898eabf1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7827318366ae15d274aaf5e0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ba1fb7fc3ff421a88094bbf1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bd4f234135c5045826ba1549;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h578c79fa7555b4a5490619efe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h162a33a0d9992485e223eff8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ccb32359ea3c9e636a385b35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa72bdef7f03111e84467deb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3c165b0ba84f25284641bbd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf829aa8b7630d812a0a1fbb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33c1f15a08b280775112b0d55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2dfe4b492827d9fc4aa9f79c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47df127c9fe2e9f666ce7b0ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f8daea0de0d20cf6db7cbf8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5299a2a49d1d8ba68e70bd1d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73d43da307bbfeab3410464e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9787a14c347a497fc803827d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf503e83109232d3fb1d01554c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb307aecabedb135d165c33376;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e0eae7f1ca9ee222552e1cf2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f825a97f1ce929489ae1be26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0dcdc1f74739680d64ea601a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dd02e7560d41f23ba2f7f501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6258d3f7a3b351fcf4edca54a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ebeb6d8de4d85645c1cebc4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9183336f02453d658d15830cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha69205c6251bb82cf334ca64f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40b9271c5e92ea9cbeb8b3ce3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd80d603dca7316925eab8f0b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd51818597ec9f68870db58c22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39c8104c88933f5f403f4b723;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16e7e238a78dd55bd6f58e067;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c1b7c0ca2ed28c299a874a84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda10be700ef8c5e533c40e838;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccbf3cf532006bf74048eded7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h536c9b9c9e15f0f63fca021f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9889779254c34bec76821a4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h923f4f21a776842e9f4401b63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4f5851be629e11b6feada80d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ea430c77c8625242ddf1a04e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h224b276a1bfa814669c0cbde0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h241f6d3d0f812c18945941c25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e219100a9e85d88f328f2727;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5eef2b227c00ae8745959f6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0c53cbea2df277dcd703c5d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16a787e11018848806ea56846;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde6ee954a8397c2c8330c4f84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebbcc278330ab9e9a934b5e7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8be5779e5b07faaf9f0587c8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f14e321599f4fcf69c703d7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb246ca20ce9476e0535d0d2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h719ac95c1e0bd61ca3ed7d4dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h618485d3b21fbbad90377097b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha96ab1ddee69bb20f80e9ed5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc81344924d2b959c33c5848b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff7cd58c5552e51d5dc191aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ebe53531becb8702716e54e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7065345db4cac5f2573fcc88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55def66f97475b33f918eeb6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc036b2aed53a63418ddce9a4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95e6791e7512893b252f688dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h473c21d87290d6d0dd7d9c269;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74aded64b2c6ebe2ae69076ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1334f6449ae8374a3e83964c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32da73cb0b5322ee360bc01df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2a338d0ff633276bc38753e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8965d9d83c97d5b0f585af71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8881fceaa9b9df4ee7ec9f6c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd25bbbd9274555ca154c4761a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28502f0db3c39448f16a9d239;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h505039bd820c9c9c0e4c43354;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b8cf9970e27c16f3d61d9665;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfed358b378256457c6adcb40f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84b3352bdb337208bdde86421;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc469111e5b62ab6e886ab620a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3df0bf9511c971af102d9400;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6590cae3a07f5ef2cca53752;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb1595c417e6fce3978eb4c3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadf019518aa145db054297ab9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he02877e37f2f937e7c3c6122c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9348ad154b8dc0c394dbff63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb12ca8c0e2006fef8ff0a63d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7057694ed91f9fb5aaa8f00db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89611c9fbfee9ff247aec63e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a982e3b8a114c1707be4005f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec90453bda866bab0a876eab0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb557d0a17c8a5a478bbfa6095;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2d7b8bfe8c95a0596d421c7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa5405fbc0c2888c52dc0c87f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7409b3c6cd7b68e0dda37ff40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85147238ada3e3727fe7bacdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfafc88c24b05b8695f5b47adc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dc4ac821126925a91c95dee2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6446ba759ec938901bd26e16c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h196394b46a57a2806eedd2700;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82fe848983fcf25d36e35f979;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57fb4c936e5995822769dc4d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2ec2f8384b1eb16eb65140b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha996ecf87eda56a58a14fdbe2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1486eabb28e1e4fbe0463bc8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe4a60c77e8b15e8dd2cdb423;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41c2b54302d37e7ef00a91fc5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc13eb831cfc9756af5fd97a52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedf4a39f0b8988fd4f0d44e48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b9e462ec51f0fcd16fcb9b12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb89de96187077718323f7dc8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c99845584f4162c5f4ec6319;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf12f98729b454ab6f00330893;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fbd99b8eaac0bd027984f5d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1cdadfdeafda1767fcdee662;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha40293a0f0b2238fcaa145ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f6e8c229683f0bc450fc3a30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h579a05108bf00f125a1ef1cd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97b694fdbe9787e49e0f87fcd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h824d38d4352f1116103d3f47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1e22bab07824cca0c66f4677;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb058170e1682781626dd1e362;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a112e830e0818d368869b626;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25b1a471c6cb38e722f586ad8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cd7a20994f73fd7a1ccabf5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hded7129d8f0c0637f4e48883;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5578cdb2e5979b15bcd42c4c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32b1c856d0058d4ab9febf4aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a7b3d95071930867c1a88a94;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88e933392629fcc82d43e44a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb2d674014477be4f68f0679e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc364d451043d0bb072f8aeea2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65b085ddf86436cba333be626;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e7268004e0b597010745ae01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h866b7590c842c1f00276d57c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2466e2359ddb10b3a8a4af8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3efa4c4fa785f8b59cef747ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5afc10bf947385b10d78fb845;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6852cf68fdd26c926a0e043e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2c02364183347b2645c45c37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3594b4a0fcfcd335a0f82e0e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h398de7c9180f7f70fcccd20a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26ebc0f71591e88eac0083c02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1abb5b698b240a0fdff8235e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62d07df0c7d2b7b4062597332;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2ee72d6b5ceb611abb64e33c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h762786ddda5fe5a0755ffc1b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2087224ffd8422b35f6dabb76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcafd3dde303e81e691101aba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf624b3c3adc6a411be89c8b0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7662a82717a00cd5a2d7b08a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he191465ba3b73de9ef1038d83;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20bd9e6ff256a4e9b47a03c4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2614a16046037dd720c802c23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2083812785495f991fcd18ff1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6054cefee35929be4c1a7aa9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf167788e4c4d45cbfa1a41b1d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffc9d56df0c9f46a63b9f238f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ea4ccf5e41025ffaffed72b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb50a93abb78611b122fcda3ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e4f8fdb76fdbccfcfb1aac4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51c5d457d78f70a3263496c69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa5015068c06ab39ce52a8241;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8044c8bd6e417a3483cadf3db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ca97d66a33a2f7b654757e6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he26cc55c85b80ed2c1f8089ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9412bd50d2611ce49d87eb69f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97acec83c38a1986d6af5a6e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf97af536023504517b4c808dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d5320fc8e7fd7b1ca341fdd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h653af7fbaa940d825a3aa4f5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46154a782f53ca18323ba9942;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33943e32eda0ea561014ac217;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb56a854f08741c3044ac1603f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2506b5450dac1d26e0eebe44e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h958146938bf02cc3cc89e944e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19b595ba8edbf2ddc7efc63f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f5b5cf7fb0182d123d3b965e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he07b5d889f198c9674af3cda2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87f09c99ea938aedfc97ece72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76c8a897a04f7ff9c2e10fdf7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd1ffdc012e8634add56b9ac3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15461db7c0db33cbe0b849057;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h222c40fe6c3e0d12278107156;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35eef700f3613c5bd3914dd36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0ef679413cbf2d33f9a3de8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93fcea0ed30adb6c1e116993f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6700a38fe34665139a31e4893;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1cef045b144972ed2ba5ac32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b0498bb1f1e07455a4fce568;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d01c73bb375312278fab7bef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e105664b548f71deb2cde7f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19028fc0f8db47602d7cfc2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf76f27b9161e9e1b0647c8131;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45a3362a5b1e639a84c53e3a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d358b5ce925cde24bfcc3f92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcb1d351e316c671d29c6878c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed6a1342837e93884b7f74fd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c6a1d9aae040a1b289a029b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d1016ddcdf0fa860131de60d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd46e9fe62898b03910908bdb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b891b6986f9e9289b6cd7c99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a431aea8ca197fc103f15fd7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11ad4d0066a21718f8a4cf644;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5b4589456e4dee3b87063f9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d07708f7780ea39a1dc79be9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf646b1a11cbe14e4cbae2aa40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8151af3fb503282950f0175c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h475bc4221a3ee216790c505c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d6b2800cdb64ac004fc8b46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14c26ef098fbaf3455c9c18aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h278ddb213cfb785bb8e857ea7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8e1c730a2e0c9a34bc5a5aa4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59723dbf6c533bf4bc02c5542;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3258a53aa9145260cc5058308;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb596f8bd4a97a9a9c812b8b15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9b7579a0fb52067e7477e39;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97795318f0d751eed1796fa14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1867b7b8f02b6aab8bda8ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee9c4a0303a52961520ef24af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb9c859bb47bd9a53b35a4461;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b1a6a5d85a69492f47d55145;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7ba2737df747d241a1e6d223;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde092d2755990f23a763a6233;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb442c27a814f8a4fb6c1da580;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h363f8e1bfff391ba7ffa9e345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9b9e8b3e8de840b4fcae4555;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d9c575dcdc6de4dfa17bbbc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b2dfa41d7a3763d2dda70668;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h808ded5d889f7a0617b5a114c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dde542615ff8c561fb36d615;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd2dd1d33277e0f6904c36686;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd68e9922acba77490f91ea48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39f3aef0b9bee36de7aa8ff1c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc822b0fe2e2658211e60f358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76538fa359b925c4f4fe1b92d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c7bf8cf462004009e7ccae18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1526ecd8c813baf35df1a9f26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99da294dde1b946fda10a019d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c6d042cabc506a4180d925b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f071f3dcd32452c183b8a804;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8524c7832f6710014d57e45e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66999bddeaf40a4d59e8a4a19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h856e685636fdd701479142880;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ccca8ca2b3117fc005d608d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9639df5e47420bcb9beb38066;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2ff84f82517b153558d8c6b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12ec8470dc40235107608daed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87066950827702f9d6ef87968;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25eadd5ad1f7e50af18c17df0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4616ec3ebe25890e9a50f7872;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h839f344c22b75e23f70756306;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha04ef0ff1199b8a0d86e826c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he13cb61370b7079e02b1764b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f93fe28c0589af631a08c255;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c4ff0f58071d2dd1371edfe7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9e9136e2ba6390bc206c9e55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4548884ae061a3f3c718dd88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha51537e0afcad8044c6030e65;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h734fc1511690600899c909246;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h758d784462f67fa74b25b87e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3a8a664cb03a0d7419b19d86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h639bd8e866b9bd470889fb893;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc405820fd26daa77d6ab5d20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9090db95eb059d63d9155faa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f109cd822b88c2cdb693edb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f448f5427466d6018a3f4801;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae0a9d0b3fe0ed862106ffc01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf92ed3d618bb05d6b7d9e6944;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff7d3af2429c1473193e69074;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d2d3add7747dc09ece7570fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9602d4e0cfc57c56860f6e9af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0a96d568014e8668f9173623;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb15084275376a96c93eef6f88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99baec4731e18e448b49b8b4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1cd9c4ad5910d52dafa433d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e6f8ca1e4cd680bb7c6bcfaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3dbbfc5a81ab3ef9a7f7cf56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2af25ce6b9994a2fe6bc3a9b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h758ffcccd9353ed7e23ece32a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b69bb4f95d9679764dda6934;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e7b4cb73031b9cec6ba17fe9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b370db069d8e5eb1588a2d76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcff4a4a9031ddac285da11d8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94a7ccb9ad64329d08138d02d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef269d5548a2a365fd9d13a46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3413d78e709d12e519ec2c3d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c3e3b22b3c192cfecfa8203f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a49acf5e59f8498549a51254;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1d96644fccdd998f00a9bf82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2e8da7cb4401538ea4fa8b54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h967d2730b32ffdfff1b569e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c9be746e4af7f0683dba1ca2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fb6cd49a061ad56dbf3bec23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf8f59cfa3823194d68ea88bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82d6fb1b10fa4618d1a37c7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef1a87111429421ef2ad69b34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5541af3a7a5859661eac16253;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h486308c08c3363133ef83bf16;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f0748617a75f0f5ff1991aea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcbc3d07457ef678aed2ae48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd41c7f1f50fb1c380023d438;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h120b7b22ddd0be7ca0cd6afa0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7563456f6474aed0b28a76fb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h724c6655b1270a3e6334dcb54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43edce04c451f2fd469e9bf1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7174e237bbbaf9dadeeefd6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7fa424b9fef3c5bb11cc0c75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he05c34eba6d93d68a017aacc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf8d55fa684ed7962b6988966;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fee4ad8cc072c7a04a06a97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h469c15a0680f28cd678e407db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h841b09decbdc9356494085ce2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fe8d83cecfcfca8f66de96ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a9aaec9a76c6993ec62e5fb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8574f3b9ed4256923d0b1a95d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1fda57e71f82b911573c4dd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf5ed0286376bc2d53870570e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13b688a8e6380d4b1bd9dcf40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79a72dcac12a61b389373b76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80ef43a07feed951351999178;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h404aaf7a2a044d62fbf8de12a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71f8a2e02aefaa615e7447beb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha079b4a7f776f2311e4ae68e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h266fa3e32d91a3670d77f1941;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84e468ad9f2cc129c135a6590;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0bb486d14e1ca34788b17acb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56cc344163dce10029849796e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9cbf6fc4e79975f48f806f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha811a73f8f41cf6c41eda38e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h324e8bbb00a4e2ae64e1fcbdb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49f56f8011bd5302d018de8e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bb13f0389166fee002ef9b12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74b7df30896abe49699c8d85c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9677631ab25b4a6567ee1fa8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac32bc9e0b62755f0ec7c45d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f9b6623d847d1e39a78bd2b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ebd4fb021b0c8ee62b8876d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76f3b82471959a2b13b5d0918;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c0f6be249d4150afe6b8492f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53490075997bffa36227990f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d5e9ea024ebd50241ca7775c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0f8ebd24e8603d9c324076dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3e94056547a506c165d0fb7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39b1595d5a4666e3b94f20708;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31c2cf1ff6e96124f11ee5ffb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92dbc2cff7ce6d79f25fa5a9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f01e1ba71e790d32baeffdb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11b4321f870b7d5734ecbbf34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0341204b2a54c8b611cfae42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc414ec233020e9d45c9d0363;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1af250351b1e3895cece34062;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h910bc7433b291ed095490ca0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e19e4e9d3c06a72129413477;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0e4362b4629ca9e6521eda52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15b6813706213d6b019af98a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heca06c44c9af9472a5dfd2829;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb418d31a04303cc7a4c0be01b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccd2b04bb49c455a0cb3ab9e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42fd90b3087fc93c3f755f575;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ac5386b10219ff90f8aa70d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9216749ac77af15d582400f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68baaa211a8bd551f3f33791a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5307608392c602c13bad7c95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eda2fda483c0a20444afe042;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39879c85a3536de8a3163de3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h478bfe92e2d9521e7ce137963;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd70732b734c35e2d7c3a54cd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e362d3718b4ae1a1f94f32ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcf27597bb1a16ef7dd15d48e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d5f909e4a14b92566f3846bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd1b25109dab25db11208821;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfe9750fe78bf68b94ca0518b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h431e40ab1d6312f5936bbf99a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0610a542cedbaacfa82754ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a698f007f7357acad2418cdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee5d4a636de8bb93e40c969f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6227893e3377060c51b90fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5889822de34142608a8d86686;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dd1c4a523f39e1f86f36a909;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he258512cf392632873b6f41d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9b620068ae477af63a77c3c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48e424607184bcd7633e6cdfb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba1060635d5df0104193034d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ad1cb695c4bec1fdca2a9a8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c3a1631e2786bfdab961352c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf31fe02d255811b43cc55f0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd490acf6a6d24067faa0044c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32c6728e7efed91a60accf0d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bb7b6d7f9cb3078972fa5a72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c8c3ad1114b908d8af38148c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda17b421f7e04c40f12a26021;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha248858106d9c61be833c9a41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha921d130a669d3600ddbf41c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3caa64e4d64739cdb43d537ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h289f255ce5dcf8d7014d7cb44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59965fc843bd951f523327097;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4e772fc6f835073d721e35e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6d8dc58238a974f0b6e2a96b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4a83f37611481c7ac8ec30dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f16ab365969f0b495b6c6d03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae67dd2d449a1e5f45f514853;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c8f1a60cf9d070b36dafe983;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e5c45b78b158d42dc95cff3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he37b817a0983eef6154baf2be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc676408636365e76ebe6229d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7fbed5d807fd430a2ec745c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1748d23ca0318d354df01cfd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7aaf635821be2797e7ebe03c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2450e4be6551b576d6de1c26a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43d9cf7ebadbd8151718e167e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb03bc6dbe5a2bd2784c30d534;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha561a1c8a9bd9be10e0510fef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf228c2db313d23ab4a54b6b20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h525d64622a275cd8117779920;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h232d5d7d4548f9936bf32639d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha874f842810fffd4d36bdaa54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2378c03dc6f8f8020cf2f84b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4fe960a39bd3f891f65c20ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h850eee9d01dc844fc01be3e09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2be0be384b61062dc04fcfd43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b6d466e4e8021a50f991b7be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5296065275d683d93a1f0238c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf77100a828c99dd1c3dcf2285;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfac353c29918ec222e03677e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he52df59a716662f5c23e0fcb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4f7f9f3f437efe9b0bbc32c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde7f9ecca85badf31fd4fa2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9905ea70fc1d0e9b8ae6ef25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc984e17a67ec20d8d64ade05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7667f9eaf11f6f050527a1f81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1dd0f05bba5eda3b9810a332;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habc5693d807de7b185f5957cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49c959c6dcbefa24fb024ab60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f2d5094a12c86381179aefee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ffea0d26189c594f97f55d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h669f6348d88036a52ba7df69f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24b3bf396403dd933a897605a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8283217aa483d132ad80f97e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a349027520583f87f581e14e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b9552acc5e551ef618d80e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c384da14f2c536ea3f24f40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h579123dc5de9376c8fe0b5969;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff057dc810c9753e03562d4d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb6fa5500a0d0031bee1d460e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8820d5aa1f405959ac4ea37a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3ea8b302ee7e2e7fed2d27fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4323061802d11f582d69bea4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca54a68b6b52214197e6f8656;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc44145ce22f2d697a85a01991;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92eee6a551282a28bf8d9faf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9f4f2819c0dcfebe96d18436;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3497066b9b83f725e83454f62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadb44c7f73f7810215aecb40b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f5c5dcde2863303690f569d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2da7356d176f6c1472f82d01f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf2208b409214db1535755507;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1e368b589cddef4040bc35f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha13f8c6c22d95726d0598b231;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe549e977d2c5570f78edc22d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77ca446cceb1fcf52019308e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b13ea9fde9680d23d6c2b7bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99c8547907ee00921ec9c135c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6018b47411113947b07b4d1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h745ef43280c0d5b3d117bc8b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a6db96cd90aad98e63c3cc7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h780176d6c6468160adcd1f9dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0a88042718ea22c9bafc29b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9900039e1cd5f4eb5cab465f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb8024fe4d98d40d5730d2b8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c49abb21145a796238fb2663;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53bb45ce78cef0cdce45a2ab1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e61bf08a8463e2f09a78abe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb61b0e71700ad10de1f061956;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha37fcb256f6695631aef98553;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe9061e4f1ae21afa89385490;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15133077aebaf6a6ebdaa580e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h204769088fbf0498ddb2f4c0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heada1e593bb9d0dadc7d874f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf89691da5aea2c12147ada3cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b7837e672ac82ac3c5b1af68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf399de8d98a32250356404bc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c9f874393be7ee84e3ea7ac2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf85073e69022c92a5f27f4049;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac96e0860af8713e5d855b2e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99791c299640b9cf0a386a0d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40c964c2b5ee372f4703b22fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3fc9e7572609eded68f499c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha41ddeaa7544e13d24b3edeee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf78a4f7aeb509e32c5d8067fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5fc4caa698aa53b434c8a2dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62c59d55b1701397de93127f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94275729139ad0ab0d66e6285;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56765a14d2215a033a2beac19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h173b1bb59df7c2c55a4d992b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6be809cbd27cb467c2b4297;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbea331e403e6c7dbd86344984;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7710b19eb18716729aa88007;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbee5365adc98ce322a5527b29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4d9c019e4a2a0d55d028f405;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcc195112ea7d32b6ac422223;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84fc77f36ec4126e38f3d3718;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb34f5e2c4f58d15874f89336;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf780e34c107e3a5c38de01471;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafb9516cdb0654a0fad94341b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc075218bc9cd27cf981547fa3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9240d664d4893f170c3c1a889;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2498262a22d800c8ae6697d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb3f8a634f36559f76af0a363;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcf22564f30a85610d7ef28a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c568ac90aa99e193a7871e64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe4f49b29777ba500fba566c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f3bdfdf897d4edc1f5ea1f2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb28e3a3e6068d5413d333c8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89249ba46b70ea33e65218043;
        #1
        $finish();
    end
endmodule
