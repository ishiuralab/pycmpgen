module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [29:0] src31;
    reg [28:0] src32;
    reg [27:0] src33;
    reg [26:0] src34;
    reg [25:0] src35;
    reg [24:0] src36;
    reg [23:0] src37;
    reg [22:0] src38;
    reg [21:0] src39;
    reg [20:0] src40;
    reg [19:0] src41;
    reg [18:0] src42;
    reg [17:0] src43;
    reg [16:0] src44;
    reg [15:0] src45;
    reg [14:0] src46;
    reg [13:0] src47;
    reg [12:0] src48;
    reg [11:0] src49;
    reg [10:0] src50;
    reg [9:0] src51;
    reg [8:0] src52;
    reg [7:0] src53;
    reg [6:0] src54;
    reg [5:0] src55;
    reg [4:0] src56;
    reg [3:0] src57;
    reg [2:0] src58;
    reg [1:0] src59;
    reg [0:0] src60;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [61:0] srcsum;
    wire [61:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3])<<57) + ((src58[0] + src58[1] + src58[2])<<58) + ((src59[0] + src59[1])<<59) + ((src60[0])<<60);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fa2d6f40f2af4833832f03e3c4b556202395360ccf1c81cf6e13abd52378e3e8825de6c1afffb39cf71efc570abfde00723ae0fefb0318e2d146dd0ad029ab9997cb87a8ba39a30ba0ff72bb59a9b01fe8b99bd296219135e79a828de4ccf6204ee869eaa6139f92c8a31af93bdfe4e3674670517f80a36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a36144fdbb81366424f7706fea7a3a23f2b3064d6a3c7df9ad1795a42379519a5db42b71158ffe03462a6cc00acc3f58486341148454850d34a298a0b803c8564ed3f44d130f012504743308bdc27ba3003e4f29e4a05176936fb3b15b54e77119eb44f627ad4fdf20a9413b53a974b34bfa42453ca2b243;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h675147654c4d01dd796aa4a256f4226f464a996d347410456c296a763279ff4f6ba735d0ba6dc433724a02b8b98b64bed9a28321c8c287c439ba9ce7edc8fa3023ab2895a493b2b4a8f09c1512290bb3fcb37bbb9163d21ca3626cabfabbcd896a8007c778581b02af933422886d881dd628d269a4dcb4db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d3d3678709bd9595fced34bc260c779e69a50084f85152b9e6710cf154218ce8179d83a585b83598fe3e5d7a6d93c2d000b379ddc8ea3200fbd7164bda02fd50af86dc782edd4a149d090e61e000629192c4736b58da15114cc64c5e33d9d54c7f931389a73232e22067930c6687464f10c359c3f84b3da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe01e49a90dfdb5777dce55c437ae03e39861c5d3fdf9fa515036e0cec205b5d85e4a7b417dc190fa28ec7a860ba468be4837bb944804953ae25a46d9a8ae2cfd0c12cc16d1da6101d95917a344c83e16b39dcb3ab7cfbb2ba7073b1fe0d8f83aa472deb03b3a4011b38bf2fc9fb3ce7861b2fa7a38b9914;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bb6abffacfd913aec26db49e2c7e11d115972fe5a521eb344097fb8a926a913c425bb084fcf11ebe989c6fe6cf605464916c84495fbd270efe1f7a4b763f5f2c71e105c9d232bd0a063a3a7612f6a1151d4b391924ac643eedc762fcaed1f323a7f318b2d89284cea7f98a04fa2fd709a1b380c2ca61734;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfefb573369d5bf2e02c96450581ca0c162aa41ace7e2cd78c696dd468d68911da0fab6d0cca56e2048d788a33fc1b6025cb410ee5282488351cc923972ba6b5d8b4e39a1f1f7c62ed13506a967f778e8571bcbfe73baacb6e2ee31d2fe2659a66c443a1c5dce7663d7c0ecd0b2e018cae42ac5bdf47a8ad7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54e3ded708d4a2e6205742b75bd466bcadf562d99c761e9b6490ad3756b39056c54e7fb435edcaf37dff2e054f01d4b2fe7d25afe702a07eb0fb983ec3b20e19e453aafeb56d566af9244fae2b2ae043a9b239aa3d4b401c44f3c7e702c7e4d80517e379c6f79b3ee7e1ff12b7b118fda3f4b02e453a4d49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ba46c4cdbc0bbcc6faca3283a36fc086aa86a893b6d8b357cb737b1b45a5d446bdb1af8d7e48980f20ac2218b6dc2171155282170b23357942a5ceac0088327d90f67683f6c6bebc78db4b83451da74dd2163eb0421e81dc08fbbaf08a0546acaa8e15e33a11e2175dafd82912bc45dd403a26f34219d9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f8cbdf50d3c575edd1badbfb2cb60df4c3fb8de00cb8c458992bfeb50773b2fae7ac26ea4bda558b61143391598806dfae2c0d1e224850481ca1abe5e4ee8863c82a6f090741bdde82f611f7617dca46d84818e84610d8962e839259c2502b6e818a274b02a015a06b9191ef35c36ec7cfe089b6e2a51f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b14c92bad33a9f53a7ff98283d1fea43261fffd72e7f7a498cf01dd3d3579e4d58e40e74a5cfe8a85b8032e88d217775d63838a0c4510f1d2aabba759df6d81ff0c27ae525ee0bf4022ddc30e242247f873c1249e0cf81024061d393f8486a54a0bd03dd1dae1cbf404e1508371654460baad9eab2d8416;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25a2d6edc572b169b5a866936d4d441c40803e3c4e772bfaf7a1de320d752398892d2c73badabcfd6b8948f5d9d62ceec7ed14d8783f88abf95f4e498aaf8b2f241aa60c3b732761939f4a2612de29deb66a00e402c5b5cf72e060749bdd577b4f65d1051023b02ee4341e4ec63582459ab18e8e019c3908;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119eaf78442116b307663c0528eeb71489123b1287c8d5c12601d8b4e1ec64943379c22e42d00480aebed4b75dd605a16f3c4e99348dba31e8c4471e15513d4a0bdcf51cb21eae976e53a90a61fabe1185969b34ae65b2abebf0059b6f6f087966b25da2643a6e23eecab929cb1422e8b8c1329b8e2d80feb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc9b47d5e256ad1f635455d59817256d8cfd8aefd9e0f0409b737646a2e2f226adbea8f58907dc4c9f4d8f81f051f282945bedffb90891da5c5cdd88712d42c55c00e25a9b1c8a4dbf9ac75877eccc05b10c427c8afa940437a9875ae1b36aaa74652ea6d82ee050a4ac86da022f8075817aeb7dcfdbc852;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d064d810057a97ebe21fed3a8bcaa03cacd8a614e02c857c8734c902eb52714fd364dddb5ad2fe3ab42f165b2c1477fe0d667e2b248761746b3310c34e1547ee821f5e8ac8d7e72089e3b494aeacae888cb5cdb089960c8feb312e8811b464f66db78e1fa6cabbf1e8fe79910a0d2943a1092d689c38cbf7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bca2435e4431671bd971fea81ddb8bd07a37a7165951cdaae6b4e5a9606bebcc7b613d7b133db533f9b2a76eadad1c5d859b7d7f9568c0c321e3428a69e80aa531b93d990880bcbc07c109fa188ab38bd12d922b0c6e062879d9c72687d699786263349cbbb969c743570d5bee47e84bffa298a95b6e7be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf397b4064538038ea1be0eef8340257656dd5b4b12928836ba9f220a213a231c489ae591607cbb76d35253b11f36ab1b18942ce5e57e0d61682805530637be26c78670b58240d5133d46ec9db13fb961410098344ca40a4d12b65e0391bd2fad2a8687bdef9e6747a12be819b2c1900b2adc085aff53ede0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7856bb4d5b00abc4129d62e062a21ba2a7ad298f28f9b20ccb7c39bd46be3198199255a74c2c2af1cb6800b2b992ad7c7ec243561ea5a19ec732e7adc720e696e0ba306b205bf761e3a1da16c730e073c9533fc6083b73d1a1501885cf5dc033189713b668d1ac26d5110f0d61901884948ae89b57786de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc534c5765279f4d339e1b66024dbdc072160f3b04146c82ae9f773bc73eb7d92170d50419c145c4debdcb877d43c5627d8cac1ce4de27da190b9877f21ecb84966f1ba9ab2a046157ff6521d0ac15f9a98248596a5ad4489e762724bec840e114c2cba5149e52b2abec354404a92a847247e512f202e3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a899e75dfc764345e580f85d5c09788063a1458d0a003f5d6538f7e8e3cdd1579dfbff015248c56bf4594fe349f52646af9903cd42c0952c7463182911082206317deeeb52a64cacf02193dc366a466dae89c0cf35d961a3de55cedd4b2d2cca9fded96bdda198cac5cda5ec63e23bfbff0d8506edd6355;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c2b22507730e5fb3d990b14e9ebd40a38d5ca759c1b451c9fa79d46efe8a12e2a6d1e5bf27b3b8d71865edaf26ddcd0a9a9bf47386a25303a19393353817583571f880de3df05b2a7cab91759dd4405d89f71b07178fb9e5598b3da3195310f9caff9b015e638858468c47e8839aa75058d0b55d494002b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2d87314b9ac5c5d5c74a7113313befaacf43afb323ee03ce31c5c010903ce3ac75493d9a44ac34cce81b576622bde33d996ba7ba1b8432d55810d1b18d32408c445308a407e30d3d7ff1490d4b635f8ad4251f8540f0a77aec0872cfcb26ec456a3ca61fd3773ba83ee8e69c6860497df914a3d63973453;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17236c7f1385f7b11e94167f281b4bec2088065e7ee1247b89ce11ca1ad0c0fbbb1ea78e54beaf7707dbd090a33287c62d2901a2631b3bf1cebf144c86d0b1e42ea88c960e9d2e163d6b28054563bc98384b7326d55caa835f887d4da259eecde0739de168cee34580652581fa140eb19d492101011d83b9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8bd78a1f5d93f2211807b447e1413409954f7fec1988ef45db660fa59f37109b947bc8ec90422c436cdf30d3252763f71732d51c87f9730ac3886db6b0dffcc765d04e4af2ab535ecf7405e052ea25a5ce5ccb38c0b10c603da214850f2f4d9c82930456c3272d828f7385db0741f768eafb532d1b2f104;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3936ce34d8eccd202bacfab7cb2c90211ecb73ca8e102d771815c4cb1f664ddbdbb6ff2a10b4214b1fa7738bcb3a327db72707aa427fb9fb0fd4c8b0b8ed77561a85d0d94b98482283f03e37e52616aebfa4a03fd15e0ee51b582da311d835752b811b7b577aff7ca4f4f2c68d1ec4cb47d54bbea0f7205;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d699e33afbf0d587541c8d5b98c8a2d5bf0e8d0510fd8d4b47595294824b13513279d0225d875cf0d023e3a9d7c64cabd00d96ca87714d5f3688cd549dfb3d8f15aff7d38132adac1cccf43124664c412e77aba9a3501900c96a63affaccdc4ccbf022fc6a091a10da3e8697744610a0b60317cbeca4329;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0f47da862bd3fa3a0d6cda25a696d940715621b2a8e3595578af1cd7ac97a754ecf8adb037ba8fd898e52effd95b063aa5439ebf7e5c2df29b10d6960045794860a7f5ba1cbeb36481d4a478550ce75931de02b6e40583de2764ff7564782c956bbc131403189e09ad4f937e0eda3ee6d8d1015079c86e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f36e81cefd73efc81cbb4a56dee24c694d0c6863597f86171a831ee3212173a0742a3aac084101826252105eab3e76481724460bae2e52c11edad661dec49c701e14c8ce281e1361c3355e5d912e0f599e7a982b81068f075c0e5e242b37e51164e9f1bf73cf41114cfa81b0db76c32703bd50b8d7b5188;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95d9aecca727d8887e4f9841677741c9b581bfa13d35b8017ac3b5faa7de3a50085e610b873145b6bc1be8a485c03647fcfe02a8eec19a94d72fc933e119dfcf4406a826330a7f788d1e8eb964033e96130ac0986b09578737c20117e9df2f82328077efbd4482839c8fe46a633427f6cbb5b0ac6619675c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ec37031766f22ce59a27f8b233071f6cf25db8bfe0684161218b3004619178a38221a5df7887a96d9181705f95c755fb73935ed9447de7868e8b1b45d80566985da0721bbd36a74aec4f7eaf8443fdf2880baa7f2f4a6b02eae7ce937c77a5fa3eb98b62ee1539bcff2bd5edb48671f4ffd72294663b9fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h801f4c93695bf8d368db9a4960e4e78d4364dc1d43c590fa4cbc67f90c79ca4929523b054ed787f32b20d7d51e27425e4547d288bcd1452e74f45d99cdf78e4699311783d516f1f5f37b85665410a588b0bc727077a36e6d8f7e29d11e45eb8f1bc9393bbd1a9bc7e37e6149e1127db9d1ba9eaad71c4025;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b04664332ebee81ae48fa78e51d7ce83c1ecf2f403f62d7b7c9c58c3cd7948d542364febd1786d0c7b32df55691b286ce20dda0e3da8da8f16c02d3121bf44bff32307729b197ebdaad9f51c36ceaf602d6fc3788ff0c61efe7ae3ec30336225107a04ce8a0ffc1b8841a6cf6a2705c049926c2d121c6c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19aa21414cede2241cd59b0bbacaa4db8b3d60d6cd7ead401e5d8f464a1a97c0b57141fce1c93325846f81733242b68f87ce1ee1a0e87a9c8ca477b8c33d7b225e788cccfe7660a19546cc54b22357f684d93cf728447e776e3d919a6f90311213a86d6ebac311b0827c80a683ed73d3eac0b100de9ccf648;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f94c37d1e724057d6c11770db0a19098d61c5ad708e33a4c8beb739a929cc3b501f256d841a3362297223ef61335c7b5200d4b5aa094d57f7d4701fe223c5579d688791e958ea083e9ad975cb4f4fed8bd46305c958719a5df5155841021366d168a362e49c509fbec7b1771469238bcf77f4497b87fe31f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7eafef4aa468fe10299cca2b76a2cd8f3ccace94f4ee638c3f1df91abdb4acccc471cf78ea5c6f2fa742e08268f2e1bae123627f806605d2713b7c5c0dae66eea21294b0b63452ccfc8a3e97c0f77bd205096f254d1162e63f0e4c95d28d85c19ad8f99ef09886f291e2514704d45b995dd413bb8fe16b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h736da13a6d610cf93f2d14db325f177819b41d5ee9458caf59f688bbfc46c0e68ef88e5bb90f2ca6bd36e36f6ca6b9870abd5166cebd8c80c82515c53e3ed054460233008c33d0748a6b8b374b4052dfa59f911907b6c24d74cb2f13535158069f48385d9d3cc6db16ee845d8355e967b97b320335fd835c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1214a3c7209844b945df8d682b589c364e833899910c793f3342e42f38e7c9001175d007be829c425c4b8e594b17b8dddb8b74c56c6878de70b25bd7c79afb7dc879d26294e03414e6ad4cfa619f20c98bdcc75326d18906fa941d3e01b406edead0f102ac471ef7e8179d11f76759599f79d039248a09f34;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12266822a54a5f5cc3c8cd1c72db8a8b1b85d8e19d78585f02f0d2f204d10e726e4d93ba6f039b0fe97efd55f14294f443fa2d31850d8df0003683aabba26261bd6fa54201315d4e10064b7a0ebd3927dcdf1c0b39a243a23a84bd5627f564fd36e5e652bcc82c758bd3f4d9cdef7b9881f3ae4a0746c1c2c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79bd69820bc70a22dc3ec8f27575415f23d9e9540c77286e2bc19353452b3e53f029782cb85ff34d7092ab1a05750ef7fe8c1e9210f82697f76bffd507e8daea804ba68673d2345093b61afdbd0ac014abc7b8d8ed2f56e69ef14c74be27922d3c44aab50d17740c150567bf8af07f208b9f62888d85a338;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf07582dd910acc4037ca61bebaf0624e028a8f97f5a822bc4cc5d7a45c265020de92496c176c2a878d21ad929a093236ba8aa30db2b10cb455e4e5d8a99fd4ff459d438681d8752f8e80045b0abbdac09986b09cc5b9c124b5160f315761d525d78e67ec54ebced4bfa0f817d3e65aaeef4fdac4ca1161e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50a116d4b5a6d1c6685447dfc52adf85335a01ae2e7e015ff3ebdec100d44547f1c23675394ea67fd252383f21649264113aa845963d7ed7a396b9e0d2237baba4c3ae18cd5006eec34a7cde23477987f4797e4c54689f8b5f18f6cc1359c511c4a78a1fe2ab0150d4c2ca0c88f0a7aa3870f074aa3a5161;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f03a89d9095777284e181772dd88e6b4228bcfbae2cb195836f051972dce0683bd0e9b388e3696b8d3c5fb3d4fa72b035496a58ae35c98363346a31653d07cdadf307a419a9219772d69ec8968eeaf981d38971faceac2a1df14cb0fabd05a0fdd463c989f119200089d4053212155a6e95b7f3c09743397;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16814334dc1fc3c189e9383a57e58de512c2a6873f46ee3abee29fcd305462e727a4296ce05d2caa418250245c973bc3219f012a6a2c4b5fa9ad9f8a2b3114e9072524de7d35d1131f43b8f32d156381a7a06002b8d4e4b0b760fbba0a290bc056cde7d671d166fcefdc1b8da5d7fe5bb829f5f6391fbf734;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7930ea91ccc64db9d89888010faf9ba81a2066020507042d3006e3acebca1a1cf188b20c84db1e0d618b4037a5be6158404adeb224effe428a886f6894099f1c1fa9501a37f9aacba013eb2a45d1333b86d9e1de76eaf301af3ae48241d7b07513c9562e0d131d734d28f7cee58d042589ccd16635b93a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c2c8ae4474a1213e4ee19c7ced29840ca03e88c09b20e2583bf9cec00204222ecd5f5994968de746e766fb737fcea511dafb28e475cea62fee704e437cdaa69ab0f97e00dd0d2274965a2b3813302b3d0c917371bf5fd2d545ba0e8acb616aa96f3a97a5a36bfb292d03fc640ee2b5e6d1b3f2da1b26c90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17012cf28b2902336042aad0a0f117ccc9ca281400e7ccb248ec5dd7ce3744f0c44282034e74d1c356cc0f549fd702e4bfbcc30c93807c23127fc693b35b98590ee80d8d7aeddabfb98cdba3b3de01211f788602d3fa93eb1ab096c183bda2f59be6cb1c17ebdcf0258d4ad2d491bfcf89cb56d706ee3b0a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85f65521d5431317b6c24791ef7b457a9bc2375ecea4c6f54a46b649226efecf67a3d701198cd5b0c8409b62f906f04d585a464924125c5e34884c0cee65475886fa2e875de07ebb2f546351423b43c30b943c666af30171a47b2989872627085c915323cca028e9cdef12bf2fe0b9aad05344ac8415094a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d2b5bbb9e643651a979365bb5d076b65e85c86244aaf1d692a3be96181c6205b5e3231e57448696011db1f19e41228f2ba91e18a61811d54da5db65878e036b473e5dd5fe01e8aa39259721423dd10fb3c12e8e805de8f328aeb20eb1ebb5d03396af8b499a28ea79cee569f5cdde88b792863e3d172c7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5029bf2f47eef06b1266d9902962abd12baf2ea344c3424c4514df19ac7c77db4d77e3ba54d9f5ae5ef6427fa71385228b66347bb18c1065a219afac52ad2edbc04369012961ef8d53bd9ee63de087a74f8359647771c42a93084f7580fa7b748315c0b0e7b8451f6a86310e3229fe197a03fc067c39126;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5907fbb5bc52ab7410e7dd342362b358f473fd9f9cc1585dacf13fbc0a35e56a6b8d074d3c687c68254d7f3f2ed995412a911cc221f3269a0c3ad48be237e63e0235ef5fcc77e5d6f5141ea697505b169af902be44f9b83e782c9e434c1ba608ce6b8897f610ef91b308a5c52b9ca61c1ae9e3dd4dcd8db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2082a55afc273cac89f649c5830252a944eed54236351370df8ac297af17d652d955ee0cb6204777c3969b88f735f176234e593e50a8625393c725ecc9270d8aaf5c8960517f118bd84a6c377b768ddbb7c106309716c964a0f1099ed3b6a116e9004ee8b10527fb7f25a32d91cb121c1f27d6d64abace7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168cc6b92d2297b8dcc9baae88d949b42ca132b7b111610fa2cd38bfccc80fe05e87107e3545d87ea0c3cd24aa59a9b675585907a21d2876617e7b567cbaf6324af087e66a59d27805c0e26a18f11ea5e9045fab9fc9d1061f97175657a9fe69e26df440b9a44d1b1e73433899ea9349d05d1ba02db91560f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153d3c788ed5b23e16c4d4d468c8cdc3dbdaf8a75bf572df91bda36348a0c0e2450f9493d5ad1970538c92cbd35b34f0c8443c7faec21df3e23a54d34337b33ecbfce449645c0b74588b1dd5b6a098c06e5db885007ccb6cf6c8a49761df9274af891d43c96d9de89c0c2d3dda7406d80e3e316e0548dec02;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18620ed3c62432ddbce3802a9c58b7417c9dd25ff5ced3523f3ebb9f30053d358c2193dbdf91f68d38636b3caa96c60b4dbf91052666a488bbdd06dab0369bcf3aa0e2cf7a624bdfd990818f3e04dd4a47918f17166e50a0eee5a267db31b97decb0dd82953901ff8090b76de4a3bee11c4d24edb0647b697;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d68ba73c6ba9d766bb5372d2ed019cdc1349cea2e6aa0504acd596bacb1f5f32e2da15cb16279fb1f97df483f7f176c01f7de33597869ac451087d62abd95a1617e271b2a2fc4ff12ed1a4abfd76b5bd529ff6ae9234a7389311e6f5bee174fa55e21d50f6cf4906b0f51cdd672fde14f2c375c48df26ad4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4ef521a2f2f2430cab8e100d9dd971110032755bde9a4d50e1f72374363a448411d00ee3bbf27f00b43d9f5ccf395a0d8c71ac3545cdae3a3037db8dddacfb06095f38d671944ef7333217c74254ca859a3434cd7ee4c6daa5759d45f8ab7213fb9cfbde3040053e311f1e7dc0d4363b0711b5e56018a9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10590e8325480d187a132c4958433e5bcf02bfad28bcc3208825b6441ceb205c5683f127d5104b09c49c59cfef3853fa71054779b1f6a4fdf46028e56f358a0499ae22a212e7de4c8990a787f83ace8952084eb2115d9044ac91928ea1b36002bd6b83578185a14aeb7657e9838d31946a3127449a6e7cd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda5488384a3e63db112a62ab076f5358bc72b6897b01b4e0fc19e3e5c0f908a856dd0456d4697a6c1365b74507cd292c157fe916bb0bebdef48fe23a66c6b52164a157885f98f6ee41c9ac948045d34222e628a1dcdba3aabc43e01a4fde0ef1711a5cbe81d3d704379fe900335d2165f060e9d94c990307;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee819962d9df0c104574064eefea7b9bf9f3dd68d95e30932b5c3292ebaa0c0db6887082603d133236984bff8dd919c4ec713efac56ed14727ae0dfac1c0761482d664e565185a6b3346e5dd8b9590489af87e74487119ebf1c02fa361402cc1aaa8add0f536f3cb58214cd687285f6e508e7ef9779f9977;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb1931a69517e9fbc029b8ea274761171ae1d2265fffd277ee032b6cba71881bc372bf8b6933f29127255b0d090f7425e41b7254cf390eccbb6dd6e6c01bd6c4a8c03f5c14dc984ab425d944604009d855242f3eebee2e669fe1b3c0b9d0871ce2db3f558abff90f8ad27da4c66f811ac8d74ffb0974fb21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125ca60f72b298cd73668d4598e52e998ec29a6b4d9569c42c27c9cd66a1861c42345a85494eb2f75d74f9c5f7fa5f682ba98706f38299c8544045531dfa883e458574d2b196b721c82c3e3831cf16819d43dd441447ff9d2f2f1036cd23d65f159bd6d8e99f4555bba0f478f3806f0b528a3eeacf4e7628c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8211d82eca805ee76171ffc1a9716dd72c51772d397b1beda6a73bd20b887a857a450ecf9bcffc6bdff74bccf57c5ed7ce6f5cd6e72b9965a92da24da5e5d09fdefe5e8a097449cf21c4537d1b6ac68e75e1dca9d76e7db26ad5eb527a4faebd2613417bb874a06d4d72612f69937d0b9fe26e0b7e7fc36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12239e51a5663a939df4fdce86b7ba9174ed6e3343c0a8335517a0eb887506d11c1447e9c4b989e74e92a5c23e1d6136c53ea6f3e39bf97387ca19e5031ee76408a0d4229bc9b7eeae6cb3ebb316051e66e3e65855b9d7653934c7ba0854041133e92d06a6c53220516c158844e51b5cd1e6394a66cdf8054;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a48b94a0fb3ddfa6d3a622e4c22c2568989f14c0b7b2d026df3b7b73394ed6e0706c516671a1c6557f49da3e1401e6333f9a48c7bc2b1fd9d80e4fbabd8076bbd150544f34fcf9e4c98b8c7b65a4dc3fc77a570daae0bbc6646def3bd851f69b1c9a1f8c774b45f0eb1357db299946b2def45c5b39ce84c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c0929302443b81780d170f1db657f1d4867725c4bbc53486d4cd65ae24a16f795f3622635f8aec60a82bcb75ae593e300a3177e4d8a3c540907c93ced61a216dd9f15156b2cc0ce76e241b8dd1446e6a36fdf22be97e4960d952f447749985cfe5587a5879d8681d017e99e8447af7edfefc38316450165;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9b6dc915801b8861faae90efe177dc0af0651aec4878289c5b23c85835a1d6d3d4fb4c252aa1a63480ebc482af71bb5eedc1ffc3bdb26c1bae6ca4088b95468b5a80e19d01508cd7073df9fbe1ef816e9839b42db9f9d95f78241dafd07309d597f3eb35fb3b33da36c56127398946fbf40236447d21d6a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b96f02c9b0dc781b43a1e5ccf809ea0d3bf1aa4fbde4fc25ec839d5c16f7242563d283cf55f041b5ad4b3a34c1a7b8a14a29555e0f64490b0c25e93037d1db5c2d6c05dccacea08b860abff8dd0a2b710edeab162312983de1bc04260aed00157da4a60a5c648d95b78647825a0db48b6f4c8905fa25991;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4a33d8f44366ca1ff6b6d859d8c01aca9cd3fb6100ac0c82c9771362eae00302809a4964c2be1c81e84646780c8e8609c75dca13563d678d278919a5bcd97ea45c7ebf7d5095af9c48e436bf4ba4599fc711e4be078819cc17aaced0f83962af1ec9ea51cce3d72868a138d1204ed00e3d03360224a64b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1191b376c9d1a9aeb6d02e819ed0a0cbc93cd70136739922f9e10fff86aa13eaaefe09c4a5db30b9c84a34b6ecaf245f3f0444ed3cc8f1280b4b81ded34ee3c4b711003a00e92e6caed869f8fbaa98edc15086bc6ad8dc97d7a41a25ef663a69db67db0bebd7edfa3e7068073f096765f44fd04f00b5c2c13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aab170f928a6812766f4a3a10af69073e6f139fbad384992d5c5da7e912456a509c988b30280909dec5dad21109bf7ab4e8e54adda6d865e16b110a45df90450544ecb63270aa352325dec9a5adcf77c1b2becefba14e22baa2de648584dc6dbbb9464c991f45b608dd43278e071d9d61890683131521f85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17edf88407f973da2750a5c4102a31735fdbabb87ac83f2a8f811ceed30e3e164af502688054a02b2e3d16c191e94b1d288a6cc6f90421e2a3b36337793d8e0f8ac172915aa645234da2e4d2e16fdd21cf03954fc95d080794e4cc50e899e456dc177e6514d34dfb957034ee8a141bf083e953eb9af557f51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f18a5f0fe17a716ed8d2a49b5a781e334c594d29c07f9362342fca5199b7331d69072b6d1c2ea197cfe49dfc9d54062949a113fca68031d39459cb8aa0253c48c17072620db09818887da0d2ae92f9d125bf2aca271f0d749841d9179b13ef2b4dfd2c14bb1ea50037613fa85c1b07ac2f77474bec22f6e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1501eb3c086afc766ef5ab7f72c25adcc049e0d3ab113d59a545152d565b53e5efd42fe5331707d5976ce23f49b65d5d1af0f529cf8a2e4c89d8e4f3ccbdd916ffff010a4f3ebf328c66055460367357aa57735bbee700da5c4283499780b34ebfc7f90571efdc994260901595d9ffa18557b501500d117e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcbe18424cb260949400335f6e63b1c61df365a2c0c798c93c70d295296f88d030e2b51b9b97a47629ad087ddaf56fd66a4c0cfe30742f2809453114cb00b6745f9581df6eb7c9c6b14b65ed54dcdc2749116c7bbe3506c0f53ac0829fb39b1c5f563b6d018efb2c962fcd360a61864f166e7daa6942bc06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c34f5b0618d053689bdae066fe661eee54fce095331843c262a103165a46a89dadb18065f521be6625eb0d1dfe476e7b2605f0e66fb4a9be9de49f70dc050a82af0dc6064176962ad2d74b3563ed296cb10fb22e8dfbdb707bebe142df920cf30609ab962b1b4abb913f0ff0e67be1fbce6086ad9eb376dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17362bc6b6713a60fcaaa9031a6cb8fc0bbc82a8b0d0cf48e9ce9e94ec057047bb0d5b0a27acb2e37c1f2eaf33cb695d505139a3e45a5e742079b6fece3df65bd8881552b34592b790f35e9ba971e349d2ef917c364a1058a61253ed843684a0e8cd5493647c500f1d13d7116afd723a9c490a435598e9ba2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd283e65cfe34424ceb9385b25a09b29566506d9b93f85bc22234b211b909b9820a150ea9e6f3c47d071e1229986458b499f103f905e428083b19e309d6f8295ef3f195e3f788fcc21f38f05b4ce6267d416fa96b8126aaa6c3abeee9d3e6e7afdaf263b178a0f4690b17770d149fcdd1a65bc724dfea2865;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afeb431adda3d60e9d0f8729a14db070fbcb6a3821ee341d713b0c992b4470c08143d10a97f2e6b54ff5ebfad3d3c55566709cba76d15caaf9a2b5e9420c1c918e29c3281b021f4c1d899a91e730f894b1892cce0a38262b3057e8e3751abe0c7883e02682f6d7f3a288037adb11a37eebda5757b21eed55;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15572a231660a6e8e3e748dccae2f08996ebcac712b5cfacfe5d09c5d90b02e12d2768579f4a8506b2d3edfd9420452b90660f52b9632790c8086618c4b075e4332280c14bb47d0bff08c53afc72878e4fe165e1bcd9285da431a67b970df67e36b71e24b0c99544fbf3524993413abcf69c9995dcac001a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26eafcab0f2fa5fc70f235e4103af23d9afd7b865e0eca07e23c7b2a1e54bd1219b9036a8f42d20b29973a30a68c0a0115c28eaf6a6840062be3310db25edeb691fb8e95f46770312bb9e9d66fca912a4754762fbdb0cface7ef8550dcb0d80b5d63c6d3dd9b15eb31a4982975982c8b513cc0fd0e987a20;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16551695b8c07c504be21364c951103a3107880c00450beaf20701f468a72be800ef0d35846eed3a5cb71e5eb0bc36a5f7091bc5a9d76df7a28c0f405e90b85e22f7a8b00ae6e8504f776f68902afce134fb15ab5e27ed7db2d20f0b2acf2ceb23c651c45fab6b802b37c1bdbc447e6d2989fc18912609d5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109ae3da0043f712e033fbdef4296caaf00c05676bc9b35697216acb6387f310e92922b0f0e74cc973ca344ce537708434bb7c885061dbd7033ddc3e597487810ee20a24b8c8110d84ea95ebba4bf006b5a6c94d7ac5a82399f79eb3e25873d9d081fc514607b53e3c8ae5174c4cc6ab27120eb42602f70fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9806766144762b1807dcd4136eafec17b89447c9ac9f477e6a6e71038dba1225f364fd6cc10ef7fab5b67185d5aa8896c4fde11d8494168d043cdecb07acf43bc8ac1640f34bfca632302c8e9bbbd33c43b02596c5ecacfeb22f242d073297c5a049e6c3085e0c5546fd2f0619c3f07a52e5e456807f83a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16153133b21e3a47c7ab278e6de1f9113677b4a865c168c6a9d90a378df161f5a9e6c4503a29e37c2c9337e07af8cc326be5535b571e5109ff878f532c37a6e2eac1019900da134fb76675d94f9244848b06654c869f104b58f2977cf893dde706d2c92f282d357c9663cfba8d64d4c1c221b488efdbe5bae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8351c3cc514963796e993558bf86f883ef1ebaeac0463a529d434dc0fb303a9db95a3403b58917c7416ba8a45c2abf17b4b138e73dfbff3fa7ab5810f166ff1f4dd951eec06f4d626f281d3c8c1d9b78563ec6e5c3184c47352da6be0b45e676283b82456356301012a7ead71239cad8d777c9b4dd0dc91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fca59818f95454f2bbd1be335fdf7a0ba8b2c62e59f3ea4faa37580d239b93e0fb188d3d3ca0d00ed9c22fa2455d7cb9588339639b6c2804e273dd48009c0cec319444e38a868d9f5707819aeb5e8f7e9d91a160569b006cf04159737dd7c9a594460648f09ee4c2c330b6d8fa6ddac4650a90f88b8b9f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f1b3694e5f26427abac2f28bffe5a92b3783b4dbe34565b607bca0f5063f63879ec263b586c61727e415d73bc471a56e7e69367033d913e0a7dabf89176270772ca9cef219306920d14a2ccd27e04661af729fa20617c2a62ff95cfc31605bb7834e2b5c06c50f512e058da7e6ca96b5ef3aec7211f844a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d67cf27b8e8bf8477f730f69c96604607a9982134a0b0b50b0bd8fb229eb726abf930f455a9eb31bb69e26b9c418776480077c261692815b346520e986273895cef10243e182ac96488a24415912cd80097259594e595935ac36df05d7fe2d7653d12d81a07ff7754b1d594bfd57bd2305bc48afe4cfd52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3636efc6fbb245d587a51ad0410f5974298db0190459e2614133b699e7c254846c947d245c7720c7b144967511c09cdb1a7d59b9dfc48d83596b9f5da0235efdd70d638cbc4b98332d2d4b71248edfc4d1ebe64e75f8b33bc03b144db0c50536a635d39d1c4b346de512724b8aa3122d37ebe237592e5d6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3feb38ed64b7d2932c4db0eaa9e85baff9b3387beac475ce01c787a051f7863f0cf9d50f68b9d1d7bdcbb5c2b775bbc0dded792895f0369eb82fd2d1a74d4e84084a9e059dda0e40b5666fed89babf8d0864ee3e6670398dfd3ecf85129fc9e3a273c168ae1c30204c26f7ec985d1253d238f78cc979ff7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19347e8451bc9230af0858390f06eca227cafeca04cabd2140a4730f91365f8a8446e79424d4e73d9256a277a639bc02c6a65ba0ec523b0a3451481c7dc64ac5185639967a4d7577605db1a7b626f107409c08de7e6478602d081b11d2d60f43f8a1e2cb08bd40398c7f5726a4103e6d29f4675a81622bdda;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d84dba326a14cb4fbb8e40610f1b097b35a8c0969f82c3da87df111475cfbcbe66a026deed6a2b50507b4a44b12c6a0aeb203852cfac258cd24cde158e6ad025fb7a0e1c38db974b40bebfacceb75d662710ad7f79618d5197bb495896578117e92b8a2a5c2d70295d9dc3b518e25980931ad0a452de0f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9427e57a2aa82878ac6a8e46131afda54b14e721bfabef32be2856b38a5254415dbd1afef2581c40877bd39e923f90073478d13e4f21eb0365950b496a8cc7d1d70ccd8469aae3e7beb403ff992a7cd284aad415571454c59cb59bbed35aeaaced2a4b7b3fac4d8452db5d97ebe56056e94e4e8fc9daffd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7886fe0dd28e0c3a4665fc67682a78be6d80c67c31b342541faa6a7f9cd9d67bf922915e8b4de2efc509a3e35353af451dcd8e7c71fb1a03fcd56ebcb0bfb9e96682e7e620b9c4923dfe6c98a9ae11ac6ceacfa93b33859ce682456f58cb76b5c920c21a96172d5a6c9b94c8dfb8aada9bad6868f113016;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h345958a931da934a72ca774d73fe398dfaf83653b19200977796fe5d2e2a4b2ead4f7f77c44ff39ee713c2f78cd9968eaea871800b5167821887fa76a91bf136bcb9cde8431a85f16503855c17e127d1f596ffd63406b04fc562250f232cfd62c3baac96018c4cb1d0ea14dbd767d1f8e5128238c5a3305b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11da814e4e65907c2ec33ea3c2171c6a09fe858c0012927414f470b409b5d8da5643951a9d6236e5c4c7944b694ee5c0bce70ad8e20ed6ec97ef9b024f0e27d8fedfafa6a9dd573d5bda6c62193f5eb220f9eec4066ebea77a8b77009b4ad01ebb6b5afe9f46ec254a48a025472d7f425087a78da2ad98b29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0e8737ca189c3483f183ea9267854dea2de7e95f33a7e0d56e7b4a1d2e02c514262eb0672d053ec5a69b33c7dc0e91aacdeec1dae5c7f4b6298f37fab84d600a6cb4ef9508670e6c95693de8e5b8b8cda3eba8f9568152b3b5c89bb8372a352d745ef49efc0bce3eca97ebcd86c290745c30fb4de53353c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109d36c46071d6969b69dc87d9769394042c58c9432093e3ca3afb7376fa69b42991875c64c15631d4f709722a9b5b79de4c490d9c57ec8f1cd72a8d57da156f4d410417e2fb4ac8f395f0bf44e6c9a3add7fd28133aee3020b6e50c13ba2be9b78b26eb9eb9f564196d66776ec7c86d6b97aa8079a5e6493;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6406ee789b6bf314f105a193f810eb7a8e1c67e68d119ca2dca5b25268b07e268428868d9466009723e777206cbcc939e8014e7b72b570e14e6f5b4b7e1875a720d225a2136afa73b37f3fb7ac4b52da8bdf7ad109427d9476e27da4afaf617ff8a5ea885347b10f9547a36cef38c4ffff354eaeed118707;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af8b638303e1482a5ae0c777daa5b641e645de59f55dbb47f70fc0ee3afb5f4a32d9a87ed10b92b1edeadaaaa97630c9a6eddf1ac11936d1e2eeb1fe1d7dd4d6ba8b7dc212bcf3335501de3228af7015540d0c4efad180592608d00c252dd3f2a39dc8ce33dba5b776f255ae038abb8b75033144790f9775;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bebdd583f3a2b3bf56439ae6e4ab641387182a4248795982c576faa608ba0504458c850ce84bac244266ce2f8eb6c5b5a7659239d73b3b9928c0e9e27765cf42a02d5f4cfd38c36269f14f769bc22fc227ab1903c6c0669f9586f1abff04ab133ef6cd00f670e7fb24fb2fb4f3e55570533bc85880190bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c487f170a4b40624ca54cb3c3f0f0b760f620e3e8c2102a251b2850a06855018e4f43c9b58868fef4595803a6d201245ff093f4eed5eba757b3950fbc5980fd6a9b06ed415856826d7a34a5def3971378ed726a1a7b7aaf12020f97a2cd95c60b425a77d9a1f927388b880025b84136ce1da52fb7c8908e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123eb25763d4062d7467a3afd850d747b0f7f99ab1d4862e5d15942f1e4440d2cbfdf64b622bc84c71e8d091cdd36d90d2e30d044a56848c4111f9bcd77c58c5307d75b00e8518fafd2f517b54a9cafc27fe6864138d576a9d7227bbeef34194b314f27c030b8c9999d7542ea4d48149deb720b342febf971;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb41295cc1f4ef5eb4a7a18952a4bfbdeb472a57d03d1cc6d394b66bae77f113ae8acc062ee5db4ab32aa87367c17d62d4b01d4ec500f808d43c31111d415b28d824197ac67508754d55d2294fc551f98ce6f3bbe73e42f84c2352d0029e3da414e6cb4123cd2054464e0c5e5bc33545f439d28caeb8b15ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h555eb2b8cf1f305d720277eca2de975bfdf3e859543eaa295ebb813e4f97773e28d946c7809e5da478dd71d08a84cf3b0cca5ac53b07780e93fad3e1a07da6cdf537d40a76e4e4990decd5309163a24d683229c30cfb334de98bc66ffb53247f60d4e804e991aceea774d14b61768e4505ab654ecadd5d01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13482ebbb8dbc6c38e9c6aa3f70ab405abba7d8cf48d73147e423d33387bc0f74cdef98f75225dcc67b1895aaa0c0eaa9eafc0f02d97a46b9cc08a13b47de021662af3f97f0211709424c7734766d90cd07b92fb1bc67e00d8f4979e908aa0e9c7ab6441508fc3000cdcf8c739bbf6fa58cd662d8a031baf1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102796abcc5786ad30aaba0ae8dd87b6cac7322c6f1a9eb5bac25efa89044a111cb936d87e8add10dbff7cc55f7c627c4e4198a430e1a4e309088fed5c85f0cb5ce2e0786f03b9f0cb66ec6dc0d9fcf40fca2af81699019e45a71e9473e79961bb730851ed778604dae39e77138956d7bf145b675ac1af0de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h484d83673e7dc7de2bf79f10e890224074f53dc189ec244f90de61aeebc8250e846d94d6d7c68285ce2523239274322981184a2ba795302c1359852552201a7306881a5c89985bb917e03f86f5d56c29940a34b7b8c4eca4545c77caab5fcf6719c090c7d2a988dbc3adae39afec128d7b6b5ec42df62860;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb802283c54aeed3b22c14ea5147d870f6e1823232461eca8f2976819801a0dfa7204d7b7e8460098bd1d125ccc80ec5757c209c420f2c95146efe1b6a4193426048ec14ff042eb607719f0537219aba0400f39a1a8396226bb9904401cb765d504f95f35b230677a383f560eb652208c25be65b872c88fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1641d63e10ae9bf0ec477d7248a6fbea23ed4c322bbda77be86bb10d33c758c4b74f5e8aa405a651d2d271b213c41ff95099c37bb378a3a556b615f1046e493fc9935184b54950131338a53d7062e32a6dbdd159b3b3c92a6eabd83475358a1b2cbe70f6979687ced2d1b5120062abb587c8d448745e8648a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc116f8a69fb9c8fd979c76c5f229131cd63bdfe6ce7386cfd2ac4bda89f79c6a05ab2f0467965fe409a0f4b37b50ed1aa6623779cc7b79025c1b18b06d93299212cdcd911a8cf8682c8dfa8972c8518cd33b38f111158a341955982106657a5de176a20bde9563a2fb18a4acc4ab6dd29d402d3b8eeb86f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175091c8a41433fb12ca9d7b5b0c048560551a7c96e884eff4a41f86eb221ae2ad9ba76749ccf66f09bb00abcbc99705f58b4e06616530e9be1665cd5524b82a1d6c86670702521ce7bd0485c5faa0ac320ec4422154ddbe609e3733e7926311c01beb3c73f996880249f329ca974eee3769400dfcf30bf16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29728da62fb246215529f545101401179661a1dc19498248cdb6f7434cdef06c3be582739ab5eb37498d1b557d91fa258d7034442e3a45d0f85b452f8ca9b79853a9c8baf374d6b98305823b16e818887861640928ad9ed5805c7a6302c3b12562f3bc6153347437130a5e3e8edcb0498b6d109886aa62d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbd525f055cf2777560efae662fc1c04b55a27ebeb5a6503c93d1cc81207d19de8bdc12494cad7346160aa88e72d98d74a31e9c352ee10268fa0d18a5417deabbcac8a9f3bf5b32f4f4e333237a78d5ec8f98b69b418cf519c4b4a323f1d6d33a893d6d90accb1d0017f4d45559b5b7f1f7f777a31aac4b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he544da86a2115ad333fffa7974d41083ce56d0f089b61a100b1f97895c80ed07198e4b1b79b45c7bc4a7b8e2592c946d8c42bc581d20374f5caf1e2bf7fe04adb31790e905d2f381ea24c5d4e98690d7b1d7a6d9de57007d80a9a1cfbb957cae4d38028d6034aa1fbda00d00bd374d4ca6ff5dfd7d736908;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3fbab6e1cf05d73b3b2fce23f1d47c68ecc1ebfab8e543243d5d552a983e6495bc02841cbc2b5fdccdc3d37941239e55833a6f421f9033a26ba772aaf924d0cdcadb1c5001b1a9456662cfc008671c0ef2c22055ee06c02d6c2bcdb9e325e3546fdaceafc915f4c74c79047826e4f7b088c5e0b9d19e2d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc36fed2fdb7714b236c1fca97815f5e668ca41ca5527b4809f15ec92e40af22e58623accd460623fcb78d6f66d354de07836a6bff69504edc956ea3e47c4185f8b69dadb5df5d6b651784051bf673f41449929a0f49f3957481e5d4d47a99df7e9f77d5edcbd253a59f9eeb5248e987eb5cc2a0dbc0cb6fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he51cad983d668ca6014d44ee876c786db17ea4b5001de5db57822fdba89b15a090286e0c66720dd6a16697975dac0f84fb5876d79f8df947ad7060e4a8372e57b6a6cc1f07cea7bfe85bca1c22e8293ca2a8c8a8533b3562d29c6d3132123be9771008107a6d7b206e6202a2af1e9e9672ed3ef10876c77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee68d5aa5c33caffed8aa149989aca7a899b160b90c81fff2ad2fcfd6af60d0b7e2db442843d12cd613b7d2ed48da28259a8ba950a70fb439d5720be5fd3509424f2b90fea2bf26b5e3766bf437218cd90bd0e449b5757c8c053a783699aa381be9a22cdd8fccb73f1bf3fc06147bba32f42a878146688ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d7d35ca1109cb2c39dad278b83bf594002d2db2faaa19425b4d8724832aa86437214aa3eeda52fb26acd0e701f986b7918bccca4c75fd7d6b1bf9cd3cfa8385a068e2acaf4862c74ff3e2865b3c68ca23dea628b559a180af8e1ee04ff5bd31c8e53a068e71334cddd2a190eeadd2e0b871d7e4eb17154;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6200124bd750d5fba6726d5ec6a5ef1b6a44c438994d1cb606e6a2756c446519b1863ea978ee1f114ff9b8c641907f4e5f9253d4303bcbf0afb1d218b7c5713765f58bd892e3c6f34f4b11939ddc8c18419834b63b8505adab15774b0c654849eaa1cd373e6832b40abee4ebc6f8f66db5cc55e464114b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc800f1fd97d46bb0eff667511e2bfa08a066fa6e4a621641dac9c384888e98b6f7b50e2bfde739039c4f1a9ed9528479bfc7283cfd64a1e87934e9535e0160d2770261449fe6ae57d48c13f642576cd968c59f1ee92b5e4063c0012cfba6f1a0c51c10293d01b309a71c4f7232ccfdb00c11a445c4869346;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1691521bddecae75dcff3ccbbefd7b964d470484c668236f1ec53c2aa2cda28d3d8c1afcbfc657a43f63d76c6952a0a6f94c4e1a26158d027855d5906b09e5be97be2ba3db15da95d94f85e11b72f54ae747b9b6c1a2621e88699fb9d2afc119025bfd7f5ae02a2d2bc971deea8adad38f2946d31f014080;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2e2e9377bec3b93e41fc1aea2d671b8f104d26e2e1ddff1adec192803f8682c0f2373723d8a61eab5659a4d731e94cee684a82e9d83c4553e75281258fcb2e0da718c51063e71532030997f366f20c93f81a11de0f0ddce9efe7fe91c83e6fafcf864e92c0c314212e725a4c614a38dde6e1c3b1828e8bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ce1dc4f2a68bbf08d11ae2e329c8fa008e3c9bea3087b1d780a47ee2baf542476c6e89806fae35e6da8af4b053976029a19d88368a28c0071f2277815c9ba6f2e5b0bf75d2b314c52a051f35c398903d1a2f907a2f8f48f12e8cc8beb5136cce89d10135c3ff191b45aac553bcc263cbea7f18e5bfe59a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90ed55b514d96c45595431523c1b76a24cd044449976010bb31b8ecf4419840947edf7c8d941aebe297a1f61b92815dd323f560eb85a840bff4f929280e34ecc6c3f63d8e6e8ed3ff1be592d800a4b6f7203aaf6f9d36900f24dcada90172b5a025b1b78d80ca6bb90632f10021f25e4489966f87749b01e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha65dbfd9cb8f0549cf3c5a8d1cf93a831d1a3b433a82e5a11a3845090127f4a8fddc8d2093e9d5fc593b68b73ae65fbe8be2e12258a54736b88040a6eaeac0ac27d6d91653421a8af0d86e83b8aba599baaed82cc04c148a0fc8383c1b190aec41c1179d1558778b030b27ff6b18c71c8c003b7cc9ac6fb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ee4b0b178e7cf2bbb54943424c8fa69e8b60a6feba03aa0532642759cf201eb15ca6cdb249885ab21ae54a76742c7bf91174c943439212679107a664272798d88a7c63f22126fb456887fe45c64d0c091e67e059e146e6c2a945e20bde6b75d1e913b2dfad0e2fdfe595505c0e3a52bd3b3cecc79a45f25;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16901159dcdd6945b5e4f4ffbb4578887a24b360afc57846199b6aeb0220b86a28d87e7f19f177dab1922f692b4672de633ec7ab5c5de1f1849ad93af81d63c105ab2f5f580ef5fb256b1b98bf9df1b91f82451e3010737bc20d94ec8be598f383235e62c531188ecf186ef0cdea60d95140b772289fa8aca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfa5b897e2f657d1223d916b83dce8b85b1836c476d74e6bf4970f06456c1a58c4a6243d4dd77ff78ab7d7c3f93c5734e9192326a435391010e4e7c9a367be4bf6db9998400c9e3727d4cfae9009256917d2b5b109562dce3a3de3827c7180e745e9e6b3c7987f6f32d3264ace264a7003e96f1c04efa15c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8a1862b8616faa4e87ba90c1c0a42bef578a4227b74ccd3de8d364072abe24e46269abad6d4515320c13cdeaf468dd2a1d63268720af62ce09a2fc5020a8d67194a07ccf58c42df9e7db2acd02ebbe359a7ddc6b8ca2bd0cdcb101e56d0c949cb13aa0b6953f1938f9bd6ea992d77ecc9049bf03a932bbc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h444dedbe4b7748395e6c1532bea9a7b8fe8199b9c649848b462d1d4b21eb1233b930c8498405a2d63ced3a3f087d820474ec5102a5d2e63180e210b4d02bf38ef27707ebc74a15fbb60c014466dad279ceba0e927ad074599732cd3f7bfd94c88031bf7e49dcd3297340a64e31b594c2a7da7a4e4fd950ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb35ec0599296b8332e16718d43f36cd4800ef475e929351eaddd7a9a89f51e4f4460b1f04a21803d9e00383899fdc3afc29f1c7c672966b0e293c6724ac49d57e3dde07de189d32a1018513e0f7b0df4ef3fc3a336b4c2d32b122286957bc056939fd45c060eaa0958b9f80395ef7a9ad1a39b82249b7c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc11f3506e732d9fee7bcff49f71b18b2056ad84a8c38aa6d94f2f1ae51aff3567c168e6c1aa4b5732dfb2d89d5d7f66c86f67bcb03c1ab006768e4d5637041123429c0bde1e1cb920db12cb83f3872c4209cba8d4c109590238b30a97662357a0642cf852b040a5a1ee315b29fcc0e61719341fd17451214;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e1f13e3721924f7d3e851b5f29b794df257b48b30a4886fa526c417027f29b2545139e9442ece222623fad90a247190b471af9673c43b7aa5bd4c256f13d66958f4d2851c1c6189ed2cc3bc3022317e182e66956dd759fbd59391ccfe9257adeed29b81edf3e33706b83d7de5ade6de3c3c75613aee55d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h547e21f239e2c86790d6fa73f1dbee4cced4d71d92865ce900a3de88726389413aa81e67e9fd0901e02893068ec0465b6dd20d7ef56ccd72acdf557907c9afdb62e9e408354367d7ef93a42e3c18a50f411b05587a9466373dd2bd069481c81f79593639b7f500800e8e516ab0e7cf79371b3a4dc65f771;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181f0b4cb6b2ca34fbec5d18d93aa4e800e93bbb926d7f62c5d055170f0378b330ac43520aca8262a6e020f38c1dc024034e2866562d78c138d4e32e802cd6505d865a8086799d53756cc304bf2d5e0664c0aab9e4b6ebb2fe8d42cc61e7101372ea7dc0c5aa86884dccbce08727af784b98fb8d3208d8e50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h941d417d0e5d81d7b53fb8d25c536d7d18382f10f06c1e423d074165ffdfc944154eb30ee2fed68edf8f63223099a04fbb2646733f001041ee364a4d187ec5705096ba05e966a2501cf056940059344ec43b15e4159a34b5d3afdfe5f656d77de6b7f5a7882535865e6f73dd585f524b8ff416ed0342719c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38595338ebf21be092363c2d8433b60d6bce07273defdd722934d5cc15e065a5c04b5cadddf490b09299b1f1968a54e8cd577cf9ddec945004f2bc17cdb9b4ea15ecbc07fb88125585ec75460165791fe8fb461cbb41214b551fd45103674e01e95965d0c0cf7c5a3b1dd1eefc75311cd5f11b7443604cd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18acde33d59c0ae3921c251b585073d62ce3d75a580e7c4af691dd222ce42832177b7546bf38c74879d050acb5bbbc611a2d12dd9ac9477bed010af4b082084136d9b3449bb3ddb913feb7364d0689433e02c1d26a353638f606557f0fe275395c44336ea2c25357d78985808ed58ddb3f6f62b0e320aaf92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b020f15764f27058832b975b3766b6cff4dfd8af09a250466bd15f1fae5ed0e97198380827f892d248bfae3a9beb90a18fc954dc1dfc157833288f1d828b9cef67a2641351ed663a7201685b2fe81ce9b1cfdb3cc82df8fec91a2d7e13f8dea434b14d49ce6bb70130479b46dddc7ab4301d61a4328aad2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha99fb2e9c46df46fd33ff92a5469889b6f1beac378be6244afd1db9e2cb98fc74eee4b4a19a3308ded87fd44c1ec861ad587e704f1d8e02e58d0312406b886b39872979038b12e6d6d7120d6d98f4ca3c78a7adb00374ffe5996e3526f44810fa305c3e66b694c2e7f4fbec3e628108bbbf2450f6ddc55a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3a5a828cb95c730f61ff3441cd69503db4b0e5a8fe1d725bfc30208c2306ec8fc6f53126957aaca608eb4c12eee55c38d942413f9aa52d05c01130673412e6e0a8bfefcc3b392a29965b12556cadd1e58503b8840aceb6e7b5a28b78de8df8692278d1f52e995e349b5662072f5c136babc21cddbbba943;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb48f24bc24e797d0fae1d0acaf6db94a303d60882a9468059beb6f5256366e3ea136960b102b4e71d9eb01f2657f9ca2acda562fec90dfa8e6bd53fd5a86a2bfe61e33db12a189353570d5ac7cc3fd04f7548c5de513b792b1a912712e1ccc32ae71c92d5dadeaf7ee8e2d6a616d7731d61ebd9e5e4c8066;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68dba521d90f50095c77b9d99f7fc2dc39da62144622a5257b359fc8cfd097a12dc0b90ecddae7802a5f65adc7c450bac0cce22163301dd8cad32d41a234b9b1c8d8a796b3c28762fe97fcb2f195421dfed5e2891b90d654058ce4c5dcc91ffa47c08427b61cb4deb3543cae5230385cdd39940e65833d08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ae7c343cdcac2afffb6a5104f5d0b18b20d516b5d3d2677432366cd5924df5fb654a04631a61a757e9cdc73595ebea94fa19731e637cc5493b5ae2f8aa84c0db44da80ea3cb4791d250c8721d0c6abd8632bfc81cc2682d730eabc99a2a225d421b9800ffdad93c1b0bf6a3c10184c00f37de4d02ac20f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heda5354e88b59bb1e0193c324d95da85b41ba60873e289099c5b39ef8083332dda4a36a56005bd7207351c9da0d2cdb09dfac520cd85a1c97e683ca38a1718e7ebef12628421b440bcc24e48fdfad7c2222e518d31d7371bed3a3e6597a84ff3706e39490710b7217151b718c47042cd5af53d97d2a7a799;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4aa9477bc91297991f669e0ae28249af4ef479e7472c824002152faba6d2bdae8cdaef0769b6bc7d4bc923e9cd6ab34dd5cf7d661fb1d175e2751ddb929cfdeb9e2333abeae2dba70f102b159d69323c5675534a58f22d294968610ce4759088858ab85852c1bcfccff425e67fe5f2a8e55510c966b228e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1056cbadad7947bf4024c350621204792a952883c1527fa6870addcc977d17ef918c292f7538307aa0b85a423f3ac3be2d4c9829d49b686239f8dad9ef895c6464055c30d62e0c5f6db0519cf1da76bedd27cf6fc213a3ec96748bf7cd6ab85c0d7779269f40d923b289c2e97b01585a6235b26d7c6b73cb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a3d28964ba027ca5562fb3d40772b8de25c58991edaa138234c1308cc0d162fc25f7588e3b6ff1a31ce1918384a2dea5592144244825d1e0ef0dad93396e1ff9834419f97c885a1d8d2fadf3181c4cf262834763048f761e7c03f5a4da30b3c407a8a3b978e9464cabc6c011099e2b6468106ac90c63a6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b84c395b7268acb1472441ab671cb9ee081a703fcfd6f9ac4cc9ed14d20db945f9087475f55dc8d26736709b95d638f47d5a808f572368b1793fd9c1fbc31f48eb88b7a3513a6297fa60b59076a1bc3747f34c270588fe293e50ba5fdb069c5fd192c91780dad78c71594b236166c7de9ba298e05c240f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb6f7d810729a1f686fc0ef9ceafee293f55751edd78ee31295ead43be9dbc69dec4431b394b33002961151f474574d79b26c444b51b3d1689d1ac28636b84ecb77ec5f60e1c7c6a260b4c256274ac8db690d3f88c9790c51d3f22925e0aed57477626435bf99b913122fe9ce6af913e540e4f16b436664d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f47e61eacf240bfa9db239074eefc94c8b49961479b162501d76d7a8b93046c90dd58cc384f98b6527734b3455d77105b105e2a5407727a52cc7cac8c99d3133f3623782266178aaa86087cdd2680bfa1164018f391cb95ce480402ba1f12a64e897678942f8113244c0ab8eb8d0e0a1020a516299263468;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188737588bfc4fe8e85a3ce8c0616c0d4b54f7cd377e5bda47f037728287c5b091f155fd06981dda96991edbf61e27d8a5844715382af7a2ed06c6a0f13d91dd742776d6a34a3c70ec0666d89dd736c0e53e279e1be25bea8a71f3fc70c147d3fd66c649b53a598cd373dfce949dda8cf3e7e9fa89d0ae322;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ab3f8c93b2c125d2e377181f3f1a417cad4f742e44c22d3a159fbb2e4109d88974622a3f2f59742bc3232ccf478d3362cb3748881e9e6df14298c793d6705d719f02f1c2d4dd2e1c49ae6f1a818d49fd4a188542d51962dd829411a9de14dbbace4a848306cb1001425261f22491d125a2f7e936db8a696;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e5a53c162d215a9710162f8751d3976acb9f87a781b8fb433783ebe8c847970269a46fe8a3d8a9702ca02bb44925e81fa63379c45563825d32d234bd9db84227d6ca23659477fcaf47aa0ad643e2d3b682cafec2dfa4e41bdf4d00cd2ed96948519ded1c3d712280e2915881899fcf8732f80fb7f051de8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a158176c37761ccd9ff58d826fd1a0b2cc09b8025cab560c7a4eba8e5235aa365211d8ff6e057ef895ecead0a23b8c3e97a8ab618027e4db1114de92ba11a1b16b7df650bb6044d9117f7b0dab37f378ca112edbe264064eed7c045f985f3292cc9ccd862c60e6c663395e00b0bd5d77c1f3dce393560;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfdeba4d595b130c01aee849c319bc8aae334eadd6830ddfabc7da1844fe013b2ba3974c977872c322e37188f48e96aa0af24da81604c5faeb288d845daad7c17cf3e7f0f52c3911ae8189385f6b2aa393b082fe4f6ffc86279f7bd31aa0f8a6ef572d1c1e72598028d2baa10dd12e2949377b00d747cda0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d8c7c7d820dbdacf15535282817d180494361f9f16d63c6d9cabdf9d7edd86d3fe5f3552958304ab5aefe6d35057c182e0022714247620f563eddb4dadc497bbd29815768084de0503947372f1f72fb346cce77a588bc6db5c1c8fa67705743d3f603bb5f6e8b891a3e500bd8681dd68aa49ba5ee8a3f98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1306c852f0202af03230ee6bec1a597b9306bfed3239873a86736172e106e984aff68a4fbc4fa46f1425a9f0a66ca29c17d78c1fa247d4aedd4553e278b4addbc2bdf425d27abe6373b19806d41f1caeeb27301f25a6b3402593120dc5e9ef8d295858b139b78d0604878d436d29969ff19276ba4bb1f45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c2d3888c901ae14af98a8699e843931fc8f1052df4fba20d738473574f4eae21789c19dfeb2e12a3701d230263b3ce825554d5df3ee1e166eea93ce9196fb1bed2f8acf3a39b8a010aa44ca44e4fdf95f076e04cd5007fe8223488dc607d6035b65f9e5346e737111ebbab9810985d36a178310c0eee288;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17afbfca6d98edce21861acd8d538f3c48a7d10bcc9b10efe37b1db6ba8218bde6fce604041e300a43fa43fad0ef961569a74212412174afbeef9b57ac636fb59597e59c479ec3fd34ed8d05ab0d42677deb94bb73d0a48c6335c694f6686e1b4f4a36051d3c64258e4f74a00206e5c9843e8b3fcb7a925bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbebfe931c7cd141bccab07f37033e51ed2f9d77226147b7cf102344c887aa38c2d7fbbc76bea4c8b820653923f8ac3f9b8f053ae8427cbe9dbef68ae6b0e367b86dd661078df8c4b3d300165aa79965a4287be15c9255bb55d1e2ff810ac411681f72b826c9a703594f44c12251b3d1d38c2858335c2d65;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a09e4e11ea54d9c77559fcd73efba916adf0b72f992b93d69e3247dab4e015579a7a809cb66f4a1548157a83f885e06d703211b201ee46497da75bee5c5dad726fc945871262fcad2c4ac595d04dbb70e60e7d229c316ed60353e9c45a8b048eb41d03fcc9a6e6e8338049681cbebabd67ff5bfbdaa1cdb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce16d7746851928e3affa1aff8b2e0a03b7f26148ec66315054bc6f65c474859f8de82cf0f2edf5b34cb4e701868f9e7d28b20b4597ca2fa68d4125c5b5e5e55c07aed66968e27d711e9c0c965a9eeb43f8800ab376b0fa1d0d647650ec75435eb98ceb6329946925985b96ebaa6dd1283e22241a69c0b17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab681e8f1326ff42a3d57ff4fad92d4dd718a81779decfd3ba10f604ff7d8a30f885484f980220166241cc77efbb3585222909824b1b912e8c721c4f21b35b8ae6dc0a208c8bddc4780d710bd79c868cd4427642066e189f01c214e489ceebba7ad386adbecf88899f856a2abc3dd9e2a510b27858365274;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122dd42cfbf5afe3f5692ee23676860d00909fa9f61a6e2098956d37a895820e73fa81bf5b4451be5cd120a5382cd1e35707da775e065c04743ee2b2e966d0da3c70789fed506117542806b4c5af54cb205076331c5fc4c3b67866ddfd1573d95133a79b8dee56a14e92438ee22ed85c37509a7289d34e4b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db1b334078d86525d418850c0f41dab45bf99ef813253f8ed2d324d1deee557c20aef5e18b07eab5f87a8ad35a9c9814501d8f6d8ef18ae1a7172da2822bc1ab8acafab33487c1347fed333a55fe0a5238413464eeccdec94c41b06649c179dda90f025242c760d9a0ba12c97e28a8354b8d6ce927909fd8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab43bc150a339ceb549d8f4a56a9686d210a332614f47cdbe4f33c2e4e17f65ca5eb6bc34ba56487e4e6ebba187fcfcf94743c274a535f73301d622fdad31444b24e09cb2677967ca235b4bff4729e0010f99e3990fc0b639bf4d796088f08c382d99a81e8ff0b752cb28c018ee8c279e1775553233fc3ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a55f4bfe8d1650672631805c479bf39b167cf4e4f1249143405e05656ba277358ca169af23cd582c3d4c2a21a89d2237f1f51c28e84c2c05f472b738f4f4580525d0298e5e4ccb031a644c7a4387d2dcd6336e902ebb70359908f47188d6522e8c224c2beb91dae07a4f50aa93e9eb898c1e5259fbac8e79;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4324546cc6f20ad3894f095d046c59be449ae0f4a59648bd91b1c47e093d3f48600c642c31fd309710bb26664df01176d1311cf95f131d20c8a7194d467b4549e1fadca859b2502dc40be2bb31494ecadac57ef70f39830c63a71891a09a42b80e6bb55f290505d00b7b271368cea3e90f756ebc3d07791d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b961e68c4a694bf7bb5aa53639d6f3eaffb67a5464b752ed12736a4c2c9e368a9aacc9755bb1be7d56d260acccb9cda3d11626c1af2e7581ef57815c8b1f4263b5d08f42d907e43feccc688b46d1bb4175f9286ea439fd2fdaba2330590578616a29c344020dd86d2cc93ab2d049b1dc9e0ac6be8598c4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da1ebff955b54ad0c5abcde684b35b25790c5505d7842d9bfdc946c26c6f0975bb8e91f9c1269fcb83274e3774eead4674f3738eb5d6faf9409f05fee730cb18cd3df92a8dd6c7860bf36ea40870106433821710c4a71800c662006a8559e46a804b2ab0d097fbd39c599c9efd8b4b2afef8052bc6fa58d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1414c51a635df57dddc535e8276c4c6621e6bb1390bcb3f5651f90406bacd1e73196abbfcc23d4fb61890ffb1c8f9e4e9169be84b32e52115818c9c42f470e09c5d1f4fa68dcf7a6acebda68cdfe00079582be679bc4f18b771c8089c8ee56efb0110aa8bafb63f2bf21506d74486003d6055d0eb39edf4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104e3c64075bb344bf6de9caf7a8ff11026c92e0a828e91d955ff479e8d23f2bfa864029bc3c00c1f1b021842dbe438b812e8e239c9e8c5726422c4023707750cca1fe2735e5297bb1e0cf26d7205bc17cc1faab3e061af2c2134527f6b30dd3e7e61eaf94728fb72c860387ec2b8b2a5037d9038407e7a56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17396e325f1c2e064dcdd049c5034e3e0295ac97ef8253a537c5edeb234ac02b269685e8a482a953e79055cd02e77baed243aa19abddaa55577ce3e65098176495fbb84c531a2840762c9515c52200c98c546fa9b24300773d17c9c659d7a2347df17ac13904302bf07f6d0ae9fb074080f74b16375d351c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a30414cde9ddf4fccdee94960bf77f4428a29272b84c3fd438534b6dfb8e131ee0ae852ec153a24dd8d6cd320822d9482dee720f5f9f0ee4bfac2701f1d6e14a054e6d3e82c7be9cfc89076cec684bcd390d0f0b5b99d45b2a22c5f9f5cadda697a426b63f28a5ab28e96d0385513df30fd22059ad0f17d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2800f3f72447b9bae8089ca7e9a556447eb9442245d66f14bbc52d4ad870ed452f2fc3af49678f8ab352c0667220efd42069bf9411892793918b9406245fe61eedc924e76cea18e7269ace2f6bb8b51728cee3fabded4ab2b5fdd92f8133daec3cc0c495ed1c4d5875fd509d579be0644c80dd8566ff20ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b5b7f0902da1d7e41ab83e6050af54a19a1260ee82188e504c88ef462f6d14494c0f6dca67e956c48a20f744e2b2dcdb6c66177c465677134d337a29acc502f102f2088419e1a92d66ce0e9c0f67b75db48346384f6d090b68135b8d4c58225139ebd1aed6d1c0f9af82538ccc392f2ebf27ba9156462f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45831770edc7360f05c2d347aade46e9518b4c163d527fdc63ebe72031b0d972c631b25db784e9581efdb1b72a70ba5420b9b59fd349289ecad545f2792c95e214a1205904ed47e70be176705e33dcb856f8e4c0a4c8bf6ac9cef90657f7bc323e572b5f945300013c3f2ce9c097c12b8d338678f97fac01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2eb162e567b98897acc065ed190af108fd9d8316b97944a02a435f83ef4fe9955433734597c8b7a30032e65a7686f0f414c2075750ee88578199acad12056119350ac090ca7fdf54d91ce785cc56c1e8330749d82c59e5fe029350f97fc8abc193b60b7450c50b658927cd6f02e005fa5c8242a58957f5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e8a3aa478baaf21371448c4c3c270c521b2f2e2821a1b5482f479b9846dac01c6204e88355d0404ef25c03a0452080b47ae86bf42b77bb92c00d826633e55d8ea210b2a51f1a1a30b2ffb04a4f186087801b9d107f8b3ca512b0ecde4c5869cd483e785782628cd502b0d0066bd9a2baedc9d12f7c29cdd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5b0c353f0ae5bbd8a8bc5e155ec1e13c31b6bedb6fe258bd73fb3158b198bec1e0ac00e89a19aafd012ca1e7bfdfe186fe5db8283be66dda3a24231803ec8e759c354b23980f0dfc80799dc58fa9991ec4b9b60b629c60245f18ce935ff06fba6ee507f80817369bb61a1dae590dfd628c5d2308508bbef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d177f514a07f9272d787687c289ff2df15da9ab86a07ee807b7ebe14026691446c144c4aa234d59cad74163bb437abdf97329ad948e7df77f1de9bc6c9186a5bd6cc0e308262735d558375074193904ad2dab2e7111105fb1642c4c14100dc47934508f55eeb220b7f914ecf91b01c36ae6549d9aa5e93c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c1a3830c3ba9f52b640f16c7e475ab9b54cb169a512278da5acaf5f1aa2b095984ab6c1bd8a2437859adce4bf75b42ddf5482b5c7f1150de82f1446448621a521f3ca3dab5bb29ed68b3659f8fe59e2f237f9d8ce8cefc65e67ba5ee77760e7e21ea1c2a3d1847fde6c3123c1da9e31529f2539fe567631;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1002ab3f852295fd0bde7c0a703583312724c8690490fb47e1a575fe5798c84aa13e0986f1dc52298b04087dcd5ae91ce13f58ef446b9428b9e895b14713096077ce2702a58ee5aa4e079af11b00040ee55551e3a6882f2c2b23e6024195ddfcd9078c79297b4717f43426609c0cd53dc341f64298220317;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67f9d437c2cc31c239cca10b47347c3de239212f46601dff15b8dffe5d051475f1f99bdf42c0404238c053934a0aaef15501fbc0db0a32508925c2aa2d9b8f87f25a11ba443d92b39a9e7c970cf6d0aebd948221b4575cf2dcc81f5ae7edb676d8243d9765dbdc3e2cba78e308458589bf7643e0128e8e8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5cbfc73e5c7b960b5eed0ae80fadda9c76f366fbc1940a3bba96e6b8bc6c841f4ac8adb4c651abd735c975fb45f3e6d487be4e747b99a69b14c50195bf8c8c59f158e22902937ccb3ef80abb2d7294e893d1e440c168225c348a0e282bfe4377e599b7f5bfd2d1ac5a108c89f1cf9e4368a7f437b681b33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac9cb8f5c32d54e7faff8fe288216280c06bab6ce659e89ac478f4e87528aac35dfcf6ad5545d444c16c1bc334f02a1578c8cb9af16a65531ecef721f00146b542a4369393422b4dea1d58ca060dbcf7f75128c65207ea65a3959a1f920345eada3a4d8d453d8049db82b98da49c53af22d6e12ef4b22344;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b852a764ce401b7bbd5bafc2e1779e0ee0bc899b7ce990eafd819508a86f706091a1f9811d6d13ff427e4c739aa73bfc8cc0bfff48953e61aaf5939acefc8c861226232ea65b1ce8fc1d57331d947681acebdee16b930ee4ae33c2e8af761441963bef135992a61380f7e8a1ed927ee8ff8ff36cf0c5ec2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h93fe4f382c733fa4c96b281dc30a46f269a48425ca857ee15dd707c00edd41d3c8f5c29e86d30165c8f9c8fb0463393889a73f61511318633bcd88556826ef8375685451fbb0ce7e54455cb09332b35a24e4fd9be6bbdcd307f6f78d0713cab3d5f73fb8eb27ce89c27ba0afcda9c4ca56a4a29d119a3958;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1d43c42bf356c97fdc9f29eccc6341c736bc3472d15e4585d725f7a3a830f703835042411c0fed506f68b899424118e109e6e00c2d86a6d8461cc751be50dbbbbb3dc5250029efe110967bc046dd2c0f2428e230a18696215737287209fc8c89e4063002953927a24d46f76ec907d583c9c1cb8e3e424a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb59b909c0f2d54441e32029fc082457700489c4bee4350376a492cf1f651bb01ad397361fb1ecee06bc884217055d4eecd214ae30ed27d9ad45f300acf0f147347244f0332339ae148a1994114071e0d31cf724b06c2d025038b0d5eb7f876561f7bc1a97edac1972d231685bf58903516524d892d01e59;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h560cc4371c0dc6104e3454f1b12a272f59061e17bf83396801d7f109b30b8ff36e617b474fc27d77657a95695ed426ce3d7e241126663a236a87ca4886abea12ecfe9f53a24e3d90fb01f19c7657aa1783c7ce2620a49782c1575f61567a886e6e10b78244e9b08d6ecb6630efa2c1b03d405ea3cf80d069;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d9decf85a797279bf5c5bb6727a7d3bc89d368c8ebb7cede907566ad4ebb1d89a2cdb2c9b40afec01b7d10c00c2c55e02a6b59274e4f35666dd4914f1fcb051ad2c21e047ad61e3f7e20b9f92734068ad9a66353ee802827553fd2429e68c0bc1307c839b51fce6c3a848a711e18a17888dffd4c6028672;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1592ed392417c016fe2229196506ace83f7a7fa4e87df3952e583b30c03ab783d0301be766dea6cd951ed524595680cffd39dabcf3967e867404fb17e3f576387f9d7422b9d8df3717629d69a1842e64feb8b2b248eb5d0c1adac137ee1b1a52ac319cc66c57bb61ba095f53a60ec5ea6d6c4fd9f67ce055e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1baa44b026adfb488a4b7653e80bb382d02ddea3adf5666a07b1a2228a5043172fdcccdfcfea4b0fcecd4e729ea57486eb6c1ad7fda73228679745fcbfed3fe4560af938918e46a73311a97f59ebd95e4fe60fd71c8d4afa9ca154ac4486dd8035689c5f643b1ca68ab747adb86389ac27f5f2c1ee744a73c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e75ce4349e21ce9603b42f3b6eea77234da6f9d2bdda64908202f09148bfa08fbf56318e07cd9f311c0ceee032ae6a6aa741fb595fd6d6227d8af89fd869e3c5cabab143b8ca24dc023ee49e32b7d6159efd245171d3e9adba66b7fd7e6b5da342620caaca4db1acb5c241bb524d8f8632a8cf908a631af5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165fdfe1c50ee2e39438545fafb2f1e5c788e4c5941045e7769d5890c2cfc1d3597cd81d8b6e534d64d4cef6635fec1ad47e303fced41ac5d7a7fe32772d15ffec712fe23f65931ed33c573006967aa5430b9cb2520fdc06ae255d92013641668b24fc9b06b396209b0c09642aba7c88cbeed3a2ef41b2121;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed5a1a724bfaa4b5183915efa57d1e528d1cd145160a0f7a562c1143865007e660039675684dbd31086207dd7dd657591869e92d121e0434329a73e023d8ed479a3eaa5a5bc55c49b06bb5e6b4995407035acd3fd19dfec34ea1c62afdc862bc4d8e8e2bae52cd036dd48c2da6fcb94dc06950787a0af667;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137b8dcff785df211e43fb90c60a3ae3bee075aaa161edc0e9283422affbe3319072c47b51d1a4ebd8c06d54d877f74887b53cff2573dcd979878cbbda21b923f6c23b45374badde12d7f10e9a4d88cad678d54325349102336e16a928df92f9e29bb0916e15908581dc3e70360ca4b784eacd945f341672;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12019b4de80d00ef146bc5151024bf1961d18c3a8621bb6361636690cad12bccd47cb4b00497d7048a39aad6a9a6a180ae152d94022bbbe63f3b045fc6962b7af09718e98520272325df41ee71a7a5971b720445b7e97ae1ae4ddb0023400f917a4446077e3b4594dc2da37031560adb77689edb100434989;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179303403e600c5f548ddc45ac00da236b46c95f16412693ad8a1e28bdebbf33f37b6fc742c28ff7a68ec45c98883236387746c449066ede215353054c4bf866db1c3a19e70cb7f5a914c23ba203fbd24125903287bdc4b8cbe05aac97d3adee2e794e85b3144feb97d8db01de433e7cef3446025cb4b9003;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h159d70f53192c0e9cb87a89e296f961d1051655e451cd6b496797a360d51c9903faea47705ab422eb61cd8e2639589dbe29cdc4d3fa6111a3b64e0779e88492c08e9999fb36af92dd29a7011ca0220881ecd7e568ea96a6be617469652636411d0f00320aca3cb4963fbebf6d9043b5e3f0582b27427f0b66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116ce6829f1f43ee39aa5eaf1f11b1cdace03bf5f7d287762b7fab6c334c5a27bce2e74a6e8e44ceeaef6e9188924a8a0c2b5596cfcf745f1c24732603b53fb9540a30226a819d54be38262c504ffeeb877b33fe7481a6901a4b652fda67fee5dab3b083d5c44058c23501368411410db730252f999caefc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14483d712df724d7b2ac3eb3131622fa38fb5f00e2379271a7cdcefa7ce3e471d85faf56f0a924b8cb29a152aadcd8a27fb6ef9667daa75b368cdfb7a36974608ef0e260df83f1f0a7f97e292d761f9de74238e3f64e5272bb27e4a0876a4565f9fbb6a8f835b4548acc3b404fff934a5e4f13e9af8919f23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fff7d678ad95fd79eb8c82bf2778e77798d20edd6d6243c844b661772f3b1a8443c887750f4b7c95dfb977215528f6d398fe398451386458527fae1a64d68264113900cf30bf679e3e31e78bc9b95223f560e2673107250557eebedea78d20344db8da640ec992199b090c5bad16abcfb304cdf6c2839d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb6ec982215231afe8897190789438618af374b4725346ae7c0b0307e293dc048a30746b54516740820ed508fe080a6ffc01ec919b02c5ffd6baeaedfe89cd7a747ae873a7e89423c733864bdabe141cb7086ec013bef8f07a0450162df8565c1ed966c4dc75e260545e623fbdf9213882285a143064837a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6a1dad4ea2254ac1b4740b8eb6e3a82d31de01643896c70f20a60492fb5db713e228cf4e4c13ea624d24a0c29060393e246212b53c71c472021e885431b2dca5aad332826a3328b9e8fe3f2f17efabc7933ebdca431460fe6af976ad0beded2149d5838642bb8c8161d1d909d04100603e7d5a61e216f33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1212a303f76138e29113af9032445eb8b5ca45e2056e14187d688a88dd178ee303e6358ab9e4df0178a231c4581bf30f570df7c9aed89c2f5003355f4196d914149abb7c05f1d998586e137d6bb08cbcfb27786101a8774825bd0eaaf817fe2e0635664b7aa5e1edc09f705af334fabb41eb168442884c188;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b4e1aec59e301bdfa68aa7760f3b8d2ef35ca3c01488f6c49db3da09ad8fee78b7e078bf7c967688926188d306a84314f6b4cf33688aaf3ef154b3ecb54474da434718c3c1be7a0097790fc41835016392bc553a1cfd0050db8d484632dd09026c1800e9af24186368b299b5549d2b480318fca55f4b5f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137d122079054a3794cd5f1d72af9e1410528ea43c38f495fb75e9c9fbe60e234e29b12f615fd235f39e731cf9e68e55837d1a80e678ad1340bef9574d730210a21db66569775b7da826160d864ef0d13108b7abe93083795b73cdeb9ffcc981b1b7a1652cd2418e191ec9c78fb06d6f11dd0e6b63e97315d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a71b066692803db6657160d855332cde6ea1b2cecbc9260101fb16f8c415a03b60a6833ee52be638effc4eaba709215f12150cb181a9534863e2f8e4a06cd318facc6c1ba0a855213cfca1a8fb0c2bcdf3543fe7de8d0c12f6ac006330634dbf83b57daa6b43b154e212fa58a37b3a9fada711997f619a86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha05971381a247de5ea4802087fb5475539924672b8da8433dd8acaed25d5a153dac134463e19c361b50d519b5006b0de89ddb94360be507984a85898f5350c9713169cd6eedd4f14abae935abb89e3f730f48dee6f4d9e8aadae0ac3ada27bad383fade594940bf41e70821fea032e5269b3e4e5de4423d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f2555c7fd839ab0781349d8ffda3a45b0447a1797796de97c1769394f7cf396c5e4e63e96bd8107fca7473c4668eaa9b2a0a01a2a04893928204733d5542814a32dbdeb3046c84e94af505d14d03d076e1deba1d1dd4c22239e773e4362352034aa82ece8fd817280f9e93be4ae6c564306df6a4cfe4615;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95561ce0233549187e32c25b1dbbd8f67918932e2970612a5cf1fa4513556bc9d8d5e8f2d1bfb29550823721fc8443e429381a97bf482602c299ecfdb04203b2ccfe677d07ff7aedd7a27b8927d183c471986fae3f8ff0f2fb6cf826503c1120e818896010557fe4efcc77d3d4c863eac9308e8ea367791a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eece2db5366420cfbc9efcb1616d1fb95b3242f54f27c8046e04bac5c110e85a06381b1e30918a722027dbbc1eed37a9587fd027ec6aa5f9055a3053e62e4ed65a127b90f903a9c2b60c1dbaab9a13cef2f20c7511537cad3687274a545abeebb262364d2e2caca203962062f1a8f347b8d9be9085c4b85b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf812a0434386b9a76455730e4bc73f64a2f362b726465f5ef3071d94e5461873478369145e743d168a7f2e137b16ed1cb680918c966c447b3efd451bdb8db699675824d13b787ca13806cd3745e1a132837e6be911123905245fc39552f5db8c779fb3ecccc6dac97def0ec98ae29a4daa64fe835a6c910;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha83ec72f4d83aacc1e053c1ea4cb0658758e36ffe0358d467780f6950556019861a8e61e4eb9fd77f3a8cbbd8ccb9867f4c339273e1731452aa473652267206608d1276b01086311479bb09f813446d160588f4d8186d162a8147a26a91b4a3e13c4cb2a15290410ed2126fe97b1ce5bc8c08de6aef00abc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cd06b93555053062e5a47298a430160ea07fd36c9b139d1d952050cc75bb6eeaa465edcc4a2cdc36aa0d5d72be5a403731d43593a7244b4607e5cf35bcc2f3c147569ed96da8e767995d6de753470dd84f9afe5e3a248a5271b7cd8fbe94d02f7ed94495f7f9820568ca24fc01737c4f2a0420fd6ec9a3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1884e5ce92c70d18eb6221721df28d0dec5fe47d43c5c0c7e03bce19f47025f66678be3e5a59d49fa3e0f4746bdf2b544ab79135330365f3e09c5ab3789cc96a16cc3832a03d775267f8bbaa4dbaed56001a4638a82281624225b3e4ee323cb27443e9caaa089831d76f55c138c749b8f4ac58b1750e69714;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h291a347f81d8faf2a45fb30a33533d4e367d4658bda8282cfddbb62b4f1509966a2f3485c9953af49e2073efb6fdb2b8fc6dae25099d317b8f2991e95204abc0a12360247f0d39dc381e06ea0a9b324dc1d102459772516fff8cc743b2432ffadf74c35ae8b96c0a14887d3f5cfedb5555b63d5288e48e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10908e31e9845c3c0e872874292160427d64b9328e88114aa226704668d6cb56e0347c0961c2fac6b1d1745040647692b53b9a03599db2198ca9c9a39dd7439736545031cf2d23ce2cd170b49433eebbfaf2386ed50d090297284831736e1c43675297190d4639074146ee1421d4e4d74be70db0a0e80aaff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h756034f1f8884e32dea8df251ffb61f5f6ae416e863a73aaff3148e8551816e801ae998274666ec01b565a9548cb6c94db17e7760c6811af4344719ec9e3ab1d89f777f557a0200e7b29d0bd09f6977baeab416bf899efae3eb69d0c136a0e9fed9933d510fb439d966ea6e9b539297368e8bfd3d225c542;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1367c35a611e2f9f0cd849d5180e1e68d7e5772254b0fc6a17ab209e9c5673afc9016c849339f4574d4a31a838e5903a51b660213591097aace77a0098812a1b3ef74dacebb443176be5b92890b6f4870801093ea9a4f64d328051f3db7a9f7be79a76dc1e5b6a64feacb89999cff9d0e145424a2eb284428;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132131db1247d77783473e442ae3f9454688e8560a5a39a5b131c5290f7f742dfc3c9eb10b0c44839fcc1b32351f0f5f774f2f829a112e3bf319f3f1ac5e9fbb6cb1d76f0fdf23c129c22c18e83e38fd9823df219bb1be0bc6bea9a90a10eac67c407fba0074578b6a6a488d6639f61e270788a6a80fbce35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ab7a11b96c1e9b2257ab79ae25e085bb649082d17d1993936584b5fa4fa050abb4faf433896e7c82acc5537a52e09eb2b0acbb8985e16d022e7b9b0ebcf8bc6687a43fcb575e6b6ee602eb5598b7901e96683b4cf39ec3ba2273375000b9ab6f5d0bc1e92246e56d7fe1145e1a47cd8e7de314ba1ea218c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1865ac5f2b4ecb1004976e3a793fc80eedb4d03c8c80cc26af507fd6713b9a750c2f726bba0320d323ba4119637fea04b5619cfd12e14c0899234acfc63b16f82cee962451bc55b0058bc7e234be14eb303de1f24c504f95b85e5b97c4261044e0dbc8e9ca8eb8ce1607495eb699a646de61e806d3f88c04e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc399707a26f0e470c0091438c649b6fc72bd59a9947977f78032df839dc8172c61dabb7ba6ce7ce942fbedbb84a5fddf87d64b6fc243418418f469542c205984ba9da9f8740bdbd0517a07d9849b93d23e52981f295041f5edab80732c6d167ee2ff7e46c7f93652ad02331158321af8eefc7d5d4edba94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e40fdc303c9d7bc049b3b0ad31f6ba38d23238bb6ae766581d9f8cfe8c3b590c57c8f428d95afb573b7bddbba9b347c7ba4770a87fbc898cd686e2521ecefec47ffdd8881b554be6da104f148b054199030d1d64fd44c8d914bddff77b4c316c1f4705519a50e4fab96459a312448efbf27d3b793362166;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16857b5e27bd8ca07e2279d48659172c406fe4fb8e907050d87b4ea0466e48c72409dea97ffaef5da1207538df5752f44987c0a07bed49d28ab2e3ebb3670576f0628316b51566f041fce90a8bbd8fd89aaeff2a6a99e74c1f56814aa8d1177c4a44a5b250cbf2419eea0ee6a4a98160b3b15c4969ff7335a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7535502c725dd04727aca527f1a6052e7f2407a591bb60724488ab5ea73ce917e55957adc8188dbdb72fb8bf448a912bda062ff3bb97bac48b5103cf1f48bad1249703f1e8776a9d46b0d59694a4c24dfb504142a47e38195a6989450787c6af1f7fa768df4cc671757f8304703cfbcb0034dda87103b403;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe5bc48c75cedfde4e38ac6f4e83d8e6c6dd5106d1e61f1038bade85ee1ca21284f640a671b8f80d550fa15639a6c7ef3dc719fe6a47a9af5d01e7a97c65a11b13451eec8bc0732b2a3490c47737db7c0a7b42716e96b82ae3d0de7988799297a37d8b5da990433bef312c341faa681938c3fdce163ac735;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2806845bb322fcd908001a5b2cb2f59f512afdd9db68536d27cca8fb6666ad68a52fe0f34f535d9ae54a58d84ec54678e0e058d45f32bc564784551d291c56b9af8cc3cdedb2c148b530bb22f3851f9b5e3c489b4eefa72d73c7dd94c9901874becdbb860e5d200d9eb43da271b1790494a441e2e51de91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85ae40ed73ede83efa426b7c0c3e9d2acb442872d856b02598d3a3db7e7d04a59791f3a3c64f3f6abfaf67e6591fcdc272d25bad2f9e97eaaec262e75193b071e9afdeac293a67d21bef2b36496ea990956c69b6164b3d1afdf2506d0d88f01927e4fb1d768d6d7ae86c49035401bcceb84d45699b177a38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f4b6f3ee47b46ca763cb338e34b374c98d261759302482034b55f00c1eb24d3e6eab014ee3412441a4c8372986f46d2639089ac54a9bb4b024460c40cdbbadbdec95d1848164a133f61b533fe16b59d4a532d3521a59dc7d71b7578c80dcde8f17f9820537c380ded4dca93240ac3e12826191c54665212;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14524ad39d487c2ba3f70e5488e22e11f7f9da4cd3cb42b0e10b1375167ba5f067ea55d4e3229b2e5b9af965b8852571f73994a037ce4f2106bde2550d9990deb4cf85759f6d5dd9bee574072c3e2c2119ec9eac707f00651c334368d39ff5c264efac0d72149a836414c8bc8de0a297189dc353bd284247b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d47d0a92081468c38d6e54867e1db3687cbbc9ef5d2770cfae19cd14f68a95c7e995fd5b0afbeebade7ac0cdd89b5eface3f33f30aef69b2f466aeb2b7855b7dd7383ad1838bb283b6746e321fd643a4b4e932d2633cca930f03ef0beb34dd6dd9cb5ed315bed0b649785ea190698d0f022a948cfc59465;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e5be3f0ae5bf7abe10ca7c831616df1b625762d376ef37b733402639095e2d10c5d63cefeb6e72fcbc5d165860e59a9a97ed838b9c8933f4795c6eb8e846344683feaeb8ab7d2827ac84d0e22d394a5545bab3882c478a92a55048c980c8c39d0c13d5025bc14ac62d45243f7c9119900e5d756f92b06bc7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1177e9ccec345db0f62c446f2af742294ec2f9db6e2ff471a23a2155ca370d4898586ddf45347678c51cc14d45e9b848347a875b2c029de5f3a82b3cd058d25cb90c4de4eb6e172a6cbfe78d7a498c0120cd575fd012eb3a389f49583602979605728fcf46a2c711435a35feda8d055230b967b322f109856;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efd91a7a780296eba3505abb122f69e917aa269e30742ec0a05fca49b2ca2aa04be733d5c7c2608bf753c3fe2654eb392cf4041f57355c431bc90629a791c99985a17193bbae4ab9bcf0f7115b2330c513a4f1a1a90a60f8ed8c516e9004f5ef28af428ab1b0b659d008ce7ce10a9bbe60d42365db2acb69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d5272188c05bb45e52e67c22a143cc7aa2470d8622e29a63e4b6f03de6e87f5ebcb14e149009a79df7cc3bb7c0c48cd5da5a52aa8f17bde3e85a70f238e31edd381c013fec18999289f7e12a2b8479f8f097ddea285aee56c0cf13d4180c0a11b76cb805345363a331f654920a7aa9d33e457bc2a66a803;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132d282a5cffb7ffeea0e12ecbedc5a242c0d06ab813c4a18a091d0237eaf495fe114aad9b2bc82624656bfc7841fae8066d177403921742e32c7c6d8c6e37b80c230426b8e9d33344136593e1ee1866ee0a4bfb73df71ae56da6d6a086c155fae7a5f180504cd5aa7274defc24bb57db1c5edc5601c6200d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd2ea97e0e232021a93d63baa0aeba66a46bafd30eb4a48cb6f661c00e7be71e521aec1bfbfb632517c9f0c5860435f5526c0a4b884ff688c9043055938385b908df18946817a95b7fa2d6310abc4a47bea2f166ec8a7c774e7ddac7a7b3da285a86fc8e564e32415b44762add5fbfd580b2bc1ffd19ace7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175c81fbc2d375cfb4452d28c9acacea0cd65be58638b46b3996540820833fc2d8429b85c473dc8434fbaae70fc92cbd586ff312722c049a83d92618a509e95df9accf59d0a73e14c14eeee41b5c6885f37ac46ac1f66039b4c38f63ca6c458b40a74be19086a635e5e8213261c5d1e3fbac8335f696e003a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107926cd6487c2cbeec480b11ef3addea4517e8616e84eb3a4ce2dd5625ff2dd5381c82990a6633623d069680ed785101db5468669e7f904fd24a02b76ff1f60153245bf2e03e6645bb785db5161b489a617a7a7eefb5ef400d5cf204efa8dc5833c230ff779483558b0b76259ab8809db33ed807a3456f30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115a3fc4434ffe5983b5d25ef7c335b948c7bbfb8a574d44283b8d0198c5de9a3e32be86185230ab4654a4856719e4017231ca397a1c1ccd215c03fea1cf95ac4236aec2695f32ed2b74986542a98e18344f00d7ab815b9d3ab54d1f460974f8aeca97ff688d9ff98577be74ff739b52695d057f3dba122de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dde56c42c06c472d31a9ba642ed52b2417a0b743e205fd18939bb3aa5b629b6d2cd060265023f56977519a363421fdca9058ed77b1a0ae77a58c309b08988c15f320c5e38bb815d26c54356123d357d56adb6974bc908a86b7ef5d1015b995f8de26d654b5a3280dcd9ab98d7169a6e1d179549e67d9217;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113534496a280c9f28ea948050f8771d3c92fcf2b9d771a406a253e90e96cb9c54b2554831c1cd524c97500b17de8751fe9612601a44f66db17067b089d4dd5b75986be163b52c694abae1292951eebf7c154ab39bb364a3d9c179662eff5b970b5726176734ede41cc9a04c3f2109aecc883411dd2887b76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4de18ddc290b32eca6db7f04f7496cb9ea22c9fd0612f9fe44c827bedcaffe5149894f2d8c3256b80698e0a259e85a29b40518498b799c67426a023b95c4665c39ba111b60601335c886f79ecfaf547215d00139762a269a6c3b48ac9a9cc5e7fd882c116157bdd1d96a88b12ffcf9e95d084222e7f0957;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1717decf6d904b42f2cd856f4c7a7b6917fc8bb4b2c3af8b7ee4c1381c6e3e6ccc42aef171c58ca1f35cbd35e81ef905bcf35a7f11505c758178eab30a8b4da97049f1f6567731a50d940b06abd0e1d0a9506a04f1e868337b6bb2632c913416f43ad0d3f363567a6e477f2afa3335d0d4fcb827200c4e7c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c485a0a029ea13c13c0dea9da7654bab875ba50cabd49b98af90bb046c52b82e4d65555f0cb7bfd7caa588041ca692904e0ca550193d800b60863733d95a0571c43307d92176812d19597a9d133f0583c9f5e0c0ec7b2879a046eede8b299cdcece0bc3f637e6365e8d5908167a71f060fcb34c70f518659;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58092a5696030fb8fc65f5640da336222398cc384e0208c2e8bba3213df907bdb4256f0a93496f775f5018fa787abf89c0f0d4195f38c470c94ae95fd1004a4acfc64ecf348ee28258c40e83864ef74b531afe8273ac2401f7e192d1d1f62eebfb628566011e52c546f0a2bd317df0dc5e27ab9d33f614d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd1fb0bf6c1c1034384937b647d02eabe7ae3989c5e402c15e07da6a95753023223e92d60d97ba408d40a4a169600f12a8546e43afaf66cca46a56023b5b5a5ad305ced6972fc7b744d1be72016817d609a1c6a65912bdac50143fcbbf8f2079c8405ed50ba71c362f331756ff16b2599d45f8f045f5d0f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7e90123a7494d43a96cfd2ac004a583a96b40f13d5d5ffa07df6f6703d22dc380e10545af3178e3cda7e423d006f7ef61cde459f16590df729177fbf524377219f9d3ebacdeb1d5e75ffacb1d98810ae2cb6d1eb4f98d49f6278a06a624d71c103a64bf0a5088c68228a7210f03df094ac3f9ef94486a1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aec03ebc2a252b94f996459579c77cff843c009a35cf9e2b3512e4c43cb7fe912d32fa5f022ad4252096d3c3b3c8143852c156de8c0e4b7abf23b428a4804b33cbb15abae6f13bcef97747fcfa9d2cf339a9f46fb47ab83309b081a9b311833154a3c855e20408ede9f4b9d5d80d011b342a3c6740ba604;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3ba47ed62c5aefc59c06cd5f9663277ca3b4e1df5b16191879cc58884f2b5eb114f95532099d44e396ab090b901aedc665963af0f96f55f174b9429dde5b8b76c0bccc4b6a1068e7b940cc6cac465e901c94b80127e69a20c43e7f3892c5ed45d9ea3f9990d4fad98edbc2c6583e739998254f6b4ff1aeb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a26cd578c9c747e053422c0b472d225bba6deb5676022ac30a4569f2cdb918fb48bd68cf3ebc3bbae50252662aa6931397fba58ee7537d135f1a91eff15363feea3e10d2b9ac4fae2a8636162037c5ee10850f31e9b2b7f1b15559a010220b33f3205a648f0b33cedc44c4c5efc5adb12a9f4610d1707824;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1231ef3404dad05006efa3be949816e854c2dfefc0df9b70e9df1dc46c4955d3559a5bdc49604e1f93a773f434669077c161c0d990157c1c3df303ed440031cb2f04c5460b3c0fe6c82ff143714765aa41664c9260f737d2ff93d7162d2e78423826116c76db6bad6c8e284bbafcf6f501ae818f3062f18;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e14180b2b76cf541edab4aa5cb2a565df74b28bc330ff53d447f45c6a54b20c8523a4a47b8c6b39004bbcf9990d607184470f43d74320066e35146a941cf05ada189da160f87af96228f3b1eeb33a7f66975e84200dda54c95580a6dd39726f7942b624f4690b0581e791c13e7132378f3e2c0b1477d39f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9cf70f6356c4cc0c26f03ebe38ed149dafef910f8a3fadd0ff698511dda8216f5eda55c62dd261c8aeed0b47db7e3bb3ea0b7017a72462ba3e9e3509fa06ee71380de50b5d2d8fc459ee24360dc62fc632f4b290005436d77d4555897a77d156af48c1c26728210b75193e48aca0eaa73110ff45d7a3817;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6be8b8a594ab2220f74d3cee93e5e286fcd723901bd9a16bd2b3dbaca916ee0dc5c143258412b3181b2532b098c90de89d0513a7f9c29f4c4ee276f7ea2adfa4099bab03296b73daa9559bc412a2035c1da5589265bac1dbf67d4f4da4f1f429a32e03a970549c3ca8a8ac072976b7504424e0ee62eb447a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h211996ff674363b269b4a9918979d90261c7cc69ed14255e8eec663b397a192ff3570e00e24174069ee8a72fbb6a1878079604edba2981a664db85b378f9de86f1e9beab20088a327997a53dfde1abe5d54b7ce305cfaba37393e54dc5eb5a59c3fe8a6d7fe49f081c34b336004b3ab52fed4b8f3d922a22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1956ae2b2b0fa773490f51ba92164887a2ef380ba5fff9cf18d5d4969b4d5c7e76ada5c8f207214dbc3a4f8dd646c77b574782dba1f33482be71432566c5acdf4cee7f90556b5b838b0fa7491426b1699a2bcb94b52f0b0e31caa27cd7177989f6cd935008ae0fac2a7de4aa8fa4058ab952b091fbb9193ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had5f790917ed86254508c02ebff8049885a122bac3a67095c6a939ccf73d65e0c7114f5f1d51b056c9f3b7468b7c66a93b90bddcc4857e21d6cb20ea2081d9f3b0f01e369312b4246ae83b683b8bac97736eeabb3e9b6e5f1a1e2fdb81d9b0f969e73204febf830b6a7ec44b1a3f5343da53746df6ec511a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de8d0eb4e53cbf5b46c855cc8607ff672ce74e6d6316a7a955c5bc5fd5fd632ab13aa2052f6e2a07703a15050d7d69dc90aac7d185a68db5717dc1c831c5a98867c3130d6063534debaf71b02f9577b40c0f3edbb86ca0c9d193d1a13a9285ec123652bb53dfe913020c404c4bf76928ba35888b3093d116;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11602def24714ab011687fd56053759a73c409d7213795ad6134e23905e846c9f08bb19c7c8c89345840fdd46fa9c27283c75fd9a134db712c975b5abc270bd530d4ed1e10b92bc1cb3b551380e8c2f8e0405d6ac7c7a9a4fc2c6a17b6c97278da1951f6318eca9fa8eb0618c50859250829fe0929a3f4a41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aeb76704c53ead60a6bfe8a61d262b0d739491112718a75003f8c5ae35de174726e383d4e553f49dbb5129cc90cb2e2133ee5bba43d3f45e6891813b5004ec912f205434551d82801e5340d9bc700663f9ea58e448764fd8a6592e1de84851ae888ad15c9182e0d6130f3f7d716a2bb867c337287f1aa473;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h777555614f850332a0c44a08290e76f2f659608400611af244eda07b2a18bedbc6f220655e9a77eea8af92b6d6525220101a011e9c20cc86b10dc10b4be5dd06e29019dde586f177ed12a53efe8febd94246ab563c6d52fd2e942ae6d49e3f24bd7e9aed728e2597eed44ccc589284458c06f90395e91876;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26a69f54440f491fc60226127de6c5a7aefc263bcd07c5b029115c921eec6dc1bbb01495f420761f69297872ce9d436b135305c68c3a310391f105d1a86a2e41ffa17adba43ee17b085bd25d64c90e2e576d8919878e306014bff3e7b6ed9f1297493f7648d4f9404ebd179c11ae4781d272039dafa86759;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175f67f2709aaad1a908a6f50113202fd2764591735e2b2e02ee282816f2f2ff1ddae4734f206f9f427349a501b458ee4efdd336d980c8e402ddf1936fdf8224237dd6fa62b921ff9d4527cd252a9c5eee659a4b00fc9d3fb30ef4b565c4383fb05050e08508f13f5b6ff7fed91146ba544750755964d9939;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191e66f5216f82f8dcaa058d7d75b9986044c1fdb816db60f217f19ebbe9fe3346e27b6364a9c2e44952d711c26005fa0da458d3351e7b309670c4f844082b0ff76e01f3535fa8ce51f32c5a82d0d2411d807addac59cbe72411b716cdd0d3d58253feb35f0c9c7513e31489873798cb48e6436f475d3d1e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19aeda41f21797c9d74fa7563c46e0b7c02ffc89216e5d28381ea4719ef35de1303f67718868c23cc0d43fbe58b7d06c1076a3b0526439bb5c416d6dcb8d0043a79f5d30106c07b36a09b9bebb98b4156c96ee07f6f305f0dec51c6dfdbfd4c2ac07ede04f317be88a4cae1faad6e43490952b2bb1372a85f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6da3665a9bf26b169a928aa5b0a2e8603010e77e799ff32a4814dc06b66c09d0350bd03361efe11c4e9d540059d3e8ff143d53b6ab9b978143ebbdb17f36e0f90089be64e693eba01537ce51404d007f0111bee01eab23ba9ac8f2f193c52b2e9adc6932f6a1b8cc2ad8bb9ff73b5abe1edd8fd44c63982;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf80d5ee6c174f4e96ec1832d5da92f57371ba849ed2d95390fee11437d2b497d4519edd76fb03327d6b6bc46c3a487747d8cd54cc35b0fee30b563e1c5ef8475d1c1fa85c3e9aaeda6b5e56643c612e6a18009ba618510586b620c74acc0a08aa860876b5f3fcaf981eedb6fcbaf6e10928efda71dbd52fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167b4157c9bb424dc24efe7aaf471ad90ade5bea56604917f75f5efe3b6332356e43eeb50807463388c4b832c810170484febb995fda96d2cf51e6df31677615e1abac3d31092e16e11241545705e4ba92655603227fda3b570728eb7dc39bff07eca36353b2c704e8dfc231a4a6746b47b37a704fd50d418;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3f1a221b9abdc4a92d80d254f8d35ddb252ce5bb9dbc8b7c3a4197d25e8b1d46243a371c87198f19fed5039965673d667fe06065b700e89525f8e9792ebcc772458f3571538a3433dc07dc6d0c21d5093e1ed78cecede0724d30befe644e3cfe365e217899a7df0033260e5a5b38b1ab53bb81954667766;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce83b5538e7f8de5f17418f75e0bd52fcfe6caa8436a7d726bf01ebaa076be8441b7e0b50bc97561abf46fc6eaf28be521995d543622035a22ab1f5eb66a7086948367960be8d912544a0452e94bb537930c5ff42942fa67869a0e5a839d7ac7f9aa59de05ac41b15d72f2149a1c9d6d8530296ccc0746b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107474eb6a4d43da8276e803be57e3010fa7045788276b47790f7495c58be0edcbcf964770eea5c24e182868999f1b3e726fa3c8541f448720af21cd3e4d5992cc8a44da66fad40dea8b18507966b220789e21c27866934120ed9cb787c45fe645e22cb98c38f577fa948655714b17ce7b9bb835d8f5145d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7891884303ce092be911ba2f571b429cd1e840bf28d5969444d3d32aadd6fbbb5d7cc275b9220b90245fd3d87eb8a4036421982cb5c1cb3be96c9748d9a749e652bc0bfbffa704f811c7335e83f45c3b336078f0dd3f379045d9c26388c16d0f78ef3cd1a3c5a765cf94291180185f4d0e222f4b962ce5fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1716ce762832a77db118addac34ee7b2b9ba1f435e0cf1f88b8854cec5bdbff33f9d7d822df7b93fc175d9a8051a61c3d613dc56e1b8df8ba14d3a2a56dc8ffe47c0e226251cb52b13aba8dbe70f1d0a83958e9171d8247539ffe7adc5ef06aec6922f7b0d7b0bb25b7a90af269efb417df4731c783353ac0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132d92f9c8ad527e5fd87fb4f18905ee6bac73f5e0fd43ca712029bca37f02c0c0019cfb50fb8207a96f5674fdb751d66b25f5aaea00ad277c4c42cd1eb42bf694361d12554e799459fd51e7f404a549e2b67a4964eec6b0d59d8a76b25a5b9058079ab1697ab9d23519b692190301b63401a6932ddf72fc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da7bc3068374d25138d825ea21f84380ad6ef72c52783ae29869b1219120a3fb4c079b10ca1205f04fc0d56d3807c2375b1a8ca4992b3669c20fa3cc054aeb6283a0cf0c79c71f51ebd6992b329b2960afec7c98f44b3d8d1eab0426e31b6799683a5edef4baf9c128faab99a2e4dd32f6a73a54121fdf51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h890fc6586f3b20214155b6faef65bb467374245a044433220b998318285977c09d3e8f71a29e14ec5980cf4497b8778e58526a04fe0f3e4f769dad9e0cfb229df3675d20e36642bf8a091abe4b3f67e6ac9d5f3564623ae26a88fffdc861884e1c2b4a0c11861b2d09a9ca3dce97993cc55e539fe6397e91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd860bf4fee8e3515da92297d2c0f0302dd9cbd4a5d086f81dbebc2184ebb983a77d40d67834eb488f65f1d7933de5331602aa7d41f606e29a45539bced51bbd70571a4cb6562b7bc1c093e39bf561b9999de97eaeb175bfc9dc80c086a0c5d587a245d86995ede78c34aaf7e71c7b7e561f6ff667e0bf285;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195118a2567f867b5a4c8fd2b3d463ef7d0ff02ee1a5d972c9fd1499265033401a2a42a0564f6969547a335f68c370c524a4e39c9c045eac720486c1ebad4c1c51899ec6d303ff7726ea672721e8d00e1892e8e98301c196b932e3fecc20bb66044974621570c570a5510e9fef676c4f07e7d109dc1011be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ded0071622e8baaec84c8009dad67a35990ece6ae2d89b4da597f46b2bd6378f003c686c79cfb4f5e7a5fdbfd04694dca3d1d06f9050b77f5f6c2fc24a3ff3686ff3b882e393e6d0e1689705741d0ee8538e7681aa2ac262839c7e169816f0734630dbee051f3dfbdafe836faaa274a43e2cdcc12f0bb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a4022721e1e98a2784458642866d9ae916c5d3c78dbe30677cfc2e328c9a2aecd0d6f31b809a3eda7c87aa5273b2d93e21781283c35af844642d80f670880279a0b7c63336f31b88f670052ed0599c5120f34a33cbb6c85fbb53ffd2e49d6904166051d3fa5d9ba1dafcc192bd7ca05fd0874115025e9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f048f54300caf9b913478deffc3c0d437d094029ae98e63273e6f3065ebfa7d012bb42cb5fd4c54afc5e2a368d9d9a3c071ad1c6af30f978f03605386bd43b70af0cd4ffac96edc32c5732e04743e2e8fbd717987a7b25f926c001c496b22b94805aa5e56c8091730f3aedb0b491d15d17d4daa1ed491e26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c71c4e9e792ed2aff807fbd5b29bc1136c56382a419c4c30b3478620ed890a495c0b02bb5a775bef57d5eaf6837c5c419f37db271c0ddb4b6d8364a7fc71cf99b87141a2e8324f7cb3097508b5c7da423c42f30057b75175d04e425e373d0703ce6b994b13e2606c0f701a0bbad127568ad9c23fcb94c54e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haca63b2d93a421a174d1f3d8009bf186eff3a16394f2349c24f9124340b707b94917ea5f24c3b2e136e2bfaef16e35a76c1d8beb6bccae1dd2807356b5ddbcf6329aee775c7f2d039cf461f2f78266ee2267b215ef8c758e1c5c55f60ef8b011f92046f20e7257db58807d5591114425cac9db22cc043cdd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d4fac65dbcaaba1f97e69abbfabd50947708442dc0a7dc6e051910622419331a3af903f1f862be92010f28f536f43924595de346f9a208384b56a604ed4026032486710a6cee2475c4d950a4565a1c14de06bdb03859ef1378562e6459c162dab57cb5e9c90e325eb0fa4996abbd0ae90ae376f5fd1c3e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3ce9a1b38553d80433b0c6835e39ea515a92ed62dd638031365e9c35f37742991bb1c75704ed5435e2048c58a97ff33e647a05726849b24dd12c80b82980703ffe3eca783b60f5b3e04c903a52118af52434f1fa45feabac98f4985259757d71968fa20bbf02255e8195bd4df84597fd419a2c38075c3dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62e6279995a9aa249726bf1bd28c27106a5c5278516865937516b92e561d9cdcea9742b82f72d02a52bddbbb98ed0578954f0eaaec2b86578cd44656d94446798da37e37adaf187b4f9eaab1ce7709ce758cb4044532ad34caaa85f97a2c170527260b302fa8f66be65cfdab0896cda4f73a00b998fa3066;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h177b34db40d5dae5032dc82ea60b3632660e717452e09a17ee22bc526c1f22a5d2bb3d39c29b7a05237648b222435065c3e90c0571c5b85a5d98d09d5cbefe20b665e49d73ddb4357f62f72f622a322c40421b0705fd9bc4f69e5883735cf5d2b0aa43bfd7a3562ab6ecce1185f5b3510920eaddb52a4b4f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3d4afb8210c3cdb465fcb1e22a52a5bebfbc86b79d83bf55cce92183d07165f6fb67ad5d5625e5002031f2b3853ba64b250738c5c4a404bfce871e635967f06c9d222eb5b48a375abff7631e6f15ea04312f49cbaa8a43e437344280dfd0e4801b30c4ee43302b6c3c8d0b35ae58c94f77847f40f4163ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1793020b69cad68cb820e36e6c2678216d67d68c6df214e4ea594f045030d3c657fb5a0c7e5f2e92147f8c3c9b6def9421a08532a2044ac0a1cf1a814a4413ba809f36b44c8276a01011daef8da180730447cec63a964ff90caf2ac2314b19d9d8590d688ac81e8e518ddf7451eca356455a9ebedefcd5ace;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a4a9b10e54ce4bc6f335dbe383dcda54e9d7acbbb568fddb8ccc21a16ba652e44d9de0e56062d54a2e1c9a5f3940d48d75dca9b48c84f6377cde7696083594950af8c5eee23f7b047b75b83891cb0a22a7ad57751515e7258ebbb4c2de6504472ac683e6a1e598a3648ffa5ef37dc10bc3697bf99710db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ab5d9a06562a89833266ce7ddb9671a4fd04c717806156d60b8b59c7c609959a59764cd67eb0272ecc5080648ca84c201f06e52b7fd310f16dd42f6dda2cb9c1bacb9560771a785278197b0f8df94cac7c9b9dc9bcb59f0b21ceb296adbff39dcd0b1c5e2034f1f1d6b46c04a818a29d972ce24ac978add;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf404a3c7169dd76ad920ff1a86cb55893c319cb4b8cc28e4f3cc25b0425d0567112fb6c2608212735c15a77a5dc5eead6320dbcf36f7f2ff07cb5cd098c961b3fe31d006b415ac8adc67b184b049398cdd5f43f3168fb0fe5d923b5486bf1f4878d21845963ce1a5bd0f573db3451f536e78a7ff4032fc0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2801a61913c1a945616672a489a435c7245c915745894bdf8dfd2994950a35322e401afcaeadbcab6c2a12b2488526303e091e6a87fbc42251ef6bd0206ac7953f97bae37edb6358c0cfa86fa5ad356aa4a107334c58c305ff77fb62a5c488de072fd9a48e30e4cbec575f546b064082520aba17043b8114;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc8e7ad5a01f863c534f0dabe67f9537f1a639b132a559e95c457c614b4b92afd27f8a332a12679c0c615a4411b494f5d1165ffe8f7613bd7cef1972d84bfdfdab2f3ed7ca0d9baff67b96294e8f20de0c19d3a84625247b7fbc2a530c7b3f913ca6f9e4b79db2c80c6ff18884f6ef4195197b3f67c32fd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9eff46a72101f04ac437d726860943c0dcc9ced4b024f43cad3ea5a85901bbc60a51efbc9256bffef7e57b0bbe88ae928a6107d409f6f41a68551f7d80d347cee5faa302e2501e025d0c6c9a1aa506d04d82af777a241d51832437da9aa4f15aacbca3c4c2edb3483ee1f8b8ae3cb5e743ba33e0b0aef83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17be2d88953caef36bd75c136000eecf7b70b7b3e7b06b2f4891c20f31f0f2b1420f682cf6861bd86270fe900011dca6a0f645bc976da5cadbefe9a5c0427bf05d3240163acaf2306835d247e80d09d8546bffd9e5e24f9299c04d0b78ebe8264a5ae4d06c16bf34335a5b850dc40ca2aac98d221c302b3ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1208855c64634fb227f716a19aad0ff7cb5de4f2a86031be89e496216f866d24847cf4125768671a9ae6a88d9f0667871aca2c0cdf41bd79f9a5dc6de53e5bf032864dcda1d1ee5c6ca9299d90439aa907bee7e6f361760351900dcd4e82c6747ef0ef6c13002ebdbf227498c30e754202fd260bae19d01a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aee4829df5f60f8ed0d5fd57501ee7118c538b4c822c264a47bd14ed39bc58a4e6d1b656a7b7fc7602f4a48e8246c0562569a47e1ca23a8cd88a281425b65cfcd35c40dd439a01db30b988f6812e67174d9bc9fd352db5e769ca17e606b446efcccdafd81bc903ce3e38d3ed1e60403714bb1eb97e452392;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h424ce48b2b9caad01ce06bbe39372e8ab4ca6c369dd98c6ede1fe8b3b38c88d7930a946facce6728753a354e6c31978b1047c900927c70db701508688d71724a8cb55f13c893b0b4116e7cd8b22528c5d705713ddcceb7d919fb97cd33a42259cc91e4f3036e3478f8d2b66b6dd6b18181edb4912f6e88ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e248d9366287597187bbdb09d7560caf704534151d3ba1ac3abc915498f51fc9e7044110f68302a5593e3f4a1d61a6f9f2bf73d15077e7a6c4fde1fa569ad3c0e8493f3051653855b248764a28b5e2d7009f3c4b6fbf5b37826521ff34fdc2ad709e3b26ef943ac36b65ead4faf9644121d96d56e8463bfe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94ab4fd715fcdb2d135c0ae4b5c552756510c2b481deb530b92b947bf43fcc51717fbf20b20f57c191f65f0c9d86d68434a683e1264052de9bfbe87bb0ad2fb87893a664ebf7d35ad01575c440c4a853de106d7bfa51b0e9093cdf87d4cf18460ec7c511013377f86519e5d42d5bdff4dbb3a8a6de79882e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a14d96dc5e2f39bf0bb2c1178498bdf522fb9ba6a8dab52123c2d10bcd47090a54be0e0cb0296300f6819b0c26466e580fdd6ce0448f3d504b308f2f522e927ceb2b00e4068ce7ddf97972c24b649f8229a82d5f719a26bc7b0ff3608f3caf6d26830fe3f12916d61c5557531d7574f836a120d441173cf1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d2a9ad847dbff478b9f42fbc8cd7f6df02cb0a661a020575d9d44d698e5980fd207d6ca50f963c0a8c00fb76f19d9aa84bd20b6a198583cfdea33c3dc987193bc7ef763ff994432d840311edcea14583a36e477e6b3d1d7bba749901a84550484c90de816e405499810fdc3d76d87f6cecc3f6e18ef6c36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef842fd919d60c5e99a52c5b7892cc99fb9788b402693fa1a9f240d5c9c30b51f1989686234e90103799e3f97d017f8d1f2cafc40d8d41642d64175e5de4c10263cad959e023b962706e7be5fbf123dbc50cb9f1ce5b949f4da09beede727314d151c90ab1de5aabba37b6d70c9afebfc42e131695388aed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4353c04569d9be2cc7617c6d7a832177a8273f650df8f727e8c53248aa5c7cf5c40e4b0cf8d4a28e0cc859955437e1c849c6fc908fa82abdc494c95ffb834b341d004292def8143b084c8b77d9dfc7a7ca8fa93596c5d7c02e58b0533252dfc4f3c82a1903ac44d0eeb59ac86fea67d8e535bbc7f5b41be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27e9cbd26599b2f5d5377c63687096db30fd5074ca4058127805aa64b03264dfc72ae28e6825db14551f8d41723179469511e2cb63e1833480ba86bcd90d12948dfb4a8419d3caecbf7cb5df54e00ba80bfb8ac45aecd32552b5daff7bf332d445909deefef125879c0a4dea6f97707d47cddbfe32f0abbe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8789350dabae83aeed3ef25c915c3313dc39cb1e4b7d04a3f07b2832889bca80c760a332434d290ad427299207da3312f2261590edd3290d4208013d07bd7014e40ded254aca0f37d8cca0a2d3c6d8e4487ac5451c38ced4d8a7c91aad7d21aaa98de7b612f5c38dfcebb126a99d197306cbca0a07e3e2b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb111892191be07952a18d9d360a1a33c8c9b69c37bd6643e7ca768cdb4744cd6e1cb93da3c553a3adbadfa14887b526f7a8f9d6a350feed7c69d61af4ac73b3011598e94b5630a99a53654004ee87f0b13f54376b1eb4bd782c24bcdc5ee32f24c9b6c651b03972e1d4fc272710fe69af8239c3fa1a07eaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e85dd0f421c4d6ce32e1bd3f55e6a7a49c271c655fd2f0e8654435cf7f87b310745496bd1ec49ee47603e488cc412db7b66f31436ef9cb72dd20d25237a323d5c570ae1531126e954f18b90cf4fe900ee6da3b4257d6fb03a93d9aa5501edda8f1159465ee9557a3971fdbdc1a4edf2b1ca9ee6ca9e68d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c5f8372b1d8a13630b5465d648bf542684aa64cde0ab01cb06c8ed7f110786eae3fec591039fd518c471dc608686e41b1bbcbe1e936991559a4ab53b4009385e28f512fc0053a3cf5fcebab5ec78fd2efe7123bd7ea8d55e0a0064db33178bd5d449c92cb3a62a2ed356a090c0bca2a0991333157b5dda0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ebb48dfa78ce0b8baddef21f9f6a2392f613db49d3599231e37663f00b27d70b140d2df1439750bfb7674b54dced3971b4cfb27e9238e1456a474a55ba0a73116ed9e54307223b6c347776051b01cd7a250b8ed88de7122c71c11ba48322be149d9e4ceca512235a0e853f0875282edcfcde0fe43dc6879;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7aa4feb196c5999eb2defb695d6701b2455ec9825e33350cc5e5fb946077c6cbb670282663ba634f3613414a7dbfe884ff755a93fd2215dcfc951bf118d93d80e6719bd3ce57ecad5cd7381deb6069e4a7820e79985d9f91c39d6b16efd2e3543b0a36eec8885ee802c96c9c7cdde7ad7a6709d2f5c342c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h885fd2e358f4a66060b988c775913cf1163b6e23ec6278a1e2561c5aed6d62438b5beb71257ffa7ca01f185ee6fe89c0b1ad299e5e87fbe47654d24164dcabfca1459bde2f8bcdff7dae480a8a65c2d8ca9d508062f7a59db0490baffc27d329a47be6a42831329b12c64b2c22078d9d2e481fd3b8b0a9f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179d65e2a10093b8a42147681e7ffc1f15cc0a844c3c8a9595d9e2aba692c498aa432993662c659129ac4a9951ae287f77e790ada863243e357baaa5798e0c8cfe9008eb68310a45a9a21382485c7036a01e5b95eff0c248da57ecd7df6194a75e84a3c35023db89f1bd551e663aa0b219d2d5b12a24b53ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d20e3a77222022b79737238c7249c49c3f0d3d22da130edc0b800dc149b632296e6f0454f46e74d151fd350152b637ad979382165b91c5339a6c3170235f2c0b0fb54d9178a4f92895a482fc7f6a838ebfab5ae29ec877e2e41e70d5f0937cdd8dc93c73951273feb91909aac8cd3a2f32a86f97a2aa457;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb7a050e97420fa7491233ed301d3e40302e197e64ba53065686b8c21013bab12643296745879ab4637bc4f3e13a7414640f0ab6addec7adaf3c4ea71e649f14e8367423f9f223d5a22a424052428cb0b3a37d2ee1c04e56d4830ba58ec4654ae7575474cac2a8b5f8fb55e3147a918d68b643476abcb654;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d81c671f9e189af1d6f18c8ffee7066c06ad60cf741c84a7aadd48ccdda8ec37fd33a1c3552c52fb358ecb19530dc4db9f1341e4c2442490e8b44fa270f37a43332f1b2813db41cbe0490219246cdb133c1a35cae15ff5f18b4dd906f12f102549b63fe424886bd835350e7eb1a6d443b7ea7f798c2d89f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cde7478cbc2d3ebf5e1aa7115863cb0be698cbbcd9fadcd9c607eb2430aca3698c8993458fd88666ba0e5037533da40a3eb9e4ff922264387af538387fd8decbf019144f341e113c42ec57d368cc6c3986b69352b913b42bc945e4a9004ea4abeaad4e495bcf6337e0203d7fcb36754c045f0f891c3ce8b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cdd3a39f6d13045e104f6e659c50de1f6bc5d82d7c79830e100bdc3c4068cd8dd15dfd1ba28a87098ed49caffa0cc1a535cdc4fc3d48cfba5c49117e6cb8edd107a31a4140e9bf37edc0e9490d4d9d7f584c704ff09984842b5705c1c8718360612ff9f014e8d1afe28eb12ea2bdbb39ef1dc87b3ffc7eb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7962042bc034a85591dbd27228b3296ba9ca343ea120f1a5169cb2595f641f101a00f5d71b95bf4c843a4b4da7287195832b465cab8391b1fa0794e310a10fe3ce1a48592eafdb3a567e6a3a72a8ee684de0f71b74c9b2805ca531303a70e03b08a062c88ccfb7db43bf5ad970ab783f7fd2ff7ba60d9fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c9c605d2a3ff7ddedc268ad4587d492d9cb78f26a595edaa54728f195a013e77b23d79cee851856662ac1caeb55d81b61c3578ac498caf2d8236d27fa5d1e954b3df2e828757df5f42c10f7827fec166c61e6200324f020ecf7be8509ffd6fe11420ddd305ae55d472e79023eab978cba8278a8906ad50d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b25dfa3972beab5fd3ca86b6acd4cb78a37fba23d811bff99910a4b74b5715f75644fbbb6b000a0755dde7fabb7638ce82990212ea7d3875f24554ea827c12a79275ec7a641dca221b98b31854fd67b2b4e7f833847ecbf785ba72c684782f4c0d05d05295b146f7b69b5d94650f31b18a6ae9faba3a088;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde9a2cae25f9c3ac0636e933f82b4935a5b235546ca755660315469eeafe33781fafd9d2539d0d350b951c759b00a29b4851fcb98ff876c8e506f0bc30e9b4ac53cc89962ac723569c3c6b5515d61d90aa5e0fa9c6edb9a6b37f7622a6c1ab1f6269786b31a3fdfc6e391780af0f8c44b692a2e5c589ec89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd066988883961e0904d0b67d8021eed6a2e378438ec7f33b55099b2fb29d7eb5cd70f8c5eb98697c6e6eab5ca8f6220bbf5d6747a5ebf7cb834806cfb5e8c5b21bae3b3ba1d112e18934fd150328819641a9c4eebf03b57a6ce3e95118ddd659b65fc8caedef6656dbf687db8ffdf9b293f01ddcf67da1f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1300d780b304de24e2610379e5dad2a7cdfd7fcb5d9943ccc40f43862c30f43544c19b5b8ad149042bf21632a08f9d38982a76d26e20502b7620ad1967bc4a196b5a96c79f31ef8ff728812a97ce5542463accb442842ea3a25e153b667c1a2ed8ed8432342b4cfba1612dafc9e77b0e2efc70154708843cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd3f2111bbd5e4c8ddf00ec92e29ed663d20b72ab0a96b00b7f321624e18804d2b1867f4ae147dcdeb36feb50ecb88132a2813407fb70019e41b3efd6a440043d63574d0f99d9c3e98055c2d9cb1ede0fc1adea05eeafaf59718bae6e667c1c2d94b7966527317a0b22cb11bda714241bf0e7176cd3c8831;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61272726637d2f2ea9de94a0b596c9b79c484e8e23a8287c418d7735019ea46e4b85c29392f8836c0a89ca4ef231fa2480db8da18a54cf8ca5b6d92704d18e18988529f59327c26c7c5d2046006e465ca7224c1e06ba499af1b9386fd6cd00034931ebe82b7a32676749311b3677397c378d7b0396ccc57c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d7c2eeeedacd52e74ccfaba58416b10b450f7461e03d23dd28667b653ae32810fa7c1296ddbec56cf407daceaf9cc47e9d343e491b607ee1d90be7c9356b5f62c26cee74adb836a4ebabbfff8e570a4e4b368e23c7f62406a8b196923808e717d837d97b78a21540d1025b67129fb9ea7237e2665a8ccb7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h527ab77d9a3e90f1bc0fec7e2ff44cfd609503942ddda174c5c9508d9a279210edce30a6f255da212763a687e9ac167286d5ebdea4ae24a8de5e850578165e6522894e7f209183ec52eb729e790dda1cad29f0cdc3dcfc872724cc58ef166054124fb6b287efd3d56937a7210e23de6798b0cde1fea96a96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59e77b277e9895b8071ebe47f471a18b40fc7ce3c60e4d79ea2e44707174e091db6f8dbf6f675ce666174a45a609afbad406a9954a52c03a9231018625b4bd1f5e4f3b4ae79ade3f2072a5584236f1ba2491861953d7e97fb8d25f24742d9084808e434f3f1af9a96797fffc2b1fded20cca3608d5e699c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e2ba0fc6e0d40640329056904140ebc03d8a1eb7f7bc679fce0c3b04c560327efb63ca200180c00f3656dc027c7396451acf91764ddfa98f7cfb6431d0b7b89d46f9df095ba08cdd1f13432fedb9575f8216233cfa8b2eade3e20b1d10dd9aba16b8d0ea4715474ac73134d42bfe504bfb647326242ba0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1a8015d5e09642ca27ede80972db99f090bc4aab484adf325ea4e5beedad6b761eb6cdbc08b836a98844731169448798072be86a165fa46fe483e35f4bc50bf9b9066cb39855254e5c9b64be1637d98d9c81861c74ac78879bdb4222e16e91583686f73c0a744e4d69960b17bb8a5a1ac1f14724eb299ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecd8ffdf969f7255f3d6e039a7d6fa51d2ea9b8d8e181e6eb6f23e8d0a152a10041a82790a171201f49acba9fba98bb1485cd3123174d99c7b940f3cb2f6978c0da030ece34fb33376a92e9d13bcbfcd52249cf5d5f2854cd493358de64b79052c69a864fd7dbd52275426b604e6ba8c246abe2efd94751f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ea1f789217156d4ae82a8c9e7b12ab308d8378f22929e51f89c301506987c2f4410d035b7b1737b3578bd1b365a2b9bd27d486931ef012f2f0cdc88aa3f4c14991adaa9b283f9be40d88f0ee8ecb05db82ec61d0a9ad90b382a6473c97eee88d5bfd35ce8a40b92c9e267dc3896b2db93820e0d7142699a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f463035c073662dc86484183b4349a0f3833402812793b6af8282e069e2131e3b51cdef36e0accc4b0d92304792752155f6e30cec741706b4fbb0c41b36b4f1ae537d42a6580ddf9dc656077c96d5aac9f74cc114b25ad4d5e75704e2b5ce303f0f3a893d430f1c39f6e011f440bd2334da351d70ea8900;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0813df708d8a8da83bfd86a5382f75c6b9cf17cc7dbdbc8cad85023aa82ef2909e2fa4e17da691b8f0933e462fd3633feb0b5cb860ef4053309a4617a598783f6eb634b2cc9bdc267e9790a75d1641221d48e47986e8b6011a6ea5d5552d287d55df86c4ddd8334e2be56489a054097a8a97985394d52cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1698c24d7898ce652b879a131c5944fcc085403db0fcc44a3fb7d86fd7e76cf54b19915ef374c6ea63599021f36506216aba2795cb704fbfccbf53fb1b439c6977315bc07d7f1b39306595e38287af83076e4c4ce3b0e4ec300a42e2954b19547226211e30a83bd0975e152b6197ea69790c3cdcd12b7b8b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bac9c9dba2d324de85ac62f127136c2ee747f92c6fa3456c6953515bfa87d123440fe6756796ff55b66b37cde6cebe8b06e81321c6536c63d9e3548f789d2834103c7641947ff2f60e183f964530eb67b5e3fca4b305f24349b886d342935e0fdcd4c5c50a323e7b5f9b04fbd330829b93c3cb2861e7d040;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e59b2a870a0cd9226d29475bd3d366f9157f3434b9186aac023f2312a492bf02403f227d8e5f464042f7c31a2c2b3982361e8526ff731d18bce077c5dcf568a229e28eca90eb5bfa3dd255979ccef1a76c109189015ed9921f88d5c2ec95c1c8d3b83184d49c8dbb33b42c1bfd803c3ae8901d68fc3aeb6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40acf26100f0e3838d1384ef6208df7bd7c70922a2c11995aa0818d83393ef609bdb3291ffa793618042eafcdc5e797e661289929c74e0936ee1e725b863f71229943b26bbf3f6440aced6108ae62074b0052c7d24cb639b3a8732aec9b76dfcfe849d8676dc2ed348fa99fa72b510e26548d9536893e02e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cdb001f8b4605d1aa9fc11f396dabc941d992411399584b82903f1f94c148d7777cae3b48a39a4aef81bedefbba5681d57124f34c5174a716353d9a7d5577b063be7265613dd77d91b1c9e95e8537029d72800bb730b70953ba62c6c8541d35e0a13ce382eeffe934fbfd57994559a1f8102dd1f466fe15b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1894d366715548c50b9699d61f42e2b2cffbb9e90ec4f6a5995d9de9ce3219ba9ee755463fb487a7d613c055c12df466f9bc8e087e68dab969219552c30774e7f5382d51d9c1577d2cd0d667f9e020bdf110da306b1a36c760dcdcbf6e517eaf1ccd0d2ebef2f090b0f3c56072a797ad41a4a4eb6b0e79dc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4e2549671cd7aa89adef7c6c8f128fa6343ccdffba3f8e33870e7fd46df7622a87d0be78497593983fadc8873f7423694301aa15db6caea9d1b2e9219df1afd107e0bf8667722e3eec987c92b5957d83191e07835fb8ff0a8bad2de393d39c67de4a25d0bcf5d9c6290550ec96c2f8cf853cc755620ef7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1921a5bb49727c9427d3dc3a5e8b1df4f56b49ada34058f58440400af2803a144b55db7b46835673dcc086d54d73ef3d9432defa8925d4a4c1861eb1e7fc9ff79a2e44bb1e4e986bc496edcff86d6fcfcb568f2ffd480528d0cbe5c1ef1d57f5ce11bd1ca6f16da663e0408c1ee22843f3a364ccbefd92b42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e2b80b9a34a78f57b09d87f6dcd956390241c9e827fa7987adfbf6e1b206506a5e34dbe22e146eedff2b0ce208b866d74b17be53742461fd2ef4f697f22cd666d3f3146ad9f918905815cec1657f4dedde9cea944eb52aef8bd99e123bf6493c7c8cb6da0da53da3281964925af2333e384e73a7aaf1a7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c58f59115c4e74ba666920bdd4a2b1cd629616da113b993c5bce67bd8bdd1e88db9bc37460e0bf522620300b9cfcbc96f84b70f36f1a4de79d88136986ec906a797d581ccaf69ebdcac96b6385e789a36fc9380cf9574c23ef615eab20af0fee3209bfd865b7dc94142c582a1f1b9f67d02fa2fdd3253be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6d3ba75b5390f1cea373d7155939afce8b8f5ac34c79c21b9ba6250e124065c0dbcaec4f6fd9c056d311ae3eed955c3bc320cbe1716f5d43363022ccec67e6ae5bfdb1c953b0029ff6882a8c12a8fad94eb6db5f3b506570e539dae51ed3ef01eaeabe6906610018ebcbaa12edbc7722950d47acec09510;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2cc4c960adbf7bb5b170527ec64fc05330a2369eb44c17ff16edaf2157f03c6f4d7258ca662defa25d5d3dd3542f2b9f54c2f6c02ba2258f9badea6495346c1700efdf682d8284e0628b48087fe0054faad1e245036adadc94738b4ac139ef8a66969ca22a4a2c5bb0a854be1fb7472301bbaf488fb50031;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc7e916495af04a4d368529c6bc740fbb9a1383a7fb34c90a085119938c57072a7ef05e35bf028cae6b5d673b2daa15409d1bdc03b08854a412b16447a09c40cce347c2a8ff703f1db11e04da843d4cdd93ed3536e794d623568bf2722e7b06d56b13232b23049b395645610b101a4ae5b830f058e55d5d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddd95b4fa9b85beaf5d435a4ff033fab4a9c9bcdb60d7cd1737d9cc9e4d79bb6f02176f5ccd2679cec17c5711f1c17b3aa8ab4605847b474aacfb794d82a5d030e216636556991cdef50578495b3a56fa88f82baf4b596d0d27761a29c12940c8de400fb576779bbeae60d417cf28dd9148c326ba1b1b227;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ade650094485e439789edb21469f84ad7fef37afa59d13981c0dce60ac46b5f5a89b0223233f826da501f231b0c17a5c78057c6c3b723b2b424d80ea66f3bf083f54c2dd6c7556150eb26e021ecc41b331b3e59a87b80017c09ad88ed77f7e2aeaab1857739dcf190e204930d151c85b9ce021d0d0def85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e8afe65703d193b0a7b12ca3e2632d8fdb41a06fe2c0c71dc9ef13bdd2eff32f699d9b78a2359c3a88d2dc8de328d7873179fac17b6f34ae137235922a4a09cd739e2e5332e085e08a353d3626c585962ae8b29efe25027e1fda2231fdb7454adf7dd899ad39b67bb9ed5958ccfefb88de4a0b722fb0698;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc351b93d16b68badd349d8dceea41f36e1c374172f1dc3a56dfacb6ffb0e6efe8e52f2eb34382bb06bebf21773f21778515e606241c85420ddee819f17750474135ed393324f51181564e6d55734d27d365b3fb588c4ae83a495b251105e473788ce6b50c760279981fec319488a63962c9c6aefe00eb046;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1474504e9fb2a8af73db31d4ef9e21cb2d47abc1ac200ca29e6a610be89bf24d0bbb9b4798804753d90a2ee9ea80d0b0b2ab008ff0c3461e19776b5cf4262818987e59c028bb0ff1c8f6431eb992dba50a11443ff7c77254603c1b7591f46e186e192001b983ca9cd20ebb1e6c7b9352b6d49f4f75437487f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda3add41a4dc9de7308bb6f17b88f1bf13d88408041fb52a8b00a677186297a0b571b0e68864cdbc3fb5cf227334d648af9adf3bf0ff197c8b9920268b4fca0c1f55298b401e2b5833c996fc4e27f5c7507728946942135feeef0cbc69fd77df3307620480cc11ea82fbd23231bd610961d650434ac8b072;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15976f45524fb96797bdb5a1329e865a2d8586607d98073fdb890a27fc685d4e6f760ff6d6009129e718727d4965e8a3eb5c34f914a29c9614a854d078ad58847e706ac89a7c3584c43f0d55956eae995c298429b15696557503b09f18ce530a53cd3213dcff6795ff1dc595820bf3c8f4be3e228b42f977d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1942a7dd9591f96c899be85237b5a5c6f6a0a507d32407114a3aad810b0eac74d72c92bc27590dad73ef63f928aa9fe76fbd681655826c166084f9fedd47013d4edc00bafe560d3418c95da7d102249f68957ce2e6da640770731e2de124053a690e5823fe9f3902f5ad15f25303ac59cbd29f59f1c148ed9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38faeec04e782cdcc1c4d44c2c2286880eb0ed5790e2667f9733a6ad6517d5c847287a913777e1859e95262727cf9a6c80049fec185afb4f982dead6cc74a4136af1a687b1fac5c3e00561d0799438fa11a97e10db1cec3c53502dc26f09e2d9b8445a191b01e637d374d6d80680c45a93624af1ca47f54c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd25f49b76e6bf754efd24217a0e41540a1be242234730bef968b4124c9725f19c2498773938af8941155d3e239aa63c9ab8925d5670dcffc9f45368cfc1177404f62c87ed1d740f01f69d088ab76acc223610505c6f5e072cdd7d2e940e97d40bf6d0cbf43ea1835194e8025a4532ad32c5fc0c383f843e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dc95b6013416354244d661fbf241d08d3010b2e50719bd2db40a591b70c42aef9bb0e4e340d3cd1688c04c499c15df51bf4b9157944aa2ff045070ab9243c32d28180b0569c17b64b5b6223620cf0bd92c8ea83ba4c25089386f50027b653611a40c10defa7b5c6096a9c77dd5920985792fd6e4a1e61be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190ead4c1121ae1ec25ab0f8a3a7fc832f1ffef30aab97ab287f22643c3faeb7456fd493eeaeff471a26484ba85d0f09f75b36429b9a3de7338c1088fa08e6550f238f00686dd86826bb5439e85afe4d2490ccebe1240c76850b2a178ed769684eaf14acb2045e611ef6e46f35269bbd17c5986f3218c2a9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfd31333552172ee3ee24762c434e8acccc056edc57178af73373323f73645f6477599920228370a59ace6c485641a5fbe4a0c4fc4ec89fa9b98e612c0888e862122c1a76d133a3d0307ad8b33c9419c398c845c085228ba2257dec6c4598dc6a922543c2be9900a4a6cce0b9a1e2b1173497ee1aee2ce84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d30940cdffd4fb4c6e09145e83b6f29d457c723824d3184ee1524121bab2f788f3dd2c78cba0b66b94ca999050cf026b8ae38a03c1d53ce5167ac50904027b12a33ca6036741f216929cac02a5cf8264e9c0d5959eac0826ca2f961ba6ff12840bb067b72d829850d49c7228f55ac13319bf4b9621811a10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdaa20344f698d011cf860fce268bcfd20d2dde1c2737a164d9f4b27dc36845c36d2ac9643602e8560cc4ed52dccf002a6080620a6a7122a768290ee517cad48732d8aa585f7de805eee6e283fa66ca9dcaef985450bfa633eff3d70066f3834ad5468fca3f7516fb3f21c52ca93c9afdeb338576b30718e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a4133439e60ea8adb0255209b486888452f0d7f43303c399c3f6a4e0169d12f92f02bf9b19ed2dfb958cb67e465ce54c02db3a16a4daf716f399002bf53a8764c62ff3b0b1a035d39422fa3f24f9a22dcc0d6ccfba4a5abb20105824e9a4c3853250d8d78d8b74c81fa52e34de5041ac5c605b5c99be36e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d96b408a1a5a2da5d7e008f33326a7d171f664f20f4ef85fc164f8744cf1dd617c0242276fbd05c1c6ddfc5975c8af843344c70f3cbb0df220247a9658c42902158625ea40a8483c460fe14782d1068b8343ccd37fdb73b7eefda9e14e652646e9509bf84566ff8db378afb0918b6d4c66afd466b268f6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afc4ba0f4a38a174fe251bcc57056f93a0404b2bba20db7936519338ec34d03f07af4bed76328389ae1b32eee06a97d9576d9c38aa68131ac5fcf035685449e9db18c9da4bd21f2b4b6168350270de5c24aaef77e233bcb2591c94b6f32747152933866bf0cdc133bd9e6e96c3a631f48ef722936857ccca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b940c21cd1bcfb69f1be8a4f18e5126faceeca6036bf899b7623c93c3762e98d9db871c685c50640104b8509539ba0e253baf0e906a0ac198149cfc85dfa0ddcfa811e1a7c979ff2d43b81423070416eb1049705b06a9903bf5e46dacbd843644122b6ae809f3964d036620112ff020a38ae71953499c8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21d11fd234d0054091bde3cb677fe34908e7fddab744140cfe4e73450379a43e6e76c3a58c7f4cb9cba2b0091f0d14cc7e764c6ccad646aa2924fbf9ede803ea8a49df2703c0520433c470586c46979afe470ffa386b0e482bd7ec0fea018f65ad04eeaa9cb1d7d09ec918761886e80845d8c4c2752b33a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3631511337a301cf91f227d08d82c211870d169d9b51147bb412f81d23c47667d6624d312f3faa8e932ca72364148eea80f37e02a0a2a3792a37a8e17da14a8e407fbdb9df43b95414dc2796a2eebf0bfed7671352eef6873dde3d4b59a93a8ba45666b2887fddbc94f180f33d548ccb29f7415d881c0c0b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b1bda81e0a9e33d29f544ba4a78f3b4eddbdab9b0a7a09fa193f51974371574de2f7aea5c6a7500c9da238c95d784c5d839c0e5a7ee45b9af1ddbc06333c9ecfe3267e480fce22a7e746ea47347dd6264fba0479ff11e909b411e53e56f03d8c614b8309e83283bcc3d570d2c7d41cdf1ab83b2f9c97b6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7a89f34d46c8d557f4e07c710a40d6a13e4ebde8dbd070463d5c506319aaf4fd339fe806415da16ebef865de4f846284bc3f6212c7f5230b6b3a32f5b608bddb4af5bbf80d62938f7cf6a1ebba181da25cfffb74880d9c61b0b4edfbe37ca3a5d5a0efd30c70002db2be7c0ac7d87d21723a3819caee033;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11edd7b6758e51abd367d5afce3ef24e3208ff4835cc52240c32c4f4fa5d43d49042fdc6630637b74ef2e06f97d936eef9e960063819466730239110ddcf2e8821cec0cbfd9e079510f0d94ed11f53446d66cc79e72ac602836cabfc0381113019f88d627bfffadfb026e972ac6cb4288c8fa1be8a19c5105;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163a0e9256a8dd2404f51fd32728cf037cf8190e97dbaacafdf40f5f1c1f898d5bf5b795e02d079483296133e6371d5b184e7dee182b9ee94f33869dff8ab2ed030816d3485bcada2fae1fbf176958752739f9ffc6c002ac51982746988181c55c47e5cb2428447c7ab6e8cfb916a4cf1c1b3f845bce6b9c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e031daaa62b5c8c36e835a08ee8a824acfda58e7166a78e24c4498df2067f0e474f6de30dc7c51d41a5d873d52f061cd6ed23b922a720a80c98312ab9f48afff22a14ca3f7690ce29801a9dbb4adc627c07db2394e8290355851c71233ee6c42ddf23dbcb5c54dc8b06227475020371f35680d5962d5624;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133d56f8e1a1596b5ffebe69aa71dd4e243c3a9b1973844fe482b1d5c42a49d99ed16f92df5693b9c350e27d19a19f22f938d0214a534f8d9cf780d5c7707ee910fc32ff9e80dc18fb54f2ae58f6ce8189913783ccdb7a06eccb18128830e0b189e3e8b102fa2eb160aa41c3eac42fed0db31dd4ffa24ff34;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17631e084d7021c6057d4840cc138e32ff02fa9627d7a855a8a8397b9f573e86ea94bec28bdf28dc72d0c52e2f8a2b11df4bb81d89699e9a615d352d36aa23469604bfe507d71b817467b775ec7d6aacb128e87fe48babdd7f9eb52c4ab8ee15be5e8a6e136f5fbc6bf7543fdaaeee8784e275af66223a83d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b39b4fa91a17575699e4b3b0bcf33d4005cd188687b1da5901ad45b6a00c2b6335d3d9c728706e397d5573ca8510a132e35812a3fcef79658bbc90572febcb66c3623e3f6e4f76772b73cf75fffed7c59c41d6d52cc14f38aef3829b8b69dccb54b16597ad096ee0d7fd55ca29a0d9124d0677b048ed542;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b636d0076f521cb7a1582bd26d28aebed7460846c42a35ca722fb29adc782e78148a2146bff04315abaee260f8d2f5abeafc612c45cdc3c533fabad1f331e6dbe9934981742ac2887b4798f17463fecbc19bd50da4f893b1925803d02ad6b4a53daad730d8011cd345e5ee03597b2ea1b6b26bb93567466;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49043f81e1ac7c44cca2f0629d2d59721e31bcb6e3d237db9bba90acb8caabe31f581b1d8e3c8bd099edb5387cb6a21cddf7a148c4e3b1832e8f24b78d34f2c975543f256d8813c3c5246445bf211e33f41105a3f41aa270d1484252322b464c17afbc27a77ef9ed8b5aa509015ae3818e5148ae5007c95b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha002311dacd212c99d86285497723a1fa9657e16d952f3b9b049b9a39ebd80d02412a6b3b5f3ce7c6a8366838447c7cf0e8032c0e309083aeddd3b59fa37c2ed7be1992f8ceb966570e910b45def3cec6507294059f9d6606bf3ded78e8428234a503c83556f7bbd110ad49be5216ee2036d6c4f561e9e5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habd67332467c2edb2e8d2615d7d8ff2c1d0671d7b63f94b687d000f22973b89baaee84c083550a248a8f96be204fb0c2fba88c374fdd0bb6fcc4b224b5486afb4954ec4f25ecafdaa98926d85e80c89385cd1e98acd2c5d8ab6da798b3a8db6de9716790a13d6133c00812eaf19fc4266c9dd486dfc9335d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69a2e1cc97e1fe65053dbefc117482d391c3407ba15d30c10199d96094193d474c5370f6c331044f2f67c701dfbddcb80885281732364d58048b0d06fcf449d72f5ad067dd13dcb83993afcefabf1a897393e0cc9cb4f0263063f3d50bf123a8f1ff73769f0b97498ac3c86c5728b85907f4420406998ef8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1e88f64ab538e2341cf68aca3dd21b64f306fa0ea326409d75ae722d969c767db7078ff30123a9b635585eb9e0843e6d6604ae0e024f9600bbe28a2dea550f790f8b325c813b73c80198e35edcbcbb371fc58d084e1493ff4025d88ae4821ef4dff9477a9ca6144e2be5ba92382a644d16f490666c00744;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8b8739f1350d5c9f342e29750bace986b51d824e3a5cbd40c0829a121681c3cd21392eaaccac6852232fe65860430f3cf6a727f619e7853739503f455eeed994f8e11b5ec04dfbb11fa15b4d6c72da4fa1874ee723bbef60d366e7b3007a6adf8b1a760068e423841bb5ac5e72a114ca9a612b7abe8d8a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1133b45d5f43f4ec6a7dc9301cd92267b213ee55d1a71f32d7b99cf83a8dfb9525a5c230fde29b671dc04bcaa2397fe0f3ecff03133a82a04bca38ce42ad856f4c12147f8dc6425c90a60322c2d921a0a143b5a6be68931209b2fa7e385b02788fbc761ad8674ccdfa1036aa2e4e4d2b010dc7b1027001cfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11daa8ffd6dabfa68c5312dd5670ac1be4ea9f754e499b06bdb222df56ddbc33822c88fc79e59242134adac181a402cd4d3fed34f51536ad71d73e34fe7c6414505f48e87db3b42a1fecebc347b1e0a563541ed5fa9a6e4590de0031b78cbdc7f1954dfbd99e42cd14911a1c5ccd0b81929bfdf5382758767;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc37e695832300f55bd761c27f646977ded6c62467f6b5270b952319b0238346f19ff8296024913a8931d532180667f44ea66887862022415c23f14e2185fce4136b26eb578ef51387923bde07e454ff3d80c8f0d26d98c35cb243da7d2a916699d187d3414f0333a3344494b4f5ab82ff8a6ed0c025c703e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1435c6fb982c71a6c1381f9517bdc918b3d3eaa3207f9a7bfc48e49d72207551e380e7b0a41c1bc421b9d57ca5c9b223780831ef8a047c0c8c18a7625cb2712a44c4d4395a564b85dfb085f3d0450116b07f9d049a621f64c5ee6b6e6b13bd800ee36b315a1813ae9bfd2d488ef9181e318b62547aa83b3bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f61e8fedd950e665dc0c7e65848cbb1df5cf62ed616c910ecb13d134a5938f82992f411525a7a31c99daa24efdf5ff324d3b57512aee8d740fc78683fd7d6106bf1e48d90a362ee5bfbb17b4d3fc335fb4001965fb974f33f7fad45d8db62d97077775771a17fd59aecdc1a16e341f2c46ca13a16eb4de2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc31a25011c45799f774974b0a5a0d259bd0a6e5c79cccb9c76fd58ffae416921cb9cbfcb5405414409a3b35dc4cab5b8d4432ebfd57e84ec8fc1662f8fbd56e23ba5e7818b951a81595b2c4c3c24930cc858beb46ac5723a498bbce2448fece5ee41a40e6454214f407c30f4fd7589f9d637b7948ad05c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h750ef3f7fa673c9b50263de436ddfd758ef8a8c529114948ba9dda4c7c0eb67161a53c33b6f07e6a3f8433ae6917aba8effe2efedff973f31912c76880c9bbd9a4335304fdda131e1f15425cdb0a6866bee42bb6aff7c95ddc1bd871ae63e4943e883a1c21f641c910fd76b015ae88012647f127be7cc5dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc57ecbdbaef6dd7c4c95d3e6198e925547eac5cdaf163b51500170f0e2017963444a36fc7fad82430de6499562e021fed1659536fee84acd7e79fc2a682f14aaae724aae090f655486c16f9db849c8ecbbb4b036e2be554c9082c6787af8f62893996cda386f03935245f5b6d81521ab8d1f03fbab3b1165;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bd2c25762a37cf5c6409f39a8e446e5dc8102faf1f6d559b980196424cae408d898ffb76f061b9448986907141dbbadfcf2bd5638eae7e1d3ee4b0bfe1b65b7ec0f3fbf41e81766b9cbca57e89f1f9237df5c0a4fd57da8769367af361a7b8d2f7d7732e8b3527fc1349e5234ba36e963ae2b34374a6ac8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h521e6813c0bb5cbb1e9653333e088357ad782c88ae297ad6098143732d534408b75b3c76f291dedbd1b60d78f22335e09eb159634469cabd7e59a1bc80fb11ef159e0beb0e2f669c18f633b7fea77bb9c749df371dd0cf45d5fb51fc1737397ea33cde69470aa334b5dda6d7fef395cc78415102c5b85fdb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had5a88ce09ce49eb6dbcd386daebf531e1d743547f385f45e17d73522192f41233bb78efa71c516275e493e93f2a648c7a8e865d786fdf4411c58a0512881e47f5b1de72533a1c426a972788898fcfa78871eef814642acad0c47d67c9cc0c15f4162abd6c820e92d5405468fe8401c40f38ba5428bcc310;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18035c8d0add4fb8773a5e8c1acf81f4b83ec472968ed326d4ba17b69ee1fb9c0081d04deb68171daeeaa90cbda3e6f8bf6d0e89f5c68b39cb9ed9ce46c07846ef85cba0b7576fbbbba74e59818bf9a019d2c2edc0b51bf49e88d91fbb1d0dbd46f66f5b9b1cd49d5e03d680c5ced1482c6ce03b013de7d03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137f2774f496cefa8f75be722281d27db03aac625eeba9e6ac18ff138f7f5257a2b036a7ea50d5e844f41ff4194309cbcc6e2ba6a4789c6ebc3805631df3d8b568a0a47773c5c6d38052f1e41c3e4cd5ca6ce11e1f5fab38654bf40b3f1681d2d05fa4087612616bbe8f9a40eec82c19893aacbf2245c414;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2af1b78720e7f044748e96e13826c5cbcb636504a70ca5b64a33c598a1ac4b411efdd9766a0310d77b9669397e2203dfc6629eecfbb2bc2da1e05adb544af52b62a43ee93d5eeb9b1e57fd7e85605674baf0ea64216163da92c7008693098945335fb1f59f5c026977a1d8687f21a0a02aa974f3c924984d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3d5c6a08ccea62320a43a7077e5bc16e3af8a10cd5ba9865f483f0071900457f59e94b372a37194cdb393d56b590429441c4d0fdba2969ea4b2218d9c7e60b1b0dc751f2e4c327fa3530ccd785e08e0b4c466f53401761477136a71269fc56bdbcb9144faeec8dca5dc65a79fa1195e10fe852b675eca51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20846ba19da392581349317f437656eedb9b5909da912f66df49efa5e9eff37abe7e652c9ad8d05835d987a77069881182a31e45c3ccaf1e4109f016987ba534ce1365d597c6058fcebdd8fc8a3cd10003dd20bbb1f42df39305f3ca4724b4ee47411927d6a44a1aa6740cb77dea04a75dca4ba2d569d515;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d329f0cfac6d5bc73670a01aa4ccbf59b4eb1ff44fb9a9522ea2c8dac5b88fb456bf080c72d4019eed97f1209cbe8f40fe2f2c29e5429991798b2a90a5f425bec5cfeeead14a1801738312af86f29781274d796f690b8b590c633b73e1c9702dbc3c7e78cd1486ed33d1181f3dc39b45a17ce989a79748f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12715c7e98b4373cfb80e3cda71844ba5205dc1f1fedf404e38d1384aab905c1aaf42d9cc7a52c21b0442adc072f4cfcdccfdc2260c1636f1b02126f0c8d5911e673bd8f63e59f0b8f96c2cb64d8693804a7e299b2cdafe61472ec29c6917a9650ecae2e7dcc59b39a9534e8420386877541d972eb9d8f9f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc65e1d177bf1a5b7b8245b503f4fbc0160cac153072ef94f4c5b9e986bf1c2f920f87cf0485f244847368da47b442935972bdda9b2771f903af65702c018f1047e9d5d58042dbc3742fceba46241411e85075a7b002a821f35fae85f5d2f799d7ed0c42493b4d6482821a8c68dc68df35b912d0a38139bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5d34a892ae51550d4a2ab035b433b2f6a20f530bc4997fae09fccaf6c1f9167b31c1cca9f9e239c454b495c0143b8d1b4b31812fc688af958fa60ed9fe6a1f76f920eed687add15c15cce6a923ac78354e34410735041b76f511e2d4f495344a6cc1136249df7f3c1b508f9ee9808334dcc4d663b36adf3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49451ee30aa8e0caeaaaf9e90fd78d18b93f3cb5e5665aa35ca158cfd38a6d5663b1fa42fd80b701d2b2b0f394baf3358b4bec389a50a5f5870c2b36b02729ff0ab3818ecb55c73aac9beae7e1744ad3ac675ad2beac3e53124cf7ab781a638aec87aaa730dc3b31359732965018934a0fb4118bb7de8752;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26a628d55d407ed0b2a05a0afea919723da65aed7b6432dde5958aee680e5c1e29a8377aa4c6bd50b1f6fed9002f0fa718b7c5f927769e3f64718b2b644f05f49bbf7a5651e34c6f36ae017090767b805581882d5ea0646f8630d77b67cc77d5c700e0882ac65f9f9f135a985b665c33be38e972096fea0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58850163cbf354668d37a8cdd164d1bd32b023da5d9d6983e2105e314f5f7b5edd62dbde6e8b54fa8cc9d3bc8256b703c9e724fed871de123825fe5734adb51025ed22ec659ad9af9fd4c3c0886c96192f1416c594413b36643d829ed92e5018deee8c1c986f120b6de0e5a0139804d0204d5be41e0acc57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13572a464850eae6ef691396060ee0159f81bec37e72513fadba49f756405fbca86d4237982e45329b4e08f0220a335a666275515083d156c151f71508e710062d6665b07bea0552f01d8dda71f4afad214805e6aaf09b9f0af88c6f538251213b5d096d78fac42227d7840b42e7c8e605585ab66bab24a58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h527c68c1833d74e810e98ed36d234dc4cf7f81f3223ef4b6569f508b212ef340068372a86e8749d34d0c159ecbfac3063b9b245179668e30b2690e7743fad940a25d80a1d1a1bc02d7dcdab5dd140fb925f6097b12c46687e8b824cab15f105d578a00fbeaa52bc7870b7919ec0a412e1b250f894cceb0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e2051c8a532c31da490e8ad439d385fd82c1fe31d08a0d1a80b5dbc1dedf6aea469f5418dd83f22caa96fe6bb2b43d6300670704a80e54fc5ce0bbbec9eacd57a97b23ec526bdf3b666601f55281bfd4bee7cdf862ec3b455ef0bbe9b5d5165ccabd561e237a2baccf4af57d85927e9f960502ac632e1e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131104ef3792a4bf8ceb5b216b2b0d62e0ed21b67aabf916441330476cfb0c5d856893d04fe980a3adffa1b3a057819a4cc8a4c44754524ad2f457b4e7093da2b9e1e6aa2de30cfe37ff498eb5c99ad0e1fcce2b2e51a365fbda768b9e0253684abc9fd69d586de9f9924de3ba84ec51d9ba95f48ec8bf861;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddac74adfe45e0b4ed60724fa62c177b231c495f10bc1df361d7ad71a232832b41ac366e1183cf239976d0eeb50afe1d64993d9daf3c5c9320272b4ff2aa84c3853bd0f3077cdeff553272b3f2293b941c80fade71bbecaddf34c1dd1292cd1b3de617bc0847dc673fe7ce0e0565fb7a71d6ea0a603a8c1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166a90b6d87cc02b3b5aced4122cf020af89de3abdfc2d856f497343ce0bb2356442131bb4c3f175f81feb58ccb55a07f3fad1852462734cdbf18bd62160288752b3836e2b5c9f2519b1987c583737ca4029cd3cc7f726a4b4ebce24b65b5467109c3c3b665410e83028c6edd24585fdcc34cbe2a40cd37c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3a7a8ac72115aed72df80d5eed703d58ea6cfe7b8502412b18398ad179b5aa662bea053f546cac40ba9ddce9b0532ec588eee715c2883e89334a23090faeab54c507084f92607815456fceafcdfd717c3fd364e8574855a7dc6628cae0b7b13051e61a7afb64001d032f6f3b530cd9777427dd1c2c5a47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27779dd8b7ac982f50b086e8cdfdda8e4c698361e1ae720e4d88d8de8ab15de5823c4dd0c15ff106abde2f0709027f14a724d9759a16f0b9484eb79bf77aa70c3e979802c24b991afd27b1aa8b7b7cf40fcec749b4796647ff8b0e74f00192a2fdce17104ebbe9b4ade187c6adc4ccfaa75f20b89843607e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1366a43e13fbd65df24c9a0fb77b12e1404d36d32a5e644d21a9f9acf1ce0504864cbcb2fa524a0b063af44c4c7dca4ebfc1f9f3b5e21f278e7d0c6fcbfe9fa9ead64d6181707032b61abb0d13e481ddddd22e893a9a0507bf207df6d0f34bc913e763da364548af1eeb7614ce2fcbf20c9fa36d359aa969d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56c7a9b1185a9f6462aa8741e1927a1938f4ba0de70e7a72a334bf43d9ec2fb9483e5b4b9fb1b24906fab951b7982382416d62cfb70bd03075a11637cddbdc131e6eaa64f57701ef10ba3f857d13f4c1169059ea1a7bef43e5260a45e7e4c5bcb6b73f30f392c5f63ebcc3f9aea64ef213878c8ffb98e26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bb06b10f236e610e196f28eeb27cb73c6f3b05e578ae63cb9e13edb1a8efaac666c1952afb372501af21c6b80a6b560c65a4bb845bc426f2970981a66b3656cdd40877780f8589687c613f5ea36d56e04b655eff161f5c91847d887a65beb80072776f562562d22aeaf37bc883c6392ecca9189b4858250;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca07eb42ff8e46b07e4c79cf0707bd41bf61a612065c9d19ec9b74d7f211c7ccbfefba23db71631069e6f02ac7820922c59992c640a352a79aed257fc5097154ff14296af1de9616e09cc7bef28772a69ebeb71b2e3fa3ca0009a4519d41388a637e643d1a6fd706fbd0ee8ff0ad730484a05cf7cb33a7b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he801ee777b7455da6f59b4ff000cd81efd9b834abbf770bb826917d55046a72ac5e817d256ffaf851df9be37d95668803e1444f3336b8403cd0d31c479729642896c48605f1ea701cd345ea95de8f5ede6d4194e7e8bb80411cd34749d171bd7d982fcd2b1e0f6ccda707d3256d75381fcbe55c629b9b5bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc403d8375d5589c0ba04a9f499beaf6d004656b9b6e2818d08e8fee42f6f083f38ef14559d82b2a08821b68238ce42dedfd43e5fc69dba1da2b59ff91ea23c3cbed137796632ecc2cbb5bccb303c476311762cb9f613170485527a1c7c70bf8aa4fba2628cf9a6d7383486063ebe95c51222d9ee422f169;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178c5025e4dea1f45bfce673e46c12ee7558fa19a1d7c6cf9f2746d2c012aa0926640bd7d99d85041d0a62edccffd772882433b19edbd93e72dddec2b7b9eff15bc5583e97b0505dddaa23702f937f36e621a566d5c4a12d335e2becb80daa137b4cfc3251f3290d3f001c2d0ad76eab3ccf5e904c33f4018;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf099d22060bb4d4b577948b68f598476d8fe79e625e9731acbaa3b8923bf0f517f2c756e170b8007b1fc69dd1364d62a70edc41d0c8feb292765e0b93167f72b23ea264ed321df5f6575e3f90ef7dc45fd1c695a1628a60df48a4c0e9a37f521fcd3b5b359d74bee346ed5bd33724d1a0c8c12027ad0ca04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4a1a747b260e993f18e76d2702dbbf469aaa855f61bd38a9de7ec035784fbc1d4dffb079f1a8af4f759005a35c5405ef664e42b7a83513ef383b543bcb57b3ca93c914c3f622bc3ab07a90b3eaebf3664d63b4f7fd72bc68c8ccf80c3abf6a71386d972f2738d292c65f03318be9308ecc2da8d3a819dd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h578d4b0a27efa2faa5b56fe2473ed890b14df8f4fcbf95baf892ceea3f2c5dcd12d1d4eef51c945aa59b4c99748f45faa599495e1af22968ec48e68bd0cf15d34536b7999e9badedf027ce998bffd3c21763d4a8f859f743b1a095d437e0caa3b44bf597439dea34b3c0c8b5765a53a3628ed1292ce951f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44b9d99808bc9fd3afbb9637dd30d762eb74607ba15271a143fbf1fe6086394421b7b8af407f26f790187dca4e189bb060f745fafcac1b76c43c569eceef142bb6a718b8ce8b2cb9c5d197242dae09933a2e2ce9181bfc126ad01acb0ff2f65c81ab78bc35bc410556f4b191440e117692849a7c823fc7db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95b47c3347a4ee6d8dcd3beb4ee680a70928e47e69184d71ac3b90ec0ffd741b3ca89d491dcc76c12d9341ce5258965f7c98dd8aa38e70aa69ab956aa718470d295018a30877a3e49575aeeab785996d767bcf8f0c0923dfb6ff97eb54acc15e30d13b67b9e82767ff81764e2ac409578e83eaeab888883;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1130048a3b6958d22fd2f72234195dd92df4f8360cb297503a88bb5d4f00ee0fead60ca957894128b7c81c2d00805068e46c479f0dabf2daea3bb4f247147286b236e7384b6a433d506adc65a9cb7dc936f221cf253b082d1a3c2853032466475c2ceed8693273ce4c8e4e5019e3a3588a2f32113799fc16b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15eae26baff938a3671f47a746dbb4f786020946e263a0374f900c88ed8dabea955cd3238be6caf0d977e98aec6c0efaf3865471d6d3a92d622c7f430229bd01310caa66fae586bbdc5b7024da03eaf04a784fc5c2464713e6f1d305fcf8b76b9846468a356d55823ee121ea54f36ee6e6a0053b874bba33f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10901a5cc076de8c11815e14c1fc80d5ef59122183b8c979f2436e7fac601ba3bf1e2b6c98ded4d1a5b8e94067e5c1561980183f4a419de31d369d4351473a7b37f743d326053a87207205a77b8d8fac2af4a0fd9210f69b04811c42243357cc706ae8ce26a2ff2c7b57e5bb1f2db723fbcda9521a3a6a058;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85c5fefb11182cc39cabd449ea592b9357a6fff22af6e665c2285534ed0fdf1dbb245b9cd078e933cd4c16d7139ff858ac76f1b6e24176390b55310dcb71d89ae7fb2b39169f825e989e4c4edc69c2d90a8b91534ae65ccd378108047b0ff967feb383b0cf657dcb9e73e4859a6291b191c06c7d28b6f286;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4c5faa17220a31b5672b574160186709ddf8f2cc6f6d25f37d163dfe894943eea3a83f5f5d33d3ea8c6a693705a3a519fedfe05c1f60f4b191551fcf5e22c33613ddcd75cc9f6cf6f0f1f15bee6b18fa6a17235a7407a3239d53ff37c9ddc28d5f95eed62133922667c47075467a8c128229af65d407282;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da30b8abc35bb9a4f053059f30eeca56af084bc701a198971fd24db0fa996a24001911799c735b6e229c3f135dc8be55a20f5b12f9a6f86ffeda06bb50b6015c5c4c9e41cb7c0d4cd9cd16b9cad74af81170bf93867a04d4ea8c653cd8125ead68a672dcc6a7f1ea2f46750bdc3fd28ac329a921a414ff52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113e8d4da8ad7eef51da86dd96ffe14b3a6c9337078748cd5e160e86c1c39d34ec4a86c2f69822c9703264af6572666050ee1ce773b74df562efd20d178735e83dbf15fa1b070448bb2352820e8fa003691b15a8b84e678cb271bc22600219c7e7c34223724492429a66c5c93cb7c33be5c36bc4c4679289c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3c23148185f72adc1914f843de4cd97f0aaf3366c43207979852e90e2f8af2fd028b41c0bb8b4d434d521db0d225f8f72042b943981974236700003f10561d45caa19c94b529615e87390e776803576a9577f2863664d1fc46f7a05d9228cc83fdadb946df4e0754b22f3cb26727b05766051b8a46a3ac2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbd6bca6f88b26013427cd1719ab3e2309514ff06c2d5dc1106bb09c663b9cd6c5ab60a887b56b62ce48126bac2020c8cf81c1486e2160e426765de0b2e3dc32a46b826a4856054ad012fad53a1970c7a8cc17a4c5908f8c226653180029860a2de7dff90084a0872d43e1321a4db0b65548ca26972debfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156c32690cfdbed53451a2aa293cd1446f62869ebcf13fd0d9fb21efc30c065d72c5935d4e781a3acd9289bce105016712bf8b8d312d6f262814b78c579e53c5120c15b79a61239ab3207db3e9080a032f608c57ee5db8181256b5d65befd30c286ce99bc7fb78500828b22aaa136022b0374eafc1f70de01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4d5f1d4e2bdc7fd1069582aaa8c64a06d8bfbe448317dab9635fd9ddd6caad8fe170e26955d6e9f086bf3493e307bdacffe0fa37c0e2f427c465b20a06b0ee170c852388e32272dc09608bf1f942e8f8f407a5c2f5ca0392611b2bb95654ab8870e298eae4a45cd985478d9c7e02e33320693dd9ec38b99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b4b4e7fdbb69ca5bf78218fe6b3729b55b2ce108636db397e14d9e9c7dd49f1d0a7f315725d3f3fe51dffdd8f03635727d95011c75d141d35063e30535713a1abb861dc1d3bda283e0197c384682133d50b871f8d517c03f07a7b9e29a25c5a496e3e82ac5ec76a77314c60ed542a79c7287d49f8ea5c06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cf117db6c0938c281c8214278f43b08c92f87b0f57b24b9cc079f968044e199027d223e8f8a4073199fe77c0ad3bbf10f2241041f129705ddb3eaf8946c6f5f30599ce750304ad14a8073be38035352c9451f75cad8c596c3c44d484247cd583fe8d642da0d2604e001ed3abe7ae66d9aaa3bd9730af50a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8fc9f86f43f149a2ee26899bae23335c7cb218670e5903bf7126b6f4d2bfe516182ba8184a527df0ce47e4e00405848f2c7112d6d6364d01a7795c80ed0053615584465250e1a5b748898ca992fa414bbcf283d07bbf1a660a82281069985a1f76d6ff0038fdc7a19de412d03bcaf8230cbee5d73320c9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha86b74c2fbdcc05bc2153524f95891b910ec01857cdddaa92aa321698fa4d0f9990e815fe3b5f405094b7b12a0ad7dc54c5c9c7bccbd38a0556215c02119b789142cadcb323734d812e85b7c547b48fb8d9fc5fc24494523f75372df68522b6ebef3553f40e92a0960a26b1623c10cd26ee4b4aa2c044115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0201750ff3e2e955bb3d82ef3bb9332937cf00105579c821f389e6314acab8fc08e8eb64781745cf21921cf28c7b88a90b1870f682101d0fca58c4c3193ed6d13c22a34d495b1b1aecc5d0aa38c646472e8464bf2c06a99168a7c718c0225de2f7226adbd471798ac6947e4e94f44192f7f26e9a426cb07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h885f0797323da310cae32f99068dfa13f7987472a6a16aa11de811d4c280590603756fdff7a7143578f249aabaec9dfcc68a35cacbb97c11a4d3fc76b77038f871e17ac9b99256f77a99a7aa34dafd6a1ce559e5d358d19a15a693939483f53ebab07a75692ed23dafbd501b677b1acef4e2bcc0dbd7cc8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5d029b0c10957d68fa7931c91d985f6dbad65ff64c186b59bfce5297929876bc9a89055a297a00f38ea34dc1f62505622e38bd8a75faef42d1416dce958d14d7ddfab0850f132df5012e1bd18e5cb657d59606d8c60d54ee31bc715c4d8b5931597737061eb95dd4b72eeecd530fd1cedb3bd9522990b6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e38e08c6f5576f4062055f6cdae79493832f1d7ad87236196767fe7cb5e788fa62f22e677df8c19e9eea74d07946f157473a7a900f847ba0c29e2241e2c978b512fc94d60b1fe5cc31742465ff47b994a87047b312f09b7df2c1be154b905cc8c3fac12de1445d92a97ccf95bfa00e181fa2e49743dde960;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e51f0fc1a86ea33d62f00657e9a96bbbaed3cd8754d1d87e269906244ad8eb776e42451ded2c99963920d2af0dbf943acc9334a478bc2070318145edfd99a00c04e5f5b106cb0a9a87fe033f7c4c9bc275a152816eef71e91417da6b74ee8864f87b4b5beeeed0dd54596f30ca1f3d579b7147970e110298;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ff64faa7c7fa8d2777632efee02483e6e2fc0c8f19bf953fefa59a21b43f22af1d4aad244a2ea5a1deda48eecf7d029f8e0f2362abdfd342b09540b9493d59fb9aacce2ec6fa084788066e6a2a8628b1b75e7e8528f873493c1045d992f2c4cf1b7168fb23a0e2c461471d9b97374d1b71bad3863276d08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa7ccc22f59b8f1faf77f8e70664fc8c02a9a0b031b649e8a8c9679918a4324ed566656b347a35717c8f827d8fe8651d09a2f6489ccd1fc65e6603f6f5994c20585ec2730697f0d23ccb86e968045a0ced5e35a9e415ee0d06aed0e9ea9be7f9706d788851aa71969ccc7c8381f1fe0e97b4e4b30b83516b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f2bb9f0322f970eea8d3d93b69bd3287d89bf12037c0dcd5bcb172226011ad83c38eac2dbf5c15b53d1d0c4006f53d0e6bd0bac6745eeee693a4f3b047d1deb026fa786011ab8acb97931c9819fbe637083dc2e5ce1a06bd4a88349f85c829849446d76f35f1213df03132a9fdb5cba041cf49c1f9e5155;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4102bd82c6fcb5f4f2c377f1f0d1db46d5e7563870b9fa1b87721d204950656bfc2841f2b9a57afe30dffc4cfb8a89390d9178a7c52b5f2d2c3b8886b8b287a4d39aa308b76080d8dcaee8c406db667bed628e5fbac4de608765596aa927efbbaeed6015d3e57497aed5c008aa5aec0f3fe72d3930825d56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fac1d3512f53fcb3eba515325779d54d687bd201c9cd8b481eb6cdfcfe69c6eedce717c1d24a4877f42ced0e72d839c9921bdac3cd11a63c9046cab24249177e48ea01de37fda52ef1db68daead50a079d7761b5335b95eb4d1ab913e489a13686a873c2478b7534783770bacf52a1b73025ae8bc4353d12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bcbf4bb2550c35f1bc9dbb4739c86253d3e6ba5d8e48f019daa3a56a79289921a04ac1116518d6b6a1ba420662c883d5ca3816f796a1ded066a7fcfae3d3d61435f6f6e175b94d4600017be9418471a7a3bbc20cab64f314c343376b3d4f3ebf3235100a56f90bff42d1c4eb8bc6f7cab003640d5cb2011;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b5dcec3125da01f3181b710394e987ac8e45c28bb9c9bfcfcaaf83817dc1a453505db80f5fb60d4704790beed6ca5b510f7a62754956e319c90fe17e51124d9acbde31121316feb3f9cc29b21312f34701fb8f30a0a129795769e3fb794473ccb9ca724c8645703be4e60d68002559a0996e3fd62feba35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125c9be82354372a70018fb79cdab185444ab1321cd2adc5d7ac391ac2b772d2f8f9ba2754368479fa4a562569510aadc796ddf59725010a22e568514706eeb45cbf934adc1fbdd30139d05da856a4a828e7a8c2768dbfcf713ca0faa58c42f687be05cebfeba83d35ad42026fb973a237aeb4a17d3fb90fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c74f0d3c24795f361f8adf3eeeb7a157e010e58ae6d76d6aa8f01e0fb8175d67b84eae8f07a6793072032ff40cc1b4e538987a9192911578a3576e44cc77dc697ae329de78018bf73ea90751c1a5948a6b45f94b890ba1beb3151778e68447ccee6508df2a32ad8d85b62c35aef577ff6f4c297881d54f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1230117b594c0c4bd2245357d6b3044097cbdb7abc8a4c80ec379abdadee68dd396595b12ba7b19e72e9afd2c8d90863fae881fdf88eb4382ea24523ce85286753d70c82849f696af4b999c66a7bf6d273f07a61b1d48c60d84a75b86beea86615e4ae6a1c997839fd417ea0ae6f8feb15348ff5a67d51cb0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab783dda077e76aed58f98619158d464f2a8c8ba26b6dde556c28af1110640f0de52ee04e02987c5578472f59f06a86c705599983a75479fb270773ec067e032bf2a1b8c015dc6b00f5628264ffafe23fc027ed226752f9ef8d7e5610ada99fecec800c98083285ae9c846c7d98b550d625a4656d9691660;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a09b4cdccff0729120b7dd82603ac2a7bd424b753c97c205ecb4374d0c64ca1b70081d321ecaf78c1607afc4e29591c3fc3bf91b02743a3179c604c01571ff5d9d149fe20fff90d87de2e71fcb41896edd8ab80d040d7294847890e5b8eb6121f1213adb6340ae094a34ba5af56d9c47fb0f4a6f557554e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173eeafb288ad0508fe8422a317eef941f29f41ed07c098dedeefe02269dc5fec56dbc0f18bfbb814d9202bfb1235fd429ae1622a6ed34adb053668c9107d76b981a9883c716e8d0328f167726b95c9375b2f7519fa4f912d1617499198c647458cc7aeb2186c7ba4a9c1b2f5cd6c245ec8c8729cd44bfdd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3b997831c3a82f4fc0af7e1ee66bdde5c9e3d7616607c23967643124846820da69953d3446f45d8bcc171322a0816fe55f85933fadbae0bb49ddafb56fedda11f9a25587f6c32338ff11abf1e6f9d390f80cb96590e825d82fd24e5d361e6667e2e031f1ef2cda1120a025a7525db8724628374b9a425c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9975b6307ed02dbc9bc0886a622faac73feeb0515d85fe9f322f1763c7615e1f631b921bd8effc98f34722cbbaf8018b7ee90dedc2552fc35b04368538e2a11ac48c5554672dc40444c6fa8e886dcb8a31414e297f227a82c55d53e16d9d52082495e74db97ead0dedc6bf3efa164c9da3ce2afb8937b10a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1322a7f6534c5a4cd9466435ecbb1a38e202f4ecd365d018631d67e7204653fb347b4ffdcdf272285b447d70d8b820674e57981416c840f3d4a0ea88788c540ff28030453dd45699e88afa1461a8e2dbb1494ffa8b784d773d02be131f326415c77d6dc0868ed868e416b521e56dfc872702e57f255d4d46e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6d202a7dc03e7ceab97adc5aad3a6f03392066a13d51945c69f7b82596c838cbf4bb8ea0e2723ed10c9de345fab968228374ac2b5b999c9bcc1f55a0821b6bc7e529f0a5af0081ad322c297bef1e9196e0e6b12d8137c295339c30ea9cfcd8d17821f897a13bccedfb8ef480b795e8304bc808ef03acd7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178bc7e7db2dd0ac48db577633a16c93dd61a11b983692334c6c640585fb07067d42da85771a2e010fbe0c478006a708721ef23d100df92df0d15d38e581301e43ed8a33d97371f56c0342b6d089a335029f4dd459630dbfef14a36b6718381ce92a680b089e70144cae1a31868b7c99fb7636152135cd411;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2ad705d845865b05bbe2751332e23cfdbceb23ffff491194000a9ef5e25919d79f732aa1e877416acd9e8e6ffa62e0d4af5506bac44b6a9bced44132d709dfbf57840050cd07e3b60334aab6a68fcba40997314d4fb4a0aad5cd2cd6906e2532f6854108faad3d4e619dae25f168780ad91a59bfe8e7a68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd584218ea13d3b0f3c4c5a2c8fc0a60ce03a5d4ed786f5c320c7be89cc53569c7bc79eee46dd04e5d8378da420475923d6d732a562b60335a7402e6a318456358525de7ef1b73eddac9ccb9736e8aad426fe5e28b3f9b8368cb3c8c37394686391c03040c4ee8c72dc7030f07407dc923b19f4df254bae9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146c2e6fad490653c7e0bb5d623429e42ba497befbbc4c836a5be7dde76589b263439adafffd761a5bcf3de2a6425a49bb07e0242ca86f8ddf5d05baefda99b4849efc49abf6ce982a84c578360bf8898c4921fa962c98d160532503a0151640eb882fac6afb5e2185007fa379338e2dd42f89c73602d6092;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186325c5afebcd2ab3860d54122b0a0ee94535b55360e5e2589ef1dfbb8c6c2ff9124be017e268643f0925b8bc4ece9f7441c0969c6e06378bc1f2ff83a87a2d0c5d75979659b9bbaf878797a3028d4736a276ee5b00322c7b11f8d8a3c0c4999924d2269379311b6aef124816a7a124a464e1b8f1d70d79c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fcd1355eda453db7f78360f25a7e733142edc71b3e63395f3dc4445e217a9b5fcba45ee3c3f7909719e364ba881e979f24528b61f2c468f7e007393d7cd6d2debf96d9db9f1279e26bd83d25917ed3f68e03004ca2b994187ccdaea63cb4a032d297906aafb5e1ef006d76147bd2fd4662f64214ea64953;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c8f010a2d493e61c757253b83cf7054c7103ded5eb1c636113a1f33a400e74ba1af5994e5dcbfb72c4eadbbdeaee138209cf5fba3a66d4c91bda0c7beed85ed44e0be686b8839166634188d36a0e54f27c5b5e8fc01024bc9c16cbb649420034d829253d83e7c29f7ab6a7eb365dae92ecde7b48da2cb03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc90ffe58eefb4d921d520d3b74068dd9b138ba5e0684c96c55ffcb4f2bb100d0c0063ade6b3a03a1d1fad28818f30f95422e88c0f496ecb5b466b24c93f116423c583a38ec3e2237cf955d879039cd16dc7f80d82132bd7ec4a32e4acfdc1e24e281167451a44ab960107bd16e1c9c73c94727d953bc8904;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde5022d86a3de32bf15254272bb5bfe3760e853b7cc4333a048f06c7f8a913779be4a7eaee4021c66c587f2d36d758d51b97c6a716a3aaa43656b0d27da63a131d8b38c7ca5296b2ec247e9afed5ac91ca60956bc72e61574b827887cbf2ea3213b15d4cfd64971d83b9248ee6a3a2f1c360711046241211;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179a77ec91948e7891fc4a2d5c0888a7cccbc93db08b11cc4d41a871f8e73e860ada99e934a5afc3fa4d0b2e243de8eac38a9846615e2460897f35a6cc2cb65341d188ded2030107dcfa1c825d9d0a0d7975cf529bdd568dea5700438d27a9c20032f958569a3b064e3fb06727be864f44ab483dc5a7267e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc365f12ccad13c304869faeb91c39c461a1737432e167218baf06b34b0b536eabc5ffbd327919e1a0c01340c061d5cff8019f71d8cb4fa009f55ddd25f457a14e3b266e14d52fcc5cdc930daf3f47282af6439c9e31bc1ee44604b04c272de0806b2974cdb997aea95167df4869e265d58f3e73bfd503923;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15373ae50ca1d81af81d8d58c2cee580695c10b35a17093f0e196cc3ce7c90e3be2df5a6d6ea7d758f94e2f99329946b124c0984af388d89adc73e47d7cfaf5c8db89f890428dafba7de819194391e4ddf19f7417effcfb1815ff0aa9d80a4d316132677e17ca2169721130497c1b89e1fba856f0857dd029;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha96e4d2b28724a6d34da78b2843bf4423b0a3937371f5c01359ed36f621fdbab2b787213fdfffeed51f5321fcab343fae358bf6943a5c16e246810817632bf0c393eb331fa7bc26c541fdc99e5e2f6db6c7f0bc0288c690ea60a0585fe7ece539e8c5da853d60fdd2354afa9334bb9340b90b442c9a1b8a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfd2790f6931ef3221ebc46e2b77cddd65c0bac33e96ceaad92de2c6b068d32c7be780d39effd9763d3a3fd1fa3b9981d27b927c32eba1d6b2a770e1d0437bc913d077fabe844ce803edaa576542a63c1335250913b8e2f49c12aa2c51a79e9f67e7312727c3fe22cd0e40ee6ea02751948c81f89b88ffc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa473a17c3c5a4d3c320e1c15cba033932c791b2cdcd9c93fef8384375a028c585eca8400d996f1658f877430cc272d4281c6aa6e1ca1acf539147d70bb7e1bb06b6d2a59b348b35e6d0df7e9bf660b8163bdfbf225647439a7492cb28c789b156f7d9120294adbdef0f8cef0a9cb84ce90ddf8ebd30e990;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d67bc1a4b1467f9daa2d62c4798f5204daad2ceb35547a401bf40bd6ac1279830d5ddbc8d655f97baf99c261ad9c331be204a81ddf772f350d9d2cff04eb083b86dd33f01f387e0f07f3d164cf77d3eb4d32f306454c32bd8aeff31023afd646532e06c8707b10d94b3bd2a969b5d77404806bdf55cc7567;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb9f19ebf1af7890cc131d84f56b4d47b80c326889cbbee42305fa586737012cca23c4e19119f7b246b436cc31cd2fe69931476192e02580308edc6a829b821737e990eb524360f3a1254f2917cea177b486fc90779d31d6dc35988385463f5fecfe40da1e605cb24d163296db5a08e27af9df64b98be45a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82d95b2fa3fbb301fa14ff6294ba9c04c2e864dbfbf61ff381968663a945bfa72779e7f690970f6fd476dfc139bd5c18947ed92dfb55b2763c0b89660b29de84fcaada2e2b643e394a3e134f1132bad9a4a443d9b277b8b64ae75cccc44cc8bd05e517c1178edaa7ec0596a4429521ffdf7c0d055e85de10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c493e8136cc6ec5230e25993d934c3d214a2d7ede9cbf09b7a9e5b513da37c894cf311ff9f6174ab1009eabfb2781dfda6e2f4a180d0dd2668fc9563e402eba08d073c53c3b9e9b84f95cb90150e942f67c4010278fcac418ecd10c8b7ad3679ab23d20cfdb949fb37cb070adc3cba3d4a0ccc199a62e1c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4460bd517b12af43b842c7c810265e3fef465d85b426c153037b3c500430870cdcc871d1c6c477cd259e2c918a7364c306f4c44165c9ddf21232df97b2461b9dc4b1a9dea51fa5276d02a674018d40d9a5b9515077aa159c37a7a9ddf4315ca86856c1e68ed32ec11d522b460fbce6329dad41329ec0c8b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a524ae746112cf1ae375bb0f856e190a18ed20472c14d4fe78de11c811feb7b270a5251e44a58662de677354c198bf520bf06c2f458bd8cc5f06a8eba782e9394b447c4d646c5fc6e98d3738d91132cd42f599d830b8ae387dc62c2ea5c40493d583ddf70780e22987305f25e7be4f1230da881b68c14fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a959ed15243eda3f7df34e0a85f3c0359bfab280c13163117eaf5cc86c9e56be3ee8780bce355a54a1a85c340a2c93b9852e6c36f83ad3cfafe52d64fc34c7af5c9313c5e00ae195aacbfbc08561e948feeace3ed63bbaf4c29de9a76c6d7db14620f1ce479c186dbea5d8e543b080a8e90c5900350ba39;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ad927fbb05781cb9243c07ecb11d33402ee0933e735ccae365dfee86bc7c9bbf8cd3f00315ca4778011376ff0a1af61caa51bb4a96b727db846cdd8bda4e02b8a853af12d835db6a899a980dede11d9b9ec8a827a8fa2644d7baa3bbfa191130e5506408b65e9a6461530331bee7b9d5214655c0203c9cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85f4d02b8ab049492d0af03c110147f2f6eaa2da08b17dec07415031cc9ae0e698b6a723890437476154babe89ff513e9f976ec925da13acda9fc99bf750d7afa5e321ac40938ab6bd99a60b3867ed3e0547b1fa61885d70730d2663af7dcc97eff3f51db8292052b99b46c4a06af7455eb146f1a4a22dbc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18133709acde74e99175ee726f01b22c252dbb074ddd5f9817f8e6ea809b25b3b5566fdd9126261a58a8f4ad75cd9a9ea70436f523c3c7e7af5d384f9d5acd315ad7882723051d995d255f71e24d9c978027ac29d268806b8287ea0762d35f240162e8ebe0bf02a4f7c05c2cb4ec05c1b912bc2d846c62e6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a3bc4012c0a1a46ddea1b01b47ebdbe7ec59c71d03312816670a1b954f4e0bb71a07e0c1313ee9ab43185f252e6dd97fdf01d16d4f6006bc215e69141b35992719215568035315604db9f16a3877706ae70b5eefa8ea03f6adedf58dbd3859eab7d05d685cddeda5426c34cfc24d44fde9fd0aa81ecc7e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e39f1b9dbddb7cef5089011244103b487b9755ce62a09dc9d932f58eaa0f9599795e7f19c1773f2c60c5bebec235dfd2e0b98097b4d93aa5edf30126f5575032994a490499a66789bd7b5f99560a3249f7ce46c27566231623c0acca0dda3a0eff72b99b02c57f980067ca6fc7cfde601aad861404361fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cfdb0b4d8e3146ec69485bdb889d0696dc733d608f98af738faddc0142bd30b415c4580880891027569b8eef782b70d3d25ad8aa6cf6b0f2265a39796ff8e28885a01bcf2f6ede40acdd2db9fd48b07f4083a66136151919081a6446f2907344550171cb545e86fd6de39cdd2ffe760949d0fe105f79071;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19933165f17ea51a8e654b5adb46c6f65e9a12f3f8d38ca76b81f5945a7f050882abf990af9517a4b79ba0cfe3555551a0cc45b7385237b5034cdf0c0b31c89c761f682db7bf3e0811bcc3cd51c29adfe55727526554123d6b6eedc990c6bc84cb028b87817f3d5f0743d762258d5a34d2a6c56b56ec1764b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47ef8e815adeca35eb93170ce5128f3587ade72c73932ac6998ae114c1feda1068564d2d9e43d365eac379eedfe9859cdc4258182632790cc391a93e00292e09d2971d9ab3fa978d4230458d01dd881836a3e957260a2e8550df2ebe7f25043c13bd9621753212f68047aa09f36565875c1ccf0b02e5eb48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7d37d73369217750758c07db6cc71a1b606586b1a7f3676186a4ff0aa00e4ae05772ab016de021298073d00e12559924fa07e2ac573dc811c258eac85fdf6c54b9cdcc3908308fa929e721f48b768fd51e7ab5ad5b712f830b28394693b2b693040948bd00fa59acee135770c75a206335b9942c7d00e76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1925187dde7f58b2a7e63137bcc78748152fdd08d0c8b0cdf1eed73c94467a1a052106ba9199f7c241a70e6d1558cf26ad1cdfb90a26128740a7f53b8918bc184d223a6af8086c4347fa18ab2e41607ff3c6dd29f868915b3c54768062c3eef8dc16568ec32d467f8c89b9f28f074bce1431ebe0694f676c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144de13f6099f1131d6219915c795b368bb5a32cdc34f8a0111984d588afc6b8b102e4f1130d15ebe205e4dd52c6943853f31354a496062680b80f5b05264a8a52ef9c935134dc8034dca418490e2c78788035cb9ab74bb0e5873b1c4eb0fda9dfd93e772cb608f8208275a2896be68cf7527e3ec8569c7b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bca06de72623e213a907b145c5f700b0305c0cf35bae8ff2378e94901b68067d9d74d9a9f979b8996ac7f6338b0901ccf14fa69a0d7906162b9f03231e5ecd707021a5d51c0e610f9eb7a63de176dd7de35f5da44c5e1bff07b85120b72d47af6bde76d579d091149488bbf33a25e4a05ba5577e9c09948;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a49a47797069ad161dcc31823883f0114d579d77ca2efe8dd94a99a96b3586849951c8f7a0c2daa5a7e9052ad2ea27e1f45ce088bf565c463706f16c040aadfdb751e22524fe8c650f975f5dc0e4f45a82e48164e1436a34a4d87ed1e3b0d15599e81d5b7b380788e7959c6b308c0d5f9fcaa380f7895792;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35989bcb32fc240a4ef67355fedd556ad7b289ab29ec812db419cce29886492ff3bfa9a171032dbfadba9aa71fbe660191ef870f55d9ecee2f7625f8b69e6442dabdb039bdabb4474c0de17a0e0b467fc6cd0a38145d67e16c4e4027611a00e5749cbe955a62ef4a70b193890ae1e2d15a363531144297fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc6d66d02bc54a3a0584d1550f872c25ea4afb8758fd5eca76af65e1287d7738bd3bddcca22965ec3ee3c1d05d124afbfb823ea55de261b222f00c127ae55a304a9f3c5e72f9e59280553ddcb558ab8edef8d4ff4b2f469c0a12614444ff965582e2efd19332a8071ef4d750b6e9683e5eebf10e8686a46a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fda8754309ed935a5c8a3c5f812913362ed8c13e0e4fa19fa1d1d499e3decde664877679bec567ff8fa09e4b544d39ab10040b810b8bcac49618e598e1ffd5c62811589341d73d9235e8232620878f61a478ec31e1a5905bf029f750ed6d171711b6933a95620f9900eb90f353a2c2130ad38d6f468353df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf412f3561a37ee68e545128b86d7d58712a64e45bfb799115fd1f3743479fe074919628070f252c92e8ed7b804e4d826ecb3b9327e2c2718e6392d96cef862166e027ed28645c98f32e5435136941820a31e499969f6c45dec779f241a7821988693ff34e88229addbe117a66a404481029ffc94b48d23e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e5124b6c3c45d809f75b630ec46394f9942397aeb38da2471d7f894440eb5a785d1015db28181fb3153635836e3774d80806328d8bee88ca4c737ea117162a09f8ca3a60e6aab51fa8170a3cce1d7953a5982626e8b002e3c955b8fc78d4589b021597d3d29d65277a6c2916af41a11391c59b663d63c3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5220220cf8271b163ee6dfece58264ca85611f40b4b3ff331cbb29f03baa535d1b3e23f6f1648f75d1b7cb27523a6ec9d8a2f4a6bc73453d1c8624c8c8c604c1caacfe30d709a48bc6435ed72c1677797a25b6b3f243d97d7300884691c85b4499e9f609ca41468eafb2eed25d4fa5a3a24b86ed5ddf0945;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d42cb455ae509f38ff6869ef607776773cc9a17905a0381b9de91fe681ebc9a1213fc8cad005cf8d9a9d8020f4c920f8b51f7b7c825e1a68896697c14dc84a9424192995323e98d12c2a3794e9b02e9628f725f73d636193f07f5c90944968c67094b5a97938df52adfae1f3337adc3274823a6683139857;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0532787e912fc621a3279dc25d53531a0009960c3c45389a063317e8cefaa92f08a809bbfab5b8606984b8be9ab1e4c88f214c5bd0452d51bc45edbad9d2c7f0c03455d9212fef815fecbc08de39ec168a3582f3ab26ed72c905b08ee53e210067243af47d8d24129a9f1e775269f506b9f0ca3a4b2baf4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf92d81d4e08590afc69538acd449888c614995a53ad55ff50583f7d3e648ce765d5093bf7c43d5ff7b229cbc358909df9716c9af204e3e48dab7fdf295ed56990b3633f035bf184c4fe38c65a418101cc8f9ac6fd79f48ff0d0b62ad53fc7f8fa9c8ecaf7ff641af8a1cbc4827b7cbe709c3e4c2d2800d93;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h546dde708a599cb23ad4b02a5975319127a4265161cb8fbfd04572a8e97fc5d9c597ea9dfc271a641aeb33a218b3756b5effa83c27f4528e09eb79b27e0424c48da62c750da14249973abd0ccbb4b729af89eac0128705abd46a6a771d6dd33361f767950e35208c2cc92938dcee82faf452d967f2d898f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hade56b1c654101504756fed416444682498ca5e1250a5c2c76c9175ba3fd43955ecb9d7ae67fc94e55ee3154eb6a7fc623aa1f289c3734ac27d315eed6382a363a4ab373be2efe87f44750f51c2d2b315d09945a43e725987ed3a4c0730e0c2a44070a1217fa8f392c6baca086c5051d7f896c27271d0f6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d69df7cf7f3417ba9c0c49db1e072017e265559dfa57dfa0f66699e6f10d57e335789a94f87b93b3894546521aeae75c9c3c59ff93b3e544d51abf0bf3c5b691e477428cad34c4e0b4ded4c35d3e4b52126ab19b8b954899254bb8de8c0278588672384bd76e08bd05b371a953e3ac53a13aeef9123aa1e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e749573a0a78ff402fb24393fe22a8c2352f60b8d3f51f1679fb29ec254099415e6f0d15f785a3e95978b682f9308378e34ada5db160086bbd1f07bdff31975fc6def0a5c061e875030105867c492fd61c1377bc47a10acbaa1a44d319581640e19c4770d020fc179d5d9d80d392b8d77154c423fc4db73f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcdfeb3e4531dd9409758c298af6c6e4cdb9773c10a45ae0f3c1a65b13a02326ba0356011d7605fa3d155675532fe8c6221830cfcf16df51c4cf21f29a0642decabb8b52c57a7368b56f2eb4545eac01a853b57416235a16ce51910952a597367c98174ab86af8ca7e54b849b282e6d3e79204f4c6c4fa783;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb643f3891d24881dc0090317a33f987b52e1ed058ef52873eea5daede70eb3a3c37fdeb60650b9e2468a6f5a19cd65abf7b02f75d7d0bc0d221125af1dee184e66c9735094c63cd415153d912cff427625135fbacbe6dc3a798d7d0ddb47e5ae9f610a1ab2bf1708c6645bff5edc528f0edd27b6ae263ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2bcd41a447fa36e000564e4cb31978cbcd9830ef36ad82d68b1192881a0d1893e7bda4bf13ebfbb45f367cc4a1295a9c60198696431f474da7b2ffa0a459452f4786363a7307cd5376bfb7bb416f55b5a94eecd8c7bb77c7ed022f164a9a27191929109712f08fb694f38db71dc7d8bfcc8ea32e150c383;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b2ce9a8796967067a33615654cb1e322ad688178ada7eddcbba395ac862fcd4792846267b8bd2257861ba5636afa7a68e282db5f5232e82509e413a6c114edde4816f922263925ebe7a49379e3dbbd2e176186d875d930cda9774f2364c6dc1ca383c3f8aa56e913a83c40863e63839553096c339a92be1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cda7f36e2addb9a3e1f67358a6e462e427627f914d8d6a64fde876d13fc0c3aec5577a95b51e089ca2b2c1a056ee1dd02f4c8a4220e17f5b6aada946f6945d05ba8cc73c85431f3b790daf629e78f2bd2f440a4f214e50f0741d696472bbd11acc5600fac2b2c82cafd91d0676f3f8b7099d8ca86045b3d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28d50796cc75619fe03c6599c500c30f0fc3a2b3c9d47676f0c2d01752ddbee8e43b67b2a601e181e63a32f2912066918df266828c03b9bcd0d76f679888d11412af6df8efa05495e8f0135a4014833bf5a1bd5c9b6422f5d08e3a84353bf8a43dd64140806fd41deb26c06b6af6783948c1a4403bd65f44;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31afeaa3d9faf054d1b749aff5fcf809a74e6ebb67b79872b5d060f97edf2fc63a567e8ee2cb2f284e2ce2c6bcc932d2fb25c37e4f1bafc63cb5094ea58c0c5aa92225cb91c27e89560aec1a9025dde0ffbaabaf4b0561bda8089503102d22c3a6c179f1563d371cfc81003692c2d4f2157391ad70cc9a79;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h840a5d999eb8e10e76d8246d710867924bfec40acd8849e693984e11e5fd5e2adc1512442c22cb46cadc7582005c83ae91f1eba4d7819fa7514962b69887db05d8f50e0175130c828dca2d025c472c556e9500711d6d56731ae29e81b25560114326c85a329ac7fb8abd19d6187b566942b4eed124518a21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c89a4b031591a19212634fc823f8a51cfee214d189ee1f16412700a0d9330ab9e86140611f86815046120e70a2930767ad43478177556d7c3e66c11669b505d8ca9abc94adc6cb9113ab730739c87a2122af53f3c3836fcaff09141e47837383b7fd30c7daf7b38aba565358146850616c4392217a42297;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1985b64a8105f2c24c2f10e1acdec3972110da3f7e6b7c4746461eff03360b68acb612acea9363761b3c8a40cf2a99aba484bed213b750c6b2bea51b1d6510c0672c8e652484a50285d15307866697454e267fb88bcf9b3097571c9afab8108d850929fb39d023d1353b06c2354b346df22d757835387268e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118c0c0ad451c82dae914f9ed61b51cf89d6ec525fe462172b15c6367c738502d46226e11573d4edc9d777b3a41eb59b1156f89b85dff21efe20757c1d259c11d125fb23b0cbf1dff1bc2ba92202eb10db4ff3e6e16d9904587917a9a16c826396e93f28f7281bf9afde73a4d2e49811c182728ec1d8d975b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce8ee830ade48eb65c43144b59c1278f1ba711a828561352cf51cffaa8502cee9298775bb905c11c411df5046f4f3e8d244a5016db1fc3373b7e0419a34728c5ce31058dad54ae25cb28be5420b4d830c0edee4671034289f1d0c509f9b0491d8c15fa68294dea228f7aa59bc6247115d8bf599a84848c83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a859e2a43c911ace8879651d436d40a0bd9a02f6fa28e21cd4c5f8be4269bf8ff842110405d2a11c68a71dc4a61ea0a6c913c5b2cfd92c45dd4ab440f2a41a7fa31a1b2b8119a030c8bbd30ce9c1900be4c7f88bf7fcc4be7eb1ddf4b3f0fafc5658a4c6b1346ac302d141932dc89a915cf35c0fadf651bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18275d40c426678e1ce1ffb0a78d9bf47e482648c2f75dcb5d443e94bc96f909db7d81c7c602e5ec9a63939e340320fc730b7ff1be841aecfd20f0465057429bf36f83187b4c8af7493af26a5949c0a1ddc5361cd1b047d98ddeba968d71327d32e2f8df74c67333a0ccfe922c45e3117753e18c59f667b4d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188c3a6d7ae2e436119717eb3256308fddd6ed2ee9635ef707c3635df8360ccecdb32b44c1af3e053e0bac29e0a974726a02801b9348c6c40f92d9ea2dde15eb8cdb8d24aa5a050a96b3e7042e67edc142a9ed8209eb2d6ea74fe871ee135807df314206a2d23f89966021eb07a77fb67382630e8263e55c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdfa7c846cb7512fc46066bc07173117387ff8c22328f60dc5bd6f850da4fea3ee40454b9092b080ebf28e5db0dfcb04b3dceaa0928f8bd996d57429d822e5017d3d2fa706d78a36c2a9da272c4977ddeced70581de2aa4b1ab13224781db1ef5f42ab76cf6f39733ffadaaf8442d74347eb66939cf09f626;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a216c135fec710b87183fab64d817ae744ca1a252edfc4683da65e924bdb229e08a7316e8b0c44ef5c2456042f13e2d592e5e4394d8a7a97b6f479ce55dca32825fbc0606d6b802da26a129f8aede059f4510c42f999ee8d5833734b62cd4ae2bc2b72b226d142cef0c99a4aae0a6a4eb4056dd00d89b26f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fda4ee288faf00fedd3643a332a73172854cc72de6242061e998e34f7a31bae5d396a2c93c67414ab9cc09a2e5df3fad2c20760d06f6986716a20fbaa3c8e16ed54da80af885fc10da965a9c2425a9c73a0eaed0ad682a4a6028ef594e0a9f83c73a9d765669129411eea14e15048208b254c886d8d086c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17be51288b3389eaef615e00a352d3e490b9e518b3258b10cb0add29452c70aaa9444ded6c578d20cc2169f0346c2fa4c517c5afab90c5ae45bcb39fe647e1e0d29fe47ea3b3c2d3c3fe448b104834c03e16dcf985ea8f8ce642b5c5083516b71f2ca3643b193574237e10fc274debc74aca011f6d8ad3d74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1593d5c3676fbe5801343b9f3bf645277ddeca1c207bbcb32938ba4119eee2932e07a87abc812c2294a49f872e3797bb1448ff8f5dfd2885757a391e904b923b07742f3232f7a66f5837a074e13be457cac2b16343fcf218bdd1528483c9d737a33fe369cabdbffa457df1bef22ccb0f6c6aa5f43a891b834;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8a16888302640d0d1f27401f47c392b7670ede5a86e459a2a3c787f8e206f25f232c8d9078911bb14b72bcf6392e577d8c2fd8de5acf45fa839b0efcee86301b231304bae6cc8a3b4149012d345e692e107fb6743072c3379900884e0bf26178d24bff7777ef4d3395ab437df9ccc384c63308accf05b0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb89abb5555c1800191a34a328a09cd15d4482abe3a163436bb6903f27a952c63fc4bb6b2e5e967e01a5bf5762f4dec11db6171d80a326574bd09abdd4e8d4d08702f2d9ca1e649806890d90c2ceffd4cee72c29521b795ebb21884a3ae1bb1ece5cb0154cf37f4d5b787a9c573daf041d41ea09a4b2f720;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1e910f6f01f6e0da2bd71bb03bc1fd0dc2f7036554ebc84b026a8d547d370bda5e39a1546fe822d842e698061a6c5e4cac818a480ef99c8aa2b9b13299837f1f18af612d13d68e4751f64e91ba528c0267cfcf7b40760151f8bb9eaa8d744089d4f2b06a163955de8cee7c764446b0241797833cdf3bd21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b5be440fbad532d94e064c4340145348af7994160c04e101ce76b24020b3a813a873b57200824139abf4820121ccb55a1a46727ab02389422eff9295e18a11b2d3f9d50b10a93300e06070588c164975270c03e84c4b8b6a4ba5736ef119429ae85c8a477e96145ce40b05b1314e368f72d909744cfe67a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h693c375ebb855bb1221c18155994f23746368d243a31f8aa81bd159eab8d4f2341ae649697e5dba9fb3d30cf28452685393bc13bc5f0c73af04a87793c44db18ff35afefb9a830da8ec51387958b76a3a2ff3ddf3eaa9c3290970b95306278683957b683ecccb19a83fac7022d51195325e8fbb3685673ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101bf9447576a839eeee9868fcabb5a5ff845aefb7fcba61a81452d6c80cb43838eeadeb6bdcd95d7e1867afe665602faf54b407dace2c25b0fee52eac718dc39e86ce11ee588040afa2425201a121783abb546570db3fb73ed71a613ae3a0973150c8ba8b64f3b6c1062c3d3abde09b1132c0fe39b46cb33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e189e8f91dbc719eea8f0b4b9f6407a8a97139968b0e3a2f7004e80694b8014dcb75e6d8205ad39f03abe5925392175794bcc524351e413c43f550b1e1402747eafab2ac7015ed98ac7ebbb3b747668a99abe155bc46c7a01388caa9822959e8d479ba61a082cad6f84f1784adc02ef8b9929937b5425a45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ee785a3b57097191ddfaa377df4ddedcf5749d77c7c37e13359d6b908fe853850782365f0eb5a6266fdd07f0766499187cfceab5d42ee7df7be24bbb46854b162cd2c865696841fb4e74747b5eb8ec3c4074642dc810cd335488deb8cd0f58755c6293abed6388ec4f793c27c1ad634b79c448ea34d2fef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0db4ea343d64ed6804881fbb39feb06949773aaf6b45ae6000b8b191f8f1a003453b569cd39c613a6d61b87c799755f2aa67ca62e2af6bcb29570695ebdbec939e4bc79a23519cdb107b4383307d3545a1d661656e00115e6eee06bbf27662cce64af76912d7ab2d6b320bc6ee742559433a4ce26e934ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3abdf970189356f1c41873b81f2dac7bfeaa747ff80e267df3dcb374282dd01de4ac227a1b82af42b7ec0a150d01892af4224d67b6326e9d7f1ec63920b7d785875c4670767b879635552feb4620912c4615022af0fa2b1eb9479a8dabe573586ae2342b8dcba88fd384b6a91eecd65bf442dc65b491def;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e7cf99beae088acd61dc1b82c6321b39e72e0db8336e77adaaf8a78a865afd5fac23cdb8bff826b0ecdf549f88f30e8ccc1a919851d5e6f50b515047dd48e06d2eee5d261755fac806c721df7eb99d6d3fe69c7dea36ee55f1706862d3138fe01b65b212d6a2e239e3468869742bde3219dd5d4d3aaba9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1467f76cc82e8841a1d0bb1c38af463444b7b485f42cc4cfcc83f9c48eb1cd592cd4ad136be5857d932cb4dd55da89860ebb682aa26d614bb089ac1c4a22f3868e0550a27ad9d0f3a08619e0fdd5e1d136f11d7402c2c90296afd81a06dfceeebb463cfe94d7041b1fd75e7cc9828d8bef39b764840a506d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h922f2505935dfa9c019df6572f71ff724871bb71bcc5258a5100ad6697e4b8d8e02ac61d6158ef7e3719f07ac9bd8333d8447408a4f71b79632efbfb9aca9132f27d1279efbed47b751a0758cffe92904337ec2b37c808085c2b0095c1acf5fa8f22efc37e4303aa19bf7b032c55bcf053730f57b482f2ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9402de850d9b87438c3969401f2fa206d8bcc28ba39134df186eddcda465ee3c20f22730322cad1e62caad5b8114284e4c9200221cd36fdf81fb2f22c7644bb310425000fa0838314e3bca1eace312803610f2d7c16f31515f7f8c34ea7b45a7eec35b880bd9f3d33563e595d73fc3fc660c13c2ee43e18c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d64216a83bad9a76a1de911b1ac7b9984ef310bac567814ce0fe274496e7f02825b66fb5a1751292cba87e5746bd1601bbc93baf701045e1a110b9695c1c90bdbbb5492853b91da7e598450b3d5513e0c37dcf2e1870b69becbfa21a3b9053fb60caf8022d21751e9fd33b6ec207a4d593789cee62926315;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf65ab14fdc77ed87ba42d4d2fd507262768c23bf504b5479c1728f89d88ec794575aa7de10f9b320c3b26d057b35cde676ff032af2637d3e57b66a808e48ede0cf8c25870e931020d45c11506deb4150d6c2271cab5ade2539d9a93b0104b83cd50e811b5aacb74565992f2c06ff381608823f52340cb9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b3cf26eac659e930f4cec63f1835535767530825e0c0a94d33412b8c9eb75600012edb00eba99bace850c6deaa8b7437f39f0304208d8e14dcb825e14755c873a85aeb93c6be70181b53e5c097c4116cdd3c073b47332f8654f387ad2cd08d2db640b21bdb2597e8e32f7895dadb4b869ba2a6fb0106039;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ff7e8f08a0f8faa0a4481e0d0e3cc90eea2a9fdea158908549b2844e189f1fbc160e229c850e12f53080d61ce111c65591dd708c2dde1e192d80c26be1ca1ad5850754d64353151c7b65f82d1fc826f8d63f7ea751087a895489a694edcb95dbc95e765113174e1b1d684550da19f771d23f3dcf2e9ab40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f32b93dde3065884570059f1d378f1e8929a5c66c532a0327add1ee73e569a565c815c590a3805a85bbe874aecb15511bba5f29237c6cc5325a5608f37a370728d700b54587520cb4476529adaa175301b74df1167dae91db040dfb01175a90b71d0c875e5844e516059cfc1bff8baa90d9a21dd25c3570;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5380830dea2007524f909ce9e51a4246304134e353419bc4b7b8a4fb280973b4444bca61bdaf21722257598aef8a9bae40bf10dab609cf00c87f7056deccc091b3ed898638e16ed05b040404b0704dc07090e9968a5944960fd85fc6857ddd0ae2619e5260d2436812c7767e98573ceb9560ca69acecab24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abaf1d4333395e028e5f394851ea847f77e7666cc7b9811679d5c0236bcb1aa4a07b4a06e3188043399172c89f6243c895b7be37a956b3730689035bda96e33c6b5cd4bacaed3ba48d8e24daaf78c0ff4792291b7f0ed713a97b7aab21e00fc0f490062b8b5b831e1af5799f2c7599d260099d4a8dd90fd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17078d4ba9188832ee9095bf3e46d5682878c618f11af7e8fed74cafbb9198093c31bf332833fdf74aa512f414bbedf3ae348ff3130032f6f692e9156eb70a7c73c2eba42bc4933c00292be7526a9e28c8e7bbf754eb86c066dcb85af8d666c17ca7eed6832b01f67df6441929b5b49d015fb6c795002121d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178610dab422d9709b1bcf6292135473f2b24411a51be9f4f40829770c9cb49fa102d8ddcf595482232bb3641dab404af94bc3800ccb3040845efb4bef0b0af31317862da7429ea0a6227a2b61f5d7c8f23908ffba72fde556b7aa37cca7501121a72fc1733b861f932edf5905ff6505cf704adbc78a0fb40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f61f6bf655fd0133d71c1f65a7d58a3b1bfadb907a891ffb18b8a63978f251ffe0cc32c32021e43c19a3a5d8ba492f47783076d7ac985c1a60f82e12ebcd66ed36ca116848be95e9f79d24c5d562d51a7e5b730666443f07bad4e3caab8a9328e71654b93b23667025d29175f62035d1c3f1b87f6ba0b7fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97dfaf23f43e11deca72bf814987a58b5c5dd51c9212c5c10904fe3e55d90bc805221dcdf70968e9c9b0641f5215736dcba85e635debd592c9604005591af9113bfae1d66eb9f67dc79d9be65ac1a74ba18c14ee7636c08ffc8c22fd70f64424e698660d844b3a8a1235c49f060264ef8dbf01daa9e56644;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf1bc710dc99ef07a070b3eefc9e4854aa84d035e94e641add66ed66ff1ec28451ebe1dd318559c2083e632a022f074264e5444bf9a46510b9a3a757984930deac2478d335792169ce5eeea9abcea12aa04f154d5dc09246e239bf3ec7cdd72dbee286402b2ecc10b654f3726582408edb7644fdbc9f04aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1328cf3b344b629ff6d2c4019cbf79fea9ca1297fc5c0a0cf2adfe545b17031375f2a9a16d28e2a45297a37576ddcc3852d9ee6b7b3971d6181a0373fd5e390d59659b6ac49b79c01d8a3fd7284c07b4c2ea310cf5262f4b727cf42e46bda82e90431c0d5e90f11b3b2b746edac0245b0ab46f3f6e99b0a6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he745a13c4cd1819c60690ad4614fe47476bf86b889cfea3d2afac0a72648f6e34a49231235429205d6066b1430838f5b7436c3df983403e47d9f9020b6f13c08f57bb5a3fcf3df18dbb557671b0519d103c455f8983fc5bdbf15df1531d0d8d19f9f78a07d1ae797d19cb56be1d5b02231c9906a521f8c04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c20ed05623845ee5fa8045d481eb633fbf29c1a23530474a289d7fadd790d963f3d3e0b4695ac935e85a0e836bcc59d7da3238474a691aa378984f89988a270fe4c15796416acf8ed6bbf46252ebdf009a1243087edbcf14636e2b2701dd156f4213b6fa76f70e6c6b5a574af08994b8c2cb5d3c08838453;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c53b2d8cb3d42896a11babdfa51a8af9ad3956ce9c22727e491a44739c557025ad94c39b1770fee073adf542c955395b72afbd6ad83bdb75c37b34ab49b43e1a817c6bec2f6aa9deb23dcef80c48fe8c211bb692f5941a2735e657fae4717728650f0dd8549088c68ca770d92fc7706f0e85c1edcfda64e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118f293fc369a55edb311439e8d7433133cc3c93ca4b7c8b089181230bc516c3728c7804dbb3ae98805701eb3bcdd5e7cd9469b1ec01907e70f694a77dba4053b19a229c680998d865ae5a9d7ef6929c9e66122c2ef7328efc06f9094c175d64101d512b0f78509e42b453157e8732b52d99e5d552ce2d69d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fcea45fcfca8c8db9976efd67f8e6d22d914d5764a8cfbb42e02cad558d10c28c4101bb37d63adf012c791550cb150a0c6d9e4daea84c54be39578951f16bb7dc2cc186dcb8844a029683ac7cc3fb373b27fa45dfb51d0a77e09d4833221bbbc32900c0fe5a6cec0e725fe85f10ba9c24a0c2ab79db736b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1686eaf6d933935088157618190b8833d77023fee3559f0cda3b5466ca3534837a0beb1dfce5d894f10d80cafe88d8979404a3c57d1ee2d4a6ca4c4e77d6a6b21f84dc7803dd5d340063b686e8d596a984c657da92b704eb19bad63925c4aeaae7970d8ddbf1c440e9b4dec2f6e0219fba201af799c736e7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fff26efb7e50e17d57d08bcc7b58248abe88f9d61452cd7e60a6c51d25751ab850123ea2ec9cd418d335262ed8626ff0b496bb8f7d0f6b9d686a27047fb0d8a0ff3819fa6a936e3e27c7c44feb43904e0b90d400f11eb81d2013f80fb9a10a0aba8847df3eb5ac12fdfc0deb654f7d8f8764d6b413bbcd9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192b0cf2ef2a81989121aecb3cd73ea254dd4af49bd381cce269e72f37febcf531eafc68f3d952f937c24c09f7c630af5758b3525b5e2cfae24881277c82d1d62a4ca26ef68c34b7c8c996b57a2831f60b7d8361c45a2967835230e365a01b45645538229be7801ed71b14f1fb45b8855090375b3f3c52abd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10030e03752d065a0b56db377eaa929ee4393071b47ea1a4a5cc3f43acfe084909110390fb8c2cc4b6570991bf4cdddda6e0891b2c782f9cb32fc611c4395fcb485ec62a49e85ac5fb4df13ab86a7e58611ad43037dc2cf05fc98ccf0679d2e487ec978570ed63be41ca80897c8463461318307723829c06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15657f991c434e9ea5828a3a2c193d6d134b4ae51e6a22f36974f4fcc5c19702aa8f74c61910d8d5e9b8dbd9cb533886e49668c18934d84c4cc19aa984fcc19dfa3f74197dd5fd52b40f48f4f0696c1f6eaa9be1eb12f32c2efb05013c29ef85c6942c4917c0dd3d85f90eb4275513f659f71925fdc7cdc39;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184126edb31ee226cff499178dea61e469c99f3f681c3877e27b4f7de4e96839b3b40a47d500d004ed5fd6afe33efdeea771d558c09d6c25533443ba84138ed2263c5ce5b8efe6b05f614dc2004e67a8c134693be9aabf3111799ec33cc15c5536a74f72543b66c92c906a22906b5b7c2f1e8ef8bd966ed92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1782dae05416d9935ba08241894b5fc91c72a3123ae70900a9c7f08d373b1ff45994ab414921b6c691d0a39736aad4b9cb7aa6e7f806ed60a2a9b3aea3bafcb874db66b927f2418fba7fc2fd4699bc0cdb650df2ace0829cfe4f6d36dc7edd1c69f8dea3cc75d926ca7de297f239df0afd74ff65413cfd463;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5251d8699c3949b78500d45a965a2313574c052da7b96b297ed4e84cb8ae127f495cb9a1128600babeca1629de4e64be239cb5bfe4dcaed94a9502f78a3c47fe3b9e471c7daa42aa811eb372be9e45aaa2283e14747864b6cbb87c86404d086099f600e7b9bf6e0c0509959d3a476d2c4f9965a430c3314;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0c0f491f4a5f802434a05670db6d47465934c2472c41b6d1eb06cc01e01d7b0aca53bbfb0fbf8fc42d324799c505b5338491daa3cd002475a2b62857b7feb0c134f441f39c18dfb9e56d7e2a04f9b60b19445efcf947fc1cd35e692b74e77c84bbe9cc30c108682a2a47924bd160a01a8889687afc26d40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111461ef72277c1b0daa8432e488184d1a8310db4f979819b620e84fa4bbeb96f5a2ab5fbc46cf3ee0336871e7de085188280b38977948a556c945dcbaab4010a4967a789794642e524c2d1d150812abb33c08d12a21a2f8a257aa60854af474c056ccd29c83a8eaa86cbb1f121f96c0e33e71d51f27dc3d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166a4c9c54faa21ca9cb0f9027d81ebaca422c001e658df798c1e1b78ef000c3c2a05da5a6b7c8a192f9c1c6575337a225a5aca56ba4e53cd16986dd1baa04593896076ce4b10ca3c4ec95e44541db7b520b16966a9376b19eaa271db7dd465f80e138bb8e5ddc3940a5d6c9b1f3484ac918533905d7ce7c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119ce9b53adc5f31e76df6b0f94617a451e0a3c5ac6070197f05668b768ab8273fcd0a8ee37dc61d1fc51e556c8b0b0e0147f01a91dcaced4231509de1afd9e241da9eeddf7da2bb545d60bc86e5241e94d0731a41356bf33a66fe92cb2c44ec66a467397c943748b14b13cfbcdb42b5385f8dec92d1e2f7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1218373dea348766f7e44b71ba09b036a59a7d836c3eeb6f62174fef10b3c17609827c67273449f4d18ca3ee428897095370b86b1be2e0371e4330e9fa58b258ce2d34ee1d427fcecc559bd660916d39a56761bad1257b88c4bb0c5b9c0d00de155ecaf3e752ec618780c251062cd0ece37a8a2be408eebd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8128a07ffa7b35246595745d2665f8e098e59d8bc26f3bcb7e34d476db0fc60f5e18047babe6d783bb98ace45201c36f01c74da039d4c26fb4ba8579ab68926f6047e70b2617819b15112f5cd679b9d1885917326298640219d21145c580fa6dc161126728e64c00efa920c365fac9193849dc91ff17c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f84390de76bbcc2e89b6127c940fde2798b996d48d18fed4016771dcda5c43b2f6a565134eb059317fffaef3e4a2eff3f04ea11da8e5e9a472c60cfb2c7116e48c3db2d90e5fc0c215f8dd308ef757987da97ad6a8df48e90712cc76f53f50d10ab35cb38733454a538d197f4c3e55b9037c18efcdbec36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18255cbe8e5703cf449a91db319649d44d22af47f580e4584537fee47cf536890861cade79ad2db5a9a396cb667b2c5d2ec9a7114444920e44e56a380aa371a7243dba43358fb63b3c392ed2dc309c0de683133250a1e575a9d49d2ede2b36e60846a86c3c7731073325530bd90012b94767c72ddc8ce2b3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc03602db64d98474b1248db09d00e6ae3d8fff50f454cfcbd8bbf4251da806fe3b9963a020e2acea7667b36d323bb09f6df90cc636c78b622fafc9bb3ba8d4e1b88cc96bee3c06f03e60d7e6a0d81386e10b4d480fc476104bc871f7c75342cb7e0d6ec01168f2c19bb39283f15c8ec66ac3d081575e9451;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15867353dfb04cda2750ff4cc08a07727ce707a3a82d8ebf66cc80506201dd1bef44e41c71fe6dc11e216fca8e24fd835f5c7ed41624fc88c18d3083be2805bf81759f716c768c54517484f1c555531a69acdb477a197bf5181e7006f25b41c2ad7646caea90c954f2386228085a5c48475382be177849824;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48da20a6121d5a9de9f831c81df01d03250e82e35eb82f578a58f52da210ee230956cf8d5f278b997bf9a31fbe05788f2012598cd80ddbc08927e39531735008d69a95c79dd3da587bd07b59200ee1374bd1f3a75d14fc06d136c390472c1674dbf16cbb9e3788a52bb88d1a67539ffb8b2c3c6f18f72e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115b349f36b59e1dac3bc3d42698f54c6f6a9d7c080c6c44919d31f5a1abacb96e009296dd2bee3396a749193507422ebe97cf065cbdc3446ed63d55a602958c1fb7d9de80c7245bc415d2ea1f2b711016993fd04da42d5fc1661454697e2239a8cbfa3b705c61b05f5a9cf5d8229f1e153bd3c6fb6cdfb14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1181aa83037af41dcf6642f7d5ad3fb11647753c996bde628ab12fe8b4443a46c9f7918625acea68f0b43898fa9c735415ea5ebd2e7390a3850ee81e7f1fcf0b2195c751b2f1a1f7d40fb42b8486fd06d425e8ae227ee31f521e5f2dcc96cc98bf662419cbc1b1176666885d32c33745cb63098d2b68702da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae3a4c6a1a9aa2d04a6c971c3a51af350b403da2c4934f97ca816a3683485b21140766f05b29d0fa144adb6f75086e2f1fabcd6d30555b03490b5cf9739769d8c2a88f3e205bafc93cf0cb356f05a0942663114ef2fe15adef92ccaa3f71fd0e3d7887c12008926b97183fc3b438c7bfb47243d97b4657ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a378f433ad0882fa7b5deead130e75d37e2515b525ced956d1bcd84633a04278b0ad1ec9fb1f9ea47cb4865e09d25c3b6245c92dab6037e49a936632ea33fb79384e9615b28b8ffbf76163c49f168d480efcb05018dcfe8844a710999ad3f2a38a4093a5c5d7e9a09181c93fe59167ec1a58d9bf9550593e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aab665ec2e3c41b475cbbed272e273fbc7ca0bd7b3cecd61c94f4238a2a4898c8352f4a479c9edd032732703adfc03b27b32db1e1c05986d79561c1e513a71db1e4cb1e34cc4677942ce4b2a8a78f32d69c75911cc2a1bac12cb4f37166e0bc6ee606f1c83285a807f5c8e5d8dfb3ed582c90c728813a14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4d5fb37ed31857b083b1e4f9532b9816bb2d2e403e95a817663932285bd1be024b7e9d47578b6c7471af90708e36b3045d27a0135742d5c03cfc3669f5c5a87c9c6ab5940ee202fc5f7df9999ff041d8cacc7463e56019ddfcf92153b7568b32c3198d6274164cd3462903a39cce9f33f33915702cbd5d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146a8a62689d38623e06da1efdb609e75a62e1fb90bb80396a42e13eeca257f51621c449b086373cd4d979ec5232fb310590211d09c63cc1df11bf59111e75cd9e32d6f1a04c724acc01b765c6d66af7e636c3c08a8a52eeefdb9dfa9990bb29aae3b09e4627ac980f5196a9174ea03d38726b774443f6306;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14eeef1d4e69fa68e1a970a868ac8997ddd658ecf1ac9853fcd80069e668c60e29361edafa7413ecb74ba623e17d6bde32eb539f7dcd03502dfb5c0fa731f1fe1f13874e76209e4d6fdb5a6156aca8f39c9725d2aaef9c3ce018ffff61f600a1357def62086d10d8662161402422cbbeba25b636f0a9d4552;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100c05dad57f63120aad1eece2a6f19b561e73058a5cc277ec03a2cd91ce16fba58837b06778521ac5a1488b0575e36f6acd16cc47e9346dcd344cff972a57983c1fe169a826696c82435562a177974b352b79fa520da265fd931952450d059f425d887f7b39cadc798f65d112985194689f29d1cf23d0b10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d12cbacf06bdc92579481793a04b8c5dc23dd9d68121c7c084cec5e3bd143406b4f9447e7ed0f7344bf9ced280c23d383b40aa6fc7dd571614b943f1eae403c2e3aedc55a11a41e56bbb79857cc6552101d1c1df2bc048e5a75c45da77186b68bee96589452302e611179809841eb9bb04e34b10acea9e94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h225e9257cb680303d2a9d7cd045f9cf5bb797858540b47b60d053da5489ecbf851576d6042ad385ceacb92d6d138e88cdc9e38250f3d28b4a21b470cd59296b22690140955eed7e6c85924c3c203fdbd45e4d74397b4678852981226450b08694582934768b9d886ae62bc92479ce887283f1b83a03151cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109f991e41d5256a0bf9affe60956e74306b33decba9677cb3dcb4d5844b7253eaeb8e3b1ea37717210f13a00011df9cee4ab2c697dbec55a3ca897a0bd0735ee72827e547bbd52df4b3c71ab529e542df4f06a4b7788e1acc77ccfd92184b5b674e61a3fbb38f2151350b9e78371ff5f33065d4dfd88243d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153abc70665b079747bf93fde5ab4c61e279e93f6dd1abfd4fa5ef76aba731ffa172fcf5365e859ddd157841fbc3e7fb224e8a8c5ce9344ae2aafd74c2cc4c8558b43f11609dc7df2cc4bdc7bb60d303ba8a0b7a6941d86e7fca1d57510082463615d0fc912ef9b0fcafdc88c235b558f1ff1f16f9a796432;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cd8f3da15ba84fbcdd07d24bac95b9dfce553fb6023cf66a070080945c2e394b8e4f342c12c78a8e25bbd32a68f3b448b1499ff49cf46db87e4d37bd31e5c61c2fd26fadc341b13bd064f52894162060f5bc4a7ae3990d078c92f9203e78a5714a92e2113ac3f2f4bdbd3cbf8f751b7a38d36e5226175fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101e931420f961b5a738cedb938dc728929555ccb38739317d7c84ec27c856ab230f36692824d56c0c8ff806632f75aedae1dd6e7687986181aa29651f6b993993c13a3fa48f1b66922ec2cac4b9198b54966ca42cee0ebfdf196048987589e8acff4129434dbaaf56c42b47b887b5cc40b19ef85810c7bad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91804ba6e8e0817a3a4c6d1e47edffa4513d1d09acd0dbc24855fd497b2810880ad3372c2a3b2d2a97ffe7a9539c78b8beed2f277dfb4871c6be1532d42e1e21f5157ec85a38338165e32978969bbb5ae9be703f2d4b3fed2e53dd99ef569a7f574eab236231412fa3b0a7f32da0b52f1ad4fda42268e06a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c0d0b3a9b9f048dd1e6d277da5b10e0d612e887acaa071681b32f8968d1ae66c5f757af4b2e2f27ff5ee28bcd283993b31272f106752aa7f2755045542a81a98639f75f63cdee2e4b1f78e3fcc0ce804d32cafc8d79f9bab905e6d3a523a63d03c7f6dbb815e3f9184d24a76142ab2c5c3fe339fbddf015;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9d884084e8529f37eefb714835b0ee699eefa626cf9f93b5ee7540af3ad367fb5e050e4d88f31df4ddc12bea6c0baf729d0fa8b4561575997503adedbb0d4da467061bb0d1517a49f5322afd5c3015daedc60f6579e1a51e1c8b3d4650fe44ef0dad75bba6fa96ea21cf7ed5a7daab3996102cab42f7ab0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h704ed159926768d3614c35dfbc79b7280ab8ffffda46910c5f0d8118666573e79c11dc99077a18a4d83df89f1d337664c130c42ecbaba4028ee64b906bc1d8dd8c2442104a1a50a4340e0fa18e05980f2e50965af7250e9f451f9f1b43fb791c10758b1cd5de9125557cd6fe56bf1b840b7f6713d91ad1b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b17ceadb34b1e026cd0fc82c1169edfe890ee80de24fb7382e6136879c24b6533add6f6a92c218b478575a964bd4322a5245fe882c933c1def2e0257f9069b916f993e85b11c95c3aac9ec96ede489e0811262311653d446d7416fd66c8279d067f7eac5bcccc70ed5dcb66c1ec9753146be9516c43bcf4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108c2bd2e6d505c5a1a9ebbb6ecbfcedabdc5927985746043ab89a4c22619be62da93f68497e1e04a4ae4341e470dc1cea37dfe13a178b92ccc702aa2d9a22cdc9ed7b6a578216561ecf9b0183a09022dc25cc974fd20803b36ca803c1daf0675ecb9b25997af64677c314b5fdea1cfe3652172b286077bbc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ba76f4878603bac2d786301b530410330d32d1d168a9d3c4cefd311ea96f6504be59b80eb4e34c5c108f82d4cb094a3c3e7ab7b15a74b484958eee5b90603d245840dfea97c6e24c716c8501e0491f2b5395cfb944a36bad01f1787c7b63783d62474293782fbe2e52a90c05a5a95084358011943e2ffb3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a59e9137798711884754ffa99876cd67bd211c7d7ed17f4ba41fdc5d197cbeff000627de53c45fbeac6f5ab0dbdaefc277d99080e3f11789b9d7e63da12d2877ef415ad82b469c232b74df8112276294e7f08def94b0b16119cbd1e89247f2b7ca6c39daef81798c4e52d1c5af7b63c06b5b88d8c85b97c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fcf83402b8aa4649d602795172275be690a6e1cb0e795d22d71787f6df1ac4a0ba1e0ab5267eb0ada6b1a23c111c1005f4bcc0fbe90427ee0f0534e7a41e229495308494cf24764d5e9a567b08710f08ff571a6ebb037ef199fa6bbf2968a665c6e7102c34d5fbec34e4676a41de383072cd56e627b632e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9853518b4dd311bc73e11a5af200e9839eac458bf4255e074d0a42333673a8be71830c22d9fca6b1fe1be9905dcec02093d856558079744ce596d5fe90a6f7cfe89b0bd76b2911be5dc6432e448a849ccc63aecf3fdd5c7c335dab129ff03766e1fe0fd6c7669d46f138ebadc82da41cdce31991e187a5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b1a09b77743214a968c4dea708ec2402ac92bccf361bbcefc48a4e8c4aa566e3b60a2d537aad89d63a56a8e68dd743a9c81022779ea7a3e499b59f98241c1204dd3fa79c28e532e9db8787cc7e1f48b330255aff54482d1daf820b48a304889343778ae721a2aef394e2901ed849eb6a5f7fb5e0c09d6262;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16765c3b43466073900fa321ad26f403ba20eb1f3ce1be51a17d682ee58b5739af0b9cffb6aae99cac2007a32dc0a8a9afcf0e2d8decfe5e1cbcaf28588f12152e99a69712fa5c87a4f0f84d769026c95552afee5c7ec9189fbf3be3e7af57afb33189c655fe4466aa8f88b7713612dfaf5bdcda9f3b5aa30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a96005c087f0b5f17b3e562d35d0b6e9a6e2421450b754f03e6938f1bb7affaed66a8ad81a7c5e3946e9b2d829767316034c1560968efcbe4699fd0ffa9fe230fdc5b1501981e7c919cbd836e92d199e23547f9dd28e0a0ef6a2abce4d27e1944fbba6fcb2309a12a911fcdbb16221e7803638e35b9a811;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2c0f40c35ffa086e350edf84d22a31153dc8e9b36c7177ee9c71ffabe294707ce3e71350e61d4b7d143e55682b902e428d63b10139fb90344746ba7f8164f6a9737cb96082946ea236af32c9c05771a2381433d3a09dd1256950149dadf7ca7e09b3a8a6f08f66a6e271e2674bfbcd22df1c65c655e44f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f65e7aca3401bdd9c8a0a1bade7a3c1d553b27f7fb9cdad6d88d75e76d1936f97e57ebee44d348e2af280e1ce84fac143f8c4a864ecca6d120beeeade18ff934fea8c36f57380661f116f9245aadf4e9ebe4e800fed29cfa2085a7d9e19cd2985c97cb3c39f84a0d3d33f32cf510ce0f83c87e6f71a6e9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b1f07c8f10b4d74bfcaf396decc7132194706defc327319aad079c6abbbfeb8926d0117ed2dad4bdcab82832bc04f29afdc1dffbb8eadf2e0e2a69108de8f80511aadfc818cb3915ccd037dee0bc55fe2a408eb4d814bfa187de82aec804c7c86b605648e4369d750c3d01c82533b5704ad64871be8e756;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb29d34b51347ad0aa55f4b1db42b966c32692dc150b99a8cb1bc5e378f51d435ba263a074194868ce51bc7f84c34e1ad35756ecee0464fb1a13a7d96621d648908685df1d5edaf73857ad119a51b418e2951197ce010e2585d0a6a6002d9c3b12b3f00bce000e39207978962273000bf45fa3c19ccddc9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7832a6db4ca02964e866f97495d77593bf109092775f6b69b6e820e9d0572c5ba9083e40b3ec3a0a4be3f2f01ecc78b250843d5e684add8c48845a2e7c8fd9ce2ff8453e67ffaefb51b39f82c4f59ebf6ea6b9483b6cfd14874189601d6a813a6e74eb3cbc0078e415dde4fe2f741e3d343cfea5ac0d356d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4d27bd3351d445dc613e01ed78ee9fcd8835e263e157b663b96bbbb3c1b707bc858ea657b86f254085ec15e0caa0dd9ac74b4ccfab65149f511eb57d56da41d9e19047f8edb249653b0e9b5e994bc3809a3c71c13c339dbc4b6ec1d011e45c6472baaa60ca378bb0f81dbf2678a617c4bc7404dea7a64a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e5a172aef8f6fdb5fec92823512e18b0606e5accc69894743499c2d7596b6828e818a2c4b54281c59e64688bf983dd4994c19f9958987d0cb4145955b2ff6460eb828d61ccbde635e2e34d7aa2a57c92923ce4ccf0579620f46303014661386da7a7366560c241bafd970b95da0ed4696bd259fd2dd5cfa5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24c6b0eae0f1a57e621e1d0ea14f594956a4d7406a0927194b5bce486630936002b49d1121dca51f058f2a6e5e6cd5510dcc35a4c42c8acf9a838238a5764e8017f3b5d81cf1a7c5e1f7a168754906077b96bbe8c1615fb63257946dfc1557056761b20b1760ec015191083e51d010c8a8006c2cd7cbbbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5823570089c4d63050db7c1db5bd94542087e351638fbb8e2755347092069759180d0684bef1003be1a427e031aa978d497a459b9c63468642d7d861455f6093d8b018aeae6e7efda53d9fb782c65614e2ae63622024c7a06d57ba7b696b82162705bcfd5d85e1e818f3cd786930d260205d30394669a48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb22ead6dd6621367ef60e6e2fea6f5bd9c5081301b51d1bea7509cb16a70b5e3213458d8fcfd6bb85a609e748cd1ada4b335ea967965cf091e63f9593c83203a9276c125c742b6f0b6077641f75f8cc8478e6823c0e6cbb4809f0df86498a8504bbb4741aaffd430b82aa0daf431699b6a3cf851bd0d449b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5aae2c2915e1951c4ea4b6e3b6182d7b1559a5452f98b1412d9caa3ac5d00c4bbaa04e3577ea6a685ca594aa440d557268dbe621dd3146e5c58be8b8ae0b4e6d855a69a5c205312bcaae881283b29958c747a75a3c042aec43b8f21a7acac30b61db3d1d4676523edbe105f142c7e048266bf7a60126aa31;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185fedb18427aa1f48a0d622c4ba83803bc322aac5bdc18296ad0fcfbbe4235305fd1dbb1a13c93cad99bd75d3a41a0066ca828e7165b205e217d331b58fee627a193b64f0c20367b29ec5a0ba1ea2885d7a1de53d7f4bfa6b3ebb8ffb2cefd78d5348b0a95249b41c140d8a93f47ac8d6eb79423e5752689;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17677e3b0cd559fde5c287ef590d9bde257a24aff90a5abf479b81a5b4f0da12205d080898851009e517518f7252a0697ee57e34a34db6f715363f8f729497b036c46425304b3b22af74b222b02ab3b40cfb93d8588d65a840997a8d5c3c2a1cfe3a1109fd4e284c8d50eb143f022525a8926484b5939ef56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1355fb3c15954f97175f8edc10355cf2bf0ad365c712d708e965baeebf35c985aa9417910d6ac26fde4db46df9b243b597d93bcda8b3b14d86184af17e03e0f4ed618bdd4f45b90b83b9a68c011578a92fa31c32a09f87d384ccb0b6795e5d9696601010e29d37dad9f418c14866c8483df880c8a1c45dd38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habd878577d9c5eb8dca56d6598f10df63c8e71d623bf28080779c243861700556d514324129e334d3a68a5b0a6890b3be986edde14fc4fc01ec13a21bbc720f3876ba19dd03a00589738dfef954a35130dd248ac8d551bf36594c8ab5beb8defdcd3eae885b18fe01f65a4a8d8cba5aaced218b890193c5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f7a05f72ef8042b3cf7ca05f7e05fab1bdd34c5c6b7ab11a0c6452d4142ba16015faf32c0c5ad92656a5495c3dfca0badf1289974cf34ce138e693d0e31f84f8f79236158dcb83b0a0b8fd70dc92bcfecba885fea70c0b5c33539a0c9e2218db3ce2a50cc93323657558cdf718114019121a4e53ced5151;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec04e63a72da9f8cb016744fc25fd9cc6fc04eb7a8631af5996860add5d86e57660a0942e6e33ce58ab11ac6158d9c30d869946738f494c3423491e268a9f032bd765c29225516ffbda4462499bb62e718760cbecdc6b0a3ff83058455762720208a27b8b7001ea2d6ee739e02acf27d745b6c7f86eb0ab8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6546fa126b41e30437f42305cd95488165c46565ca4ad2c03977aff3c051a541cde579377a77cec91f164a18ccf37a342a1e52f4b647427145b9e3a018d2696e61490b203bb85b572e5bc1b44577c925deb80c215661d66bdee7006a804b27a07de735a90d8307eadc87f8a6758eeb279dc16f1d940429cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bf2806f990c94df5425670f6fdbf56c37a496c6da4c0976d9d2f0a229118cea40c250c108cf96f3111c4e6e996974bab968bd8d2274dfd12c1ffa09ea21427aa65892ac0469786bf1729e223406d1a3a970b85e142a28cf47b4050626bb0ce410dbf054e5327b8feae817edaaaa97d148f5ae82cd6e5aae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16935aa500c71ff6e941c759980f678da4ce707f6c96879fa4736ca959d37e9ea46643b22173d5e1c54b040d686e670d78c438aea1aace13bf6238b0bee42862862c8e0e2aa850a114183061b807d9433d4e45edb63bac7e1c6087228b05d05da08a9488ae5bae6242a092b640a4b59ee98af89fdeb2ee08a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1273703d88748346ec484422f082a2e7afc6edf20072400c79cad8391c23ffb2d7e22f854423876dd03bcd9ced95942072c249fb1eacf80969f98c0b707e823218ef6605cfa0464bb4cf5a59c2e5a96e3f71e235d27c800351e68ae31f4c328f4a4c61f503c44b2bdc74eefbffbee025b1e008be0e2c88b99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1086dfa856265decaf451031b15de49653a690362cd75710db0d1418ca60cd40511baf84df81ee4db31a15e06caca1e6150f725aa35fc14111671f195382ad76019dd74bf76e3a71c86295561df3b2d644973b64081088ffa81de189325b29bb7a8d12e196edaf1ed3a96202a30cc7d7eeb51f072d468634b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1535525a8fb185c54b7000d12e182c6dca376595b84463ed2349eca11f73ffacb2e7c5f67513cf64eed85920dc2982a27140e38cbfe812097d36d6332774cf4b10a618a4f55e9ee020deff3e5428e5cce3130d57247b0028811d65cbe11cef7b44fd5bae7e46919bb5e8515dcf20b1139e085eed1dae96d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14db796e1816539611e14346dd0ea907331569b83549d842a0dbea903f83304550e240e9c316d381605c9f23a5dd07fbe3e1a4f1f06e62351619bfede27cba4ef8ace9c302256cc8f0159eb333fe0fdfad7c1ba7b79f6c188bc2116cdeca61953d6f76a9c3c30d3d7838c23055c086460cf804d185c72dcae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118f33b3094bb3db1266618617e5857f7991f5971a9feb57b40dbeec79d9cf9c1f532eb51b568882e321f0858a316d1611c3f6f5f113c0bab6bf3d980c6c5b37bfe3345007f6fa47b4d0f484488e2d4b4d45a81c7672ecb057121c0615ae9f3c8cd5f2a8bb0096ace21a2aa12b49fcc126c7a74bd8f2c0f69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a58b314c34f0ec9a1e6fb266a995a906b1e3ca6129aee8ac7aec3cfeb5b1b7018503752c0a654f3afbab597be052cd82cc86e716c3a72eb887e8c7dab4744c1b4e916239060a74d84d59d4d3a9d44d415be0be52e4529098d8471189db260c395675d639c7d1e66176cf802c2abd5b316b2c6ee51af439e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heca216886e2016dbb57aa0e9f4e56d7d340e4232e35bd2a914bd4589b189686159728b9deda3a2b8e84b910a73d413f82e0df0a6b9e97ca66c9c3ba83b5aba4f3580a7e45f730254fbaf29a7decbca29ad75231c691e4f1ebdafd3dd247d46bb9053abc349388f4b78e24c75169778781cd2675f0efbbb4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11491a2feb4e3106be8d524b565a7c06d875a873c35858fd0e4011bc96abaec9b9ed0bba15a2cad8717efdbd6e7485359f33390a793f0b0899de710ba07ef1abbc2d16c18f984b3296cf2c0c94e989b022b28e1ac794407e195727533b5f69288e1e9b25d55d516ebbe16da945e05f19c7194cb97b47efac2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf978989c07103b5911530a3aeb8e2b4d2e24299f6e17d8cc22a79e71dd3929261e94b76c4e92f46fe7315a18c0210cb6ad407352f1f984ede97ff3197e1bcc5cce192dad6d14b4742b75b3c58af8ce283c863532260fbaf6e08eb4e6bbe4367777bb63b50a7e2bdf3538927497613b68198fb34bec7a5c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1695340df84f8196df786e9425a50c6269063359004e6db8efef02cc60acb2700023e5873375c575d06a0159b334733e7e73b089a6fc55c2eed8f25c58ea2f740ba61237d2f0367973f41a4e261a755fc36be4a3c5e215ea57d1d705412696628d526170aa76b1ed3bacf86d19587e2c3e1e61c01bb67a335;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c652fbc8565eb6b3b0e2dfb98fc98c21b5bc272d9fbacc2b067a0a425535ad3b43e56f1eaee5184af04f2031aa370a28611f10749c6112eca7a6982ab1e966745e688ea11ba2c3510d115912ea7019708c592b16aa5aa8ec792611f2db5a53abdb325487002bf5f4029283322587910238102ec3a660447d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14071c4cfb8aa49a11feecbb21c5142f3d8fed2b3a7c5af8ad312afdb65d83d47b2eb72ef497fb34f34f35115a269da05e02eb5f61cf2c2a06cdd374cbf59ffdf23ab18d584185be7d18d50d2481b5b9c8b43b1a59e5cebdd8b9205f8c0cccedbf4a736e65f3f0038be37e655466175cb89e4e569b180143;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0708aff1487e0dee898dfb1fbffba2669221f916d1fea974280ee6fc7379c35b53ce09f22d49fb7145720aa0482655683e2de5fa2cb4f2705bc2aae9710df55a742b4aa16c14bae45d87c515d44de059cf3017ff86cbb074ddfc241fd015d90e76a13d92c57f64d3cf57e5c88cffebdb7db502827f634b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e53433d3ed3e9014b1613c64a672bf6d5414859b6e4f7d8f246e27992d022639b03f0b512858714c4f3afd039ccd16fc166546c8eba637e8d641d2ed29c72753156766435ca10340d32ed39ef5a70834637351642dc8b967aec1e97e8b9cac9bb48dcb73c9d2112d50b090b32160022d07d976bb19a7d9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84c70d6d438cc29eac69747ae56099cddca4a736e68c49571de974b6981e71846496774c89c1117ee6c01cd48204690c5761f73606fab243c57dfefd7e771df7201699622693d775f7fb60ddc79278f1dfeb47d3a3801d0a1230d9db80cb854bbab07a61364890cb219062d286b814a8da88ee6e4c9a7a5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h334684f50a0298cfa8837dd85ea5002e9ce8f5a8d3ee52007b6a5004c9a20f0a4a515f16e968b16f35ca93caa8b9e083d2e2568623fc46aa51670ab0f9130120bbf5c66595eade312ecdc32181a7dd1965e2a60402d369f9efe54856c46e1e708dcec132d124c237acbfbd681054110066373f621c57bd28;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cbfcd2e87a7cdfaf33a2564b3a02a000151d79b02263b66870427fbfeea7d7a70ffbce2c3affb6511f9f022a5afd55f4b68e6774329f4b206d26159b93e722aad0fb354d1263be2349d390f825a6f0fdac023de49997a3cd68110ea42866243989ca74fd4ba8ca0f06aa12602566f41a64bbe2b0f555588;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a04f8a6fbb18a05cea09a85ad92ea905e0baae6b254d4448ff49003c7093f9ba0e4f3c95431b0ac91fa779fd558b01f4591cce8e76d9b2394371485757303d3a75478ceac6edec630761af8f2ea7cb724381001c93b5cc3b72706afa2b565a88011d80e82b0b367add3dab3dfb91e773940a1f27ac45113;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c71623c5a77d9aa2e35717c1b22bb045e1df618b0dda721f0c4abb884d072e5dfb77edf6ea3a4f5bf7eac59a8fe2ed88a78067b8b2cfd0c5e7fdfc64331150074ebc0470998c97b43a4d3c7ffa5243842590bc5f8050a2447bfbf8066ff744ba704e2ced866d0b057da149567854c5d9860036d4a820d9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1caaee8ca033822a7c24e32365d57d974bafece0f75ab3370cfae03ff2a71024709a118e154bf25f556e289a2e2e7f727dfabc3783275fc448d8842c837e2629f804c8097aaff58a37b2cf5f2de9f5ed3e705ab3c9513fdb0e9a113d1a5e4baa836f4f330464c5af92a3b10c5e66c3fa1722a764f2e80f720;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169131c4eb911e9e33e3039d4c79fa9ee59f81ffba5dbb2364711497ce67202822ed38f00e7e98065f8073311047c32242025d199d18486f2fb6a63c59886112751475d66a9b921ffb497e36dcf3223284d9d442d328c9e919b9e09325576b8cb846b8375ad18557e1d7ea7a072cbcd84137c363158ee7b3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f60240d84a94e76c93ab4d1955e7dc677b66ce053693976512b09b1e0227dceca1af9a8f570e279cf62d5f5b271af1023dcaa488e4f986f89d4d817f87832aee6b0ea85fcef3622234042aebd8fd3ae170223264cbe52a6dd27447e41d9020a91769b2a188498fb7a4058ffa3f6af4b7eca0fc1ff8348cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfeac00740bab8b36b2ffa484063b599c36e906e7a0ede0d907766ca2067c7b13fa9530d6598f9a448f4cc03fb8e5fe71316eeb9da8616cc4682675b3a3b95e3ed277060e978cc4b96efb17bcadbc256fe75d1e62fb01c9122cb74b0aa2cf59a00e7dbbe2329aa3c4189c185ab7c2e41c2847aa4c6b8b7fad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b492adc7e3c36abba5e4543dd6a05181887a40bbb5a13a4ce876392815c1c43b9130c8d9a38f45a1d11e0cd7726eb8577bbe1cc18bb85d276a3b730e295666e6d34f041a3924f8146ae4ed0bf70f52ab536fbad5023a35010e5768b8b7f4e5a8b704dad6e3a77ac48a6e153b970e55dd4fa4e356e37dd1f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf365d9ff52aa90c075f850aada2ed0290703fd1cace7db396be4bc9920493407b4162d2ef410b61f909bc81e8c6023ce6498a767eaffbcf67a61463b4682a8cc89b5e5a5e5d3acfb539d5e1379b77af87273a78e10210271fd31222d706bf3c44cf2d7939fce21cc237e9147773744a2fd261bbeabbfdef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1967818b03e4937240dea5ad3cbb2024282f8be43713d287a6d00deedf9c416df8f4ec715620c173dbcf3b957dcf652bd012bed3f7dc476f62345f59d7a262acb79cb3b2ecf3474763ab7ccdacf0e829a6dd4dd816cde2c305ffd917933a6a7cba74bb2d7753430a1230133a22b87c21c1a809498b1d98e98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10925f0da6e5ef2923a22f6521475bd72d5b7cf9587835e5bea53f7ceddc8773a443cdfe2e93cbcf13009652f672bbb716dca63a48b9fefb7a78406dade18602b029440f45758677610d1e4241661c9ecc51c89f67be36047714cf330d3c693603b0c391b531b952c4be6ff0c6f53b8399398dd4479e1913c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98eeda903dcbb80d3a4bc4c28c0e211d123ed0d0b737c55bb7110daad4954e51b836dff68fa45dc4f02ca41776cccc9293c3c70b019c89bf342857f15bd50be6e5564b957f6e95012a3ab2437f293be2ec8667cfd4fcad68b145435d697664871fbbf464804c10633e0686cbe537d3c7dac1bae91aca96c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee5cf5c936ba4fab85624e713926998e0ddb9c8f5de0090702b822475dd45aab4a0f4b67dd00b3804cd185782fa515eae3c38b03c420cfeb0753c268ec28026193fb37c9ab9286b40d726a525988eb8a360c28eabd3035e5818ba38f3e8d8de9d757cd4083d500d1f9f317ec6051dfc971a9de2ddaa66be4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c2051d02acf3dc88c17a6585c635ae048d75c15eecdcb4057545f1087eec2b9ef23cb5b8bcd1c6cdc761c9522ea1230a3af20eac440d67fbd764ebf5e39fd19d9f50c599dc082ca0a31f3fbf61e8613a79a3e6f6bd35d6a0b3a8fadddf8cfc980cfe39c9915d7903b51dbccd293756ae95b0a3e2a7bc43f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1992f82fba06ee81b2662ae60a9a1399dcbe710246e336742dc9400f221c79de2074a0e3388e66b540e874bd269ef0032042bb13fcc9f5d87747d8fa25640da70f5db770ddfa568391fe328e7887bd938f58a42b6aa27d71a9e429f657bdb099d413cd79a4ac18bba19edec78c1f1ee7358da5d627057f2a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1046f029b1d2f914ed8b714b32ea4ebb2df19d00e31501f9d7cf1f683b1d0d39836105c35572a2788fbb55cd32b4328ff4aaf60d9e11f146df1b9ca44c4e2f8521e92e8d37574a32969bc4a8385b2eedf67c3a69cee8f02cfa7a61001730b691c4d08aade6e6ab09a6576013eee5583ab6c95d57e70d6efc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dacf2f69dbc623f2acf1b8f350fd5804b697d87030b808c8a1773996fbdd96705cbf00d3f4ccb74a7c6860660b9c0eb09149c08960e5f81def6c77e8f8e448215d6ac18186aac052cfc381316c297a451440fe8e5e6afa33ae5bea86306a93cb89ecfb700edba1de752d130e64f16dad4ec559a27f7ce89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4d30c87f01303eaf280852d1074f48bd4f76e8f23547ccc1defa2d3ec0a6c24b7362fbf2305f184ba9fc71db3da8a383325ee1de59b66cdfa86dd59ea76251633a634a3e7edec27bf893e968f5a91fac461adccb1612d598c9378340c853eba43aabee279034f28a3ce500ad497ee8cf76e45791677a9a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4fd14f4fff153e289647c1b115038932d8c7edbdfaf45a63b827ab23bac81d2c2531c1ca1226aea78330a24d61ad66e6e4ce17a239ce8ce38960b0e4a95155b877a84e13d3067934cc9f322c5c168e3da95054813f47afc05e5022a8dd495f54660c4f83a3b1a38bfd022bf0826def3fef7d33bdfdc4f36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140a7057fadbfc4a2f006311645485644b849ecd377dd93275c11a9afadccc8df8e2633cef81c34c4f810f25958892607e24d409e193d972d3ae751fda31e7cefba3773c50d1df13d5109ca761358687d75980afd087fd5739c22dcfd8f4163304caa26aab38bd4784fd3c58a130d2389db480843d6e5cb77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha38827ba6cf15c55cb455046dde04eff15003d5e07adb42710ed6f319bedc49d4d969b2ae6f098b8e7e88cfcbbcb3a1d7196e3ecec3c2e06c9770d771eab71a934f036ddf08a5beb3067b473dc5b53214008a63a71f6936b1ad95464a3ecbacc3acba3db7271537f6687fb1a7c5b97fc48d3e84cece069e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h904e0041705037455cd42f5cfe6091ac054ddd8bb36d27f555cec55dca8aacddc0efa731b089b1e9e2635cf2271e7888579d14c9e2749f1175fc5e463f0d14fc89d16dc98edc10d2bd57045eddf8956559f767af2eb951fa57f14569800596ece7667bb325ac301d952944580a9b54ca0dd37bb051fe5290;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ed1d5c05486010d7bfc205461acecff55739514d1918de6b58cf2156987f2506f3b7a5a76f65635b759e1648d3d40f36973ce981f52c294f56fdbd7832c19064157b68ca675f39981277d55a43a964ddcc7a61ed76303c68f3fa27716f4291cd5c141e2c7e0e0d81d45daa4fc997e77005916acaa28694;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed0859b0168ec892474fd5227c3a9b2baa4da47a44c59ba442e93bbe9bc4d06dc06bf6237981a8c3f7f564e73c285f7019bef2f439dc817b9b77600e8e7c8e462ed9340a555ec7d2c29041cf26e69aa884d065eb48806415dfc9244a7fb9df893d7c5112b7e8a8588bf4ba71e49e9dee0050c8a9e3369dc3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5c4b2cdc99917794b5f54a17376f24d53ad9b134fd33222060f3cae88b315392beb3f2fe6b30ec040663ae72384e4d6bdab1bd24b758a25e7200c97342b575a91555cd93931686703c7671b0d5ef0e437ec1a864311491a698ad0664d9fe8acf85187a1733b06dd6db9a15d532dc2c739a90556b741fc44;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1727ff23af682b7c4c320edb6036fc3b7adaf1ed5a5918a3426cf82682480f7be9eabf9427f30bedec07b3db0f75e2a3c96170f58e7c6e6bc1e3e4edebc4393db499073335e964681b3cfc648c462eaf5a0b385220cd51ea97ccf21e24822cbd9922d5b20ac69242f4644ebcd0f5bef0efa5148a60164fad3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce0ae6822ed1d99f6f3134cce7928f64cf82bf9b2a65c8bc47bcfe60f8e6cbc4862e12bdba438047376472974a2ec15ffa22919695e1a25e04afb98c1bb7d645a747d1519a798ca81cad6a8087e2a905ce5c20c32492f49385a0e9b791cc5c0dcbbc803fd3b9ad9760f70abb8e1b2e32e0c9d7ea4e97f8c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h204afffe1ceb70d35dcb5bde3d28995cc59c52fc6a0e975b1c5007e5d7b57fe0ece44fece55999ac2729879306ee181b6375201ba2b5711f9b83f4fe35d4fd4daecfaeacc4188919998522b29606a209a99470398ad7154426d5a31dc93e2f6566304f5dc0064856da297bd639898ce86f44fc8b82903938;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1831d895f7fc1ccb314f2069dda750d42feb17c17a64fe5ecb3142725302d065d8a465789d6790981dc75c1d7761c339f3d1f57204f3fb07809a709b92b9058fa1716ca88ac6ff173a12ab048d0918d8e2e12df9b5b0677282e470cafe64b254fdd0a21ecf7a6e11181bba8b6b20b1b45f1c3797405df9384;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f645ac03ca2e341e8cdd8c75f77d4d65f7480f460ba978f8a93b0127bd68a4a834eeb06fe43602c320df3801c6fbf4c72a3184d8df5eaf1a176b876354f4c5e83a7a8ae5f48af229e7928d6ba9f9f3751d89efe1188340906558a86e745089ddf2dd4279f44da6944027dc54560dd6d30749b6b0ef158fb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a689ad61095068d91fb9bb112ea8338e89c3f2297174f18c34e3df27ea7e4063c64199fd7cee30021083f06e6ef4e1dcac0a617319858c96d78fadb89288821fbc9791d05e6cfe718f69a671cd80546cfe9535e44cb2345bcb5990d47fbf4ed7b30eb89e3d07a950838804b120ae5f392bfd337782f9845b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he00574ddd94d2f14bcf9df76f0ba4dcae3709f3e89fb3dfe1ac7d57a52d3e09847466ec47ef2a6ddd0a268ed9f081a7bcf879c0e1dfef26cd5269082bd1fdb373c574a477ea3dd89a6bc933656226daa990bce62aa9f94b2cd899193344ccbac4b744c03e4c04eb0e22c9c6c156ffe5613d687a6067c468a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfbb6b2d9d2b73af2f0c9bf6792d5eb279d6e752c142365509f80f985486a16ed52764e87df06190ec14b040b90d4f709d83354351f501a9cb51fce1ee15cc214ac5c35754bfab0bf6ca9ee433cf3ae643e4e677074bd9a6b0b08a607f48f6715eacb73adac946b89ce71a19c99268d3587083cfedc1c558;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d9ce86270e9c19762e2d12a3e7cc9bb3d2fb469f21f353df9217b10709e6713d7d19feee72163b5365eea0072de95f333e888e42ad9a3bd8d8d0c020ce2c4b3b7d87ab402ae0cf4e77f8573d9c836d15d212dd70fcb14cc8042b0ccd90a7a8c54534843ff95c93e9e1a5a4e0823235aa79809301c46b3dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h334d3c671be8265e4de3510f74e15892ef09db83a2c5b9afef91adb656ac4531f4cdd414c6de250db2f5a008c4af08791d06749dc6d2547c2e3e948fae7e6b198f9fac8ba9e4bb329b22664588c971bdc5d8ddb41e2b8450904ac879e6f30dd48ceadb83eb14e9119f64898a5dfbe4cdc90a4fcd2fc0ae48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb18ef007d039ee270113b6139f5de1aa8f83153d64e2d723f60f6531eb539ae638e30e24320b24e150d4d99078fdc83d739071f788e4f4e5005542431f13bb372713d8f7aaf9d8ef21bc5e98b39ef5add40d5e7d6ecb7cfc7c59c22d8a1a2e5b21cc04d4a0b90f4c5993a97424c50611f93f094786b39f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b908bb140e5c06260535472aa009714abf38004f8829c4ddc523334b073885b38a47549a193480c4f9448188a1b4dbd8538a084ad720556d2d89075b1262ac5216ce93772d9349d4ef2bf8601946e07197c8c9803d2290540a4b3b57cb10e9b49f852a356d6a6ca6c3a4bfda165b80bee853a82153eade5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8d321c50f7e1bc071036f45e89a2156ed24b6152f6caa6d82c6d4fd0396a0c2e06bbe4f04dc57cfc0563a13c2785fd05bacfc53afe9ccfdd0e76bd8ac8a2854f0da4cef81c304ac8ac94fa2dd5f8952e3d237774a6b60840dfe9d884b1edbce41cd00863b2b56964027f644ade06af37a60b3806df62816;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc130fe31b9e052ff8dd775a90775cda9c0924e86384796774a8b83280550aad63b0a7c3dcf85634d3dd73655f9a0a8d04cbc3e81424c1ede25c965954fbbc927255bf2f91c3e382b70a38073901e5add47e5495aa439b74a8c4bed4a9322e6799f6d4cd3dc9fd189a32a70446dc7263b1007e2c779fc23d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135b02f2fb6a19d04a2a77979bfb678300f723ec0453e56bca7e72ae61b169094eae22c4ac2dff5250d9faf15d8dc6df96d56fe3eb93587f195fddb8e87931146f9ad0de4c5a95b952714f0c3757ca90fd71e6856e0cebb9981a02b351442e387b1d850af3b358766345479b8d4c51e1aa62ebca5de6d5ce2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106480b8f865f6c9791b2a1bc1cc7f249348db4422fa0b77508b661c84594fcfa8f67c7edfefe8b559e9e2859584b541a78a5f085153fb462ad1c636acff42a38f6294ade42e46822bc8e05960cd93efb0e3b4fefde417fcf9113b0588ebf83c47ea0b1706277c3b9204c9b92af8d93fd185043fd3278581b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d024d8c90f5ab0eff0af53bddaf569557a9e4ae6f336418f651eef0cb509d831d89dc960c4a4a5f4d6e5cdae42893862d66cbfc33b2df6cdab9401714e0d059998b134de538197cc09c898706c0b4eb8c174429f975452dedad1b6e2de8bde0aacf422189b75212985ebd92aef49ce9591ed0b5ad508c94a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadfc13b68f3c5370b68ef2417011d9d40bb2da423620b2a94df9d1489cd4a7a1ea294459dbe3d9d6b6056e59fe9dbe28ca93dfc1db22f33f22b6686d09fa0790f800ab75bf652dabfdd65011aea58de895eeef23ba51d1d593d67cfd188a04fc4dfc2237aa1e1c04c1bf172390fe191c8e5116b801f70ca5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h477e383b12798de1b7e1b3909acfe2b0ee94aff031582e0c5be7a181546906db0e22fa7395bbfdfc3d25f93496c00ea01bdf99cf19e71b988a85561f549397a7617063c6e72b655f1b29a098d4a44b08628c391f18044af96dbf8ad432cf8592a285c120cdf82da74ce3b0db6343569315075d84caa2efce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd099b17d40ac85b089b6aebb0ce4323ae96aebba62c50175053325a3e1eaa0ebdcedafe67b4a1978f58d7dc39c85ac1e49ebb693dcbdabd4f198f962670bfb7fae0dce7d4e6a111a1e4b55eac63c10b36f077ec94444181a63540567a4d12036cad524290dbc149623fa8539c7ca0b096531ecdae5ba9c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fe039d5a99fd93aa56fd91163512361a9acb5bd28691b8a76a30fd480a7f7cb087eb3c92d7c7ca481e65d8a96a569939d41d38ab8818afb754f9f97473f6ba01cba5da12fc22117339ec92830c04ef8f66ffbfb65ea3c7cd405f824a7746bd2f67e64d56927847ee2cea9b946eab16d3508edd64b7d5c50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbad89f72125229a8ca9cd66bc0a23d6d39fcebbe05047165c07ba16dc92edae27f4b34cda6ecc357b770d846944d949d0606fc8760a6e12537424e8414d0cb42b03f52b4220a8e5baf9e9bfdc0989a1c216bda6235088c93311f02ff684469551a2b423f80f2416c34880f93897193af775031a121c9886;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebdcee6e83d76e40600e1ca78058eb4382c0aedef8c52cd041964278f2a00593a58ace457169ed3571bde898f9d9ef1e1f34220acf43887defc125e1d64e0035feace9f1d411aa8c95065fe82d30cbda91d42df13c8119d467c750ca26cb510148b835fb3ba964ac1303e4c413af391a875231d17b9caa23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70111f03bb09fb90b3edb11c7d12e8e12be94e251aa5418f15b21435b94264b6013ce381eb9dda37367e8b45e72ecb4b1232cd41be86f25c3f548849e4d7eaba85dd9236999ff56d295af809d69234c2b895884e6f09ed18a96330959e00e2c65dfd54e91d1b24682abdea876a5c7ba59e0176a14510c0d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e3602dd4f80c9a64ed1eb6d788e8ec8fcc4be5e60dce9d64482af98cace64298f05a60a673665db5ef608f89a0fa9d0e845a303a6a54c68f760c18285886096c5d7567fcf4020b8e2e02663c0852f856eecc0ea1c0edc439195fb0617e201acc92c15199903531812f0c6fe72b183657706cc41ba0cc96c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc895d04a690d2c1b5d9d0fd3f7af8bc76769af6d55fcfcc8d4dc83e3753ec25c02ee6b54b7e09b77ebe3be13a7597ef2756551098c9cc5f116efb790005e7da61704e77d27ccd50a5884611367fe793e2aa09a771392780a5f0aec97b1c29c04fdc1d9b386415887e10359c77b02b32fec709344db5672bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9374ae1113063a4e520ecdf51e00f5ae07eee6cf1dc0ac392a4b9b73690cfb6ebdb89baab584a231cafee97e0ddb57c3ac0aff93f8d9a7de9aea2ad0670d6daa50f56cea600a0ef2c8571409b3075c3fd66c80ab6a650e8381f59c86ed63736c16f0728a02b18215bfbf925858266b0dafb4ebb8522e27e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32221fcde115f336afad540fe49d1b4ff09212e5dc292e097dff146cba399b4424bd5a48e5522be6dab0dd2a21a20c719152ff3ff44c4b4029713a64157400c4ce268f3af58e5b7384af0003683cb349586270766ee94fb00b1797113e1d6f2fa23bbf7751b4e3c04edf7216b8ae63561ab879f5df9be51d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbeeaed48bbee09071b927fde0ecd57ebbee7f2e8f40500572388924e46301d34feb80f1127679de0b0d355c63c8ce13ef3a909ae3c7a2750909a6ad4312e934eb023206dc597d4cba14e65ecdb3423e156e34d08b8ce4d097c4395c3fb5d67942adb8de3db011187ceacccbf95fc1d5fce0fd6e2739da5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h604d67ed0a850f7e4d111a6b94e0d8227a621fdef719a42ae6c8d9c32bde859a81e9b6d00108192b70d42ee50d3a381143ceb2ad3cf265182f4a44fa1c8d74aeabc1cef7d0197084fcd0809102b34822924da038442148d3d9b6bef0dd973c98f8e85526a44910376fddd7d3d09e4428fff03e76e7e41d53;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa49b29c10040717a96ba8ffb7330c7188fe00830995e933800d094441c5d9adf6a0ef505092edc541c11870b8dc755c4557f75404082545267709398faa265d299f6f4662c87ce78fbe4afc9560c2c722565cb0d02e1eb54809833c77f7bb758353da8b3a9e7f2304b34e060b9e52e9740036b1eaac8854;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99a6ce86db0a1f4f10adb8fddbd1b1578dabd3f0d77dda54098fb98ffb9c8d86a36a6e827402f832ef411f7c1b45daa850b4983b5b7e7e7dbd08ce6eaba27e1d9acd44085f0e60b17da849750bbd6ed2b44dfaddfc543269aa83252f7d31ce32113fdf546ed7755c83d8510617eaa5a21a6638f61f2e1387;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18069f1c4692c1236d1c6ab4070b5255eeafa3bcdad2d80a3f353eababf940a84063b6bebf1e6d7fee07b9a1ff75ab6f555b1109845c94bc4760f1573f5e1260d9a919d3279741ebc258f57c7e686a35707c67adce7fa3d6220778e2e1bf023e8a229fc88fd7a0a7576ab56d436ed79fd6d7d8346d9ac5203;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6748eea1d2395166c813d423b6239eabf84401640c36bf9a341c6877ed9a985f5593cf3cbc4024bd59670664984801c8d960cd96bcbd5b7f24facde6dde7ee01419f4cc1c6d0f130011262fd4b5e2b69cf97c593d74a3207f1863bed7b630b79bcb4af6cd29730c559f95433d49bdfb5cb512c42309466e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8c5aa77b92d364d020e273ade018cebea832cfa8506506d37dc2e099792c98d6735686ae57022e39203fb8d7352720fdc5bb4a06216181e9e288a942f6b44e6f02b9f10103d361d86248402c697450bd8e05e0653a8ff4973b0df0c2ceba18d31f84fc29b9a29503d2100b946d65625b43da0ca07c61fc9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3358e951c713a42af03f401be91e3f0b59760c3e9cae0a7873433457dc9efa8531a4712114ef47107c550437ee3a37b5bb091ef13eb9462fb8e2c030d2774c9a175e1e9d58455c80e9f4c2e258a1801cb71719ce3e240f413bb122f951873331b8d8507e86be3470089fb2a35a8191179b3cdf0cb0bbdd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he05ea97dd4866e087d80abd2cb55bdbc81392e6c6a31ab7e396cc70f43b99d6377964d5b83c7f1e2661b9a34b91f2781fce9c521c3e84c815c6b0baf25e09a522d85fe0f0451fbddc87f324845d12773037ca35ca4269044ae0c84beb7c3860163ff6a7c369e9029c397304cc1004b35458880084e89ed8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2fa23544d6da61c4f5c23d120b73c439be7c0a02f999e03a380df4d2d1dd0b8f684751df528baeb40bb9af64457508f4cd732cef8950084c1d6d4a87b6d1c00de5057c257cf9bef3e968787103e9857aa4a966407b40ce65df4a04fb7ce4eb27ec735bf4cfcf6db86184b8cf1f9257145543776051a5d30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157a07be38f58f4677c6c254ebd158dc53a36b492c841b076d8a03ce95c35daf0ae81cf76b447a90cea4add2541a5c03188c66dbdd5ece8b78f75a8d9a6cc9e8f5463b3198c261a7086f0d2e7b771d924cbf9d4ea5b11d059789273e55ddfc8fce9d0f08d990bf946f950b5d41f29e32439e2b2ba1f7b0c7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b912c2b1435b487753be19f5d9dc5665c46dc8015a1e80f750ffbe23e6add9c810e97a0c06f0c6afd65c1d156e377e9cb0b5beae2c422e5d63ef91ce50f35c5d53e959239345f3d657ae8fbfda0341a6852c22b541923fd613c0433d5b354accbe08aa275058e6159d2b4403642bc706c6cfa6bba5fa6d8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b78b545d37c07faff582bc19af56e18843f308d5c1dce4017b7f5ae9a08b184d5aa3f8b881880020abbc2797a4c4bd5bb9eed8d43acfde75b23bca6782ce272c03cd5bbcead4a33d54d86a10fe163b9feaf9a70394abe8c1690af70d854b41d5a9875870eeaf4a14cc569f4a93f6bc2d5651ccffa3d41215;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c2331fa30d751f6f54b7499d642ce3c3e1d2859765bbdeea4420a93a91378385df599d747bfb2a3013460e0807a15f5cfeed2ed51286d19eefc2e2aef67f7f56e3320dab8a04f6289260799ee7639c0f6cd70b66bce95d6fef00348a4362a0463de86e29bbfc75a2866a3aa8a8f427f4bcffc9d81c4e5eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86e158c34d153f64961fd1a0978bdd01f35cc269d3097751f4487ff5d71c8975f52b4e25e3a439d215c424847d4a7c4a24cb52c8de98042a240d3e7d32c0ff18f2e6e86bde4624d9c72e938e3f6ef9d078f6db8f11870b21b2511e3b1b7acbf3746e51058c7c82add2a4e557a44a1b3d7ea4efb6b268641b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8c18ad967ebe93c39d765d45a67361db10cd04980fd88229708b1190ff66ef5db62ac362fc4d06049dbb09eed2bff64a4283384914c07764feb0833b690044f978d4be57e9633331ac9448a42344cbcc0b00484a3fc65e0a78dbc52bf2ad352289a7555837a4d98190619038cc6f5c2a0f6948491422897;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149c91fa9ec23b5aecd620fe74f16f3552fb82b939f6d55c47ad5a068c9b66bb714bdd266ca66e50f9639c3b6be8ee073e7fc3324ab05daeed1c17220465b06d4fb8a87da5c9aa73f60ebbd67fc3d558bba4c1273f80dd8907e5faaae5f2c2f93761e2ff404af961b8322e6c54ad16f70cc67b1aef363f09a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2443eec7d5557f965df7e49c0b2b31e15173897f6e9633287fb82ffceda17f2ec113860f26f221a2e53e5950584e52b402d35d10aa1a97bf7e0a4f36597f75b607f2fd6993f0b027a42ec537abdcdcafd978782814a9923ce16f9c20536c93abb50268a9c50e8c222cf051d2aa1b52c9485775223348b0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181568217f21598f1c90efa0b6241198a21435a5848ade8dd3c72d05e2285ea8517e163f04776fea262099f69196ebb7cbd1c5d0c8c901eeb4e2e9d9b2b4232ba6f8a45790a27861458248053dd69bd8bc16892eb59cff574de37788c076fae0fb7aff73b818cb279c2f8ab288742189da611fffffb6c19d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6b6c42c09b6be436afed2822deab8f33c7a221b02068a8e46fc6b6f3b5a4bda28a288556eb5d40d6a19f1388729eaefa19842cae856bd1a7b7af687197f4f98cb2f3f25a64813867bc77531d5de08ce0d694b89283f52e2902138b89f89b3f54a48c4b8b1e4ffd545230adffe41a0d3dc04218fa6ecf1b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4d6abd47dc7a390a0fe3f4b5aa9f5e6b67958a099021d095f1b9e8e8bf9e53a622fa69f4d6bdce46dd2e5739465ec84b6517bf2c9ab3db289173dca6566797215b2dc529b98d3560a63582f762ea2a5d0f0f7d5d775ea76e4ead623c72aa33c07ce2ee25cb7fc2691e3786fa18fcffbd6f87b8c067419b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199917d7e0d3beb2b928aa58ef5459867a9686274ef5ff0a1095fadbbb050a28bceb5fd2df53057801214b162e8c24eed281f1ae160647f572e638fdd6983dfbbcc3079aa9f31ff51ea661fea29cd603c30f91ebb7225ced3b01aa12f6d677593c6d00fe7c2c3a9a573ab0ca2dc935a6f786464d412456cae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae40a7b433f61277f6c5d934cab67eaaf5401d3a7d01e5aed74416868f8967c1917a392c68184e45a8d38c8d82d2783822d4133e343fb48f096dae8873102386a9d4b3408f0453633f743ebaa972bc56c32507f4655cdf362b7697553c21bbc8f4d1b7574152b65c91edbbe5e1438c78b63d52e9e50870fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb92c4860502611231db7221efd40d291128f970b2e69816b0e965a7751ec716e2e2c9e50927b67ce66d0d8e360188792c75b37ee12a559d1596446ca9a6339e197284c4f813eb034fb2693ebb122aca862c71f4a4d490ebd1d111629625d6b04dc838f5d7c4f7c0cbab06e5cc65de5fb5aaece439c0cc141;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148827cb94cd5a90d769cd5f96cabe6f79679b979150f6ac5c9a33f27260fbc624b52fee8e967a03ecdc7a241f4ba8ef74f349c3b4db38e5526af260cb4d3888bbce432236f3a071304147cf76082c74b8117897eb686c7e26db74a06c24d4e7dddbb9b55589e051327e20337cf5e04cb010c5c1465f6db65;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1270b5bab6b316d7f04586d387ca3a5968c871700fc874c38ae4a5e7f0252493f2c5a1f8b267be2f6c7f9c08167bcb455621dcd2203dd91531e03c320c182598467840c0f2c54078b341a7dd981ffee3a35e951aef50c77369ed7cdcacfea2aa999f72e6c9bcb98ff0a801ba7b305346972f77de7720f9211;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f217bb0fd2e78b0fe0136132032eb0a217738263ebcf0e8094ec8531192e5ef3324bec61d588d5b2f2b51265ce15fa1c412533b012e73e3abd874800f7329689a0d02a5ff69401a87a7a0bf109d9a2b356e9f642d1132a6df85369a1c0b086f25dcba1cd26daf126fac26efec250679ebfb76f64d224127;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172e626a0112134aba9cbdb89cc6c9aa652092335d00e2cfe7e4cf538ba67a4b77d911d9875770592e83647d24371ddcde2c6442018f224086294b2e0bc67d8f85f9d6f147a97727b2e80f7dfc5b9285fb2d4c7b51a8bbc11e9c25740f45276283425c006ce8b3d6b707f32fa6fc5a494f9e8c04d53dc3cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h437f809fb86d111ee09878909525d1b2f113bf7a3158e7be8aa33fba9095026a2f34a30d228016c055d7b9c81f96e63856a011b0fa4ce2288fa6d9c3227d2cbf0d29c151cb932605061acca8f8a4367513809479ec706354f7261a905483f107fef75ec6ec8a89bf27d4bed57890d190b41b2bbadd30d6e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d452b23cfd92be36ceab0cb5d73d4c8ccc66a12ef2e3fca1b103256ca47c738a770bfb9e6edca1734a8dcc3bdd918917e02d797e94f2777f80fa1f36c79707f54f61daacca9e32b0f22c9994334544da0eb0a4d98af037936486f9b85618e431e6848ab0d7ac2eaaf2bb69802c8035f36e0be26f75956e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6abf46e6ded9466f7ab767f2077b2beaa8bbe2f4aeeb7fb6687f81ea8028aecd0f7b678c720420557dd61dd0d46cac510e2a87c57e701116c6133492ae21a01ae7e372c754b065423685dcba34192ca14723b00df750b586a457cbb009cb03984e73c6a643faad6f8871fca0dd3e27503f0aa60a86e0fc4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77bf189f0d3a4d6b118e7671d0a7af0bdd0920b0f5e5a7aa0947d795778e72662c0a2c6e83eb0ad6137d6161d49301ecf715a31a39c59610e12412f157fb20cb38250dc19b30053def70207a2bb78c9063605b54bb6daa13daddf6d414ae9bb74ceeea96b81e07aeceff3a595a60bb678d4afde829d8e7d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1035647d00af437d9650454bf58b3df80f0d4f26c106bd5618794bd5d0d0b88a74a55cd564430d1a975a97082ff4c690c562e3224ce70869f2d445c41b5ca4e3249dec9b635a67cb152863890216437772f8c1cccfe5e284e9e929a2577d9b8266039d33a3cc5c060b4d9a5aee14f797a07ae454cbfef1ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa8d14db99a9c2698db2371308446d46360e675d49b2c59550c50ce489083a773823a17e1220da28be86a6d3d0f5fbda7550cd53a5ef95b635ff2c6be4d0e49495b555282f11b78ee2966f9494d12e3fd6f000e7e1e4e6aba5904df25cbf24fa07f8040f63cf6df611dc4ce06b51119f613b639ed9116611;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181b49c7992de7d0702b9535398402997d4f312c8b32e2849aca8fee731eb8700ea214be9136646565320c24aaba8517d7d36d026a58eb45634d234636d844c2ad8efcb3eeea4e6d7c6dd0b2ea28c318c55c7d2403b026324290384d6f655a091108423ee2e9cd91804e1111968f0c4a02a0b962ac7c97ec5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc06164520145100b26b5ec3dddbdac4f2ecdc0eb4a3964032c7ff09e9ae5004248827f4c1023e65690200c6718735b928b6ed9fa215908ff8337ef4c4c9b43a93abc83d5f3e8ad97142c1ac28883d8acc7b1c4930cf1942ef6e5382f043318c3d33ab82ee35460c68d774eb6447e29000b86ad549e9829a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6668ce8129a6fbc9e6df9ff27f2d031d0e6252849ac6245b7bdeca5b62705b59ad8d18b118ac6ff825091523d57e33cd1013dc598f88e78f3f923a6cbf9d2d0a22e7b53651376d046c18e11e0184167131e8a6e4a5b42ac7d1b8773f55b126e3c7c4427f49596332c91aab87ee5547d3dae10dde9eba6bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e51057fb7deae593046aa1a12f7085d75abf654dabb5d23c3c17487f0918f4097294acfcffa1c4e9bea054568af4f81f0df8fa57c44dd55977df76344fc87a0ff3f6f15c04e8273645d07b81b1a4738c85ff98feccbed480cb700b72c679dbeda00e4a7963fc2df64484d6c807f4ce1cc1848e682840da5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8740713b928bb2a8a49f967d087aeba68e8a6437bddb1c3fd31b2290c749ba0ed3827f7a0dfb05d8596dc0244d6f4c2ed23c3278410197adbe76dee4f7aa14806859a3f283751e8d1c9aecf244dd16bb478f91e6cc1e3d58b6450eb4bb505e42f5b6451ecea82a76aff4b0cb936e698e369a813b6452db6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1057ca5a0cf85bd5efc0229eb5036ff90f96819daeffb210233111d5fe392ded101e7dbf23f613ac6f384a16f43b19fe397810cd9c292be14d9e21e366255c31aba6fe3279a4fce919d84cdaa92befce62f564c620c75be414f1c42cc1f968b3a0321b8b96fa5acb13fc16674ba90b207ab923d0ff3958c11;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ae446d4db2e2d638688ce8e41427ba9fe57ecb72e81e2bc3c9688cd80a208f6cdb2dc00133f5b3ebb21d3cef6ce6e30945d958e30f050838b7dd43428541654a1b82bd1bdc3be4cfdf28460e7013fc5c238857e052998d6a933fb4dcac7591a365e199e7b5ca5dbcc2ea7959eb8bcb1237e6911e8893c8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6eabe0ce66f05283ae428517132a2b1a928209a9882166f64a910d8e3625497269c984a313948307480376cd72c22b0cedfa0fc1cdbbb5705b1a9d0a8aacfa9e234476aed1b775bb5c37e24064c483bddbcb1af96c8e4bccb9f66ed0c5218176fd963084a702f99b713e0c3a97693e0ea956c9f0d1313aad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h332e2d8dfb2dac671543569856218b8dee77b747df448da05dd9a0a2d83c4dabbe672883b7901cf0922dc65a1641e815460cb446e1881725fdd0e3aaa2902a20cf4d211f75cbbf7a76416e844a28b08d503f9e4cb74c00b446de26e1764479254a87bdc84e554f2199bcfd42d915c8da70ed28ff9dde7e26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c860887a693d1367f4c3f533b6f7173dc3cff07f84c1d586a804b17b33bd59d82b63575a9f67a7e7fb08754e51ae7b59c10e97018c4c8ef1db228aecba8b6f9a37dc40147659efe922a68e78c462babf9119feacf8abf054da8f1adef7ecd81aa85f8533c1288819edc9d02504e968a472f7790a4ccad69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haeee0bc7b25ea895cd0e7019d4612408e70108836a3eadecc0d9f52301459a4fc3deeb211c29b4310850714fabe449d72360e255352ee5e2d2685aa9d82527656c39f8743ee0aa484e628cbc753a927704370e443f40e3fa80df02b101587aa4b8949437d9a19a204ebf274d54ba716dd94b1ea5a582976b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha94419259e990bc55045a8e3a50199aeb6b3aaf54eae3e2cee87bb8a64ac38aa4c771149274c0caceeb35b8c185439a8272faea8b58a5829831fad014928a7aadafbaf5f21683ec404df91572f355bdf1f596e011d9d1506bde55364aa8b7dc4eb75ec06dab587bba5536f8d549926a92a56ff7239319cc7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c251ab24c3db4ec512de7ce7097f2764883e4bcf13d76bdd11ab5dd626fdf1b440b254733ffb979244c9f3713700d1e23f15782faf69d21762d3bf072620f88fde5540fcfc16ab84f8692b19794aaa490bc3a9183300317c9cf74d3932eb3985437cf259e937a27140c30b84bd0fcb0e0484d3feb77169f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae43495a3e69ae173efc73f8ed50aca24319ad2ec710b057ca01d2aaba1e51f67dba7ac46d5c781c107c3e8ef4c5473dd1b3a7afea510fcc6920cdf2f484e01193bc718d069154604d8fc83114e2d87e4205260c4086ccc5c6bf6b95c0d4706e8a12feb7ec5e045e3c248185653250219bb120f77e821f2c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b1a0dd3964da0ee5f9893fd6ed0cab69747f360e5fc45e22f5b286cef6d0ae32160e3f6c8c1483772379f05c0c55820738bf31dd9f788e644814c7d717c2ef64541d8d37740d985a046beb9248ea7cad804b88d31112bf878780465803b950afa3f97101c3e31dc85ac15b55cf2af86dcd1ee7a7c04f08f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9a1468c4689992ae4ee04c2a029e2b3062acd52510d76f6117e490b9748143f29f6606f494787b46589a4432e3e04ec548d15f5dc96c80c2942fd7076566c9dba439875340a81c48d25339c0d48710962a4e38ed338661f80773aec88e84127725eac155de05ff6916c9ab5ee3b01bf24e4da6f1a1abde4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1995f55b481f45a7f262c33c256127a15a1d6851dc54b8f47a58f485341586659ca25159e304a7b8f206b7dfcfb0218bc8fbec9484301d90453ea3a536b94f78a04f168e3971970d0d355ca56c22e81c5c210c3752be2d9f48967819688199e7f579436d31e9ad3ca9ae63b0d7af6af760c48aeddfec32f54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac5f726e1116088d6259c1e311c423757e4676960f6e05c31fb9bcb4a329de285f5bba5a51650bc9a53dd94dd798dde493c63f91e8aeadc677bbc1ffca73537a73c22b736c9a31c7a3071f6d8a5fde443b7ff6dc5d704e66c19adffbfc247d2effb996a2cec9412451f34cb83b4a67be69b88e48998e0df5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c98c8bfbf969ba196e083327693b0ec61f864fae3fe821f403a028ccf9b598634ef8e44aeb82d03e3a6c7bb91493b58d61a1b1a6751a780b6bd5efb32e01e8d89f661ac87bb47d3c6b746a74d66cd2c22296721c5f5a545461b2ee8c1f36dd4fe73d0340ee69d86045352312e8e2a9884672f939412ddb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22e61fc3b86ca286af8723f3ff0e96807f5c963314b37419f2f0291bb11794bc6953519eadcb91c3be649bbd3fd2322717adc017744f1e95b41a457e24ef71233a806cd3ee796a0b964bb3d100ac39c87dc09fa443fa55be8bed62048f63bb401d33236ed07ffaaa7faf6a7f75ed5c34c243d82f3e2b430c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ab58bb80776d88139fd80e5cecae8322ef2de88720c858f927ae5dcda8692a825823938cd2e32d175be14450a3a4253a34f8128be5d8c359561f7dd0da02acdf8eef77161b4ccc95c4844a69889a90f7a15e4ae2c49144197b7a87daf030ea67b73ae9be01641ed4fa74a848acdda49752bb15a915ef3e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45c91c261a2f1683774fbd6d3bfd896e37a76ef6cadf3507193ae088f8f36b68e9f5ad0acfd378a23d6a6cf5cc72abe8c91b888447c8a150cdfd26f8a1d4f691fc8096ee647ab4cd7eecfc741e121bf46235297592cf7753fbaa9eee5c263a73c6d42a285915c5cf11e7f5f787bbd7e0ec2dd2915daeeab1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e99900f239b74fcb52da3544e30cc95788c57557ea29ca1e381c5e0db48f2264d5ca828d5b7acdc59045a81242367f9dffc1cc5eb3f815209990c2082bd614cd049ac5f80530e9566973d29f84d4faf9b05210ced2d068f9f3d49566e2076133c9c4a478ab08d1840614f66f06c71a1b566a618801752b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3d99bbb4d1202861cd24b743bf1cad48d87c814795d78d09a8120d2fec37bcaeb120abe81f8b634948d4b75fbebce1992f74686edcaaacfa28295d310f696e067b7b489ddc8ccbcd5a0130a75e2b69e6b7a4362e12f188a80eec8c7d99d948106ba5773cb29ea7754d0a88a4c1be25e0cb886e06a3273ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb9fe9a4ec038d5e2fb92b8a5a1f65b6e5f255e82baffd5b9909231199b885d7e7769efb96ba653eb547e66c6080d5debdbf03b66d88659cff2ca98a886866555cae2d0dd1f151ef82599168fc20655c79bdbd518eff7a7c25aa78c280813b8e699b0c2e6bac5f2790437507560ca1cbc266f4be65793d79;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ea46db05535f698348f2cf1265eee970cc5e3f8c4ba598e8330bfb31fe053e3192500317b3b0f2368282f8fcadc9ceb93f3c99f3b98374e97c8775b062778ea5683032a017deea7cf69fbefb171e79b5df7c32b4e7f721050b44563913fb96d94556647bc78aa3c7d59c6e2a1b4c0b3398ee5a58a13c7ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf60076664b790809fb8b3ed9865503d7a9b414555fac5f0c42a214c43c5d2d16fda8708e9c5b471870837f278ca1ef2a1f3ecd0ade294f68e688f4d9b019b6cec09b37c195d3684f0ca593e938281c42b50502967f70e841d1b7f15fe6f9f2739addf04ba0cc13fb94841156200d8ce23fea610c65cb2818;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f197fa27bd48186dba410c7a21c1743fa594f2365ca14760e8b1ef2c7dec34e83d13e29fd3dc16f8169b371b511994a0dddd47a39907359c59c1aabb0a1c45c934ac0079d67f2be93c072b438afe2e51ad156323ad53e9399ae59f86c90f4c5964bcf8e5d4e28616f918445915f42d2877d13e3c2df9e59;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40c599c35dbd2a013efc242c156f8145dba87cf5b00008c1fc68cc3701a3b5a7a991c761af9ebefd07381ad797a1b5c356be95053bfb70fbe7008a1159dcac9f78ba38d1bcd72723823b1b478484cbdb317f2dfe424ccdef57aa68385b0e7a68464f5433f4186b74e78405c282d6d7aea8d49d3385ccb7ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h827e7d08682ac21344e57bf7c5f43b49af09d0393c5ba6ee836b23e99e3e99932d9fc376cf8c010d5ea85beaa0a625417376fcf65d8a01e7932943f68b3c4efda7ade3f90ee425ab3c17387ce96fe50c58802d6bc806de979dc4ab63554935d35758f1fc3fc9685ac78d2620137640245548c6680d7a9dd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1464336f20d310e73ad952f7954d4c23c22bd6145225c3a2e2a429d6a4380fb823db436fd2f3ff9fe46118395602ad284410c76b43d64761ce33428c9f182232472c529cc33a6119fe2e1cc95f92ebad67c08c822fae04b7090650a990523e76517ec8b156e26c39f29fdeecac31d0b760019a193882c022b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3bec66319838392d2c09415b54384b7a9d6d8fbdc388ac08126895100ce5ba119e98cc42ae85edbbab329832ef042130958add09a6da7370d74391a604fc405b5b851c7629ba34d01b838b529b0ebfe6f1abce100b2234ae708633c0ddb42a19efbec0bd79b5cfe718c0f5735cc5bd7067c8e447161cc8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c7f58cc71957e1baca3e61b10b1cfc5da40818d5ad0f3ccbe76a00dbe811a737e0412c679fea1b05dff68e8963eeb5adc2b29464af11972e62c5ab10a2c5963acecf16b6857c956daa4dbeef598fefaaa872da277b620950c616b26bf2e6d08c4d28f13f6c56c39cc2d0c36da309a8212366cffcc6c67cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e7c5ec09216cbb0229b5d562cbb639a6edf704c5463e79f587745405831bb3b999ccaa791d73d43e838e889fe7e7ac78e8437ab387d4d8ba5e6dee77a8939e0ada64d71d94d4e10052d5ad5b5f112b7ae0e655d1765a03cfae4fa65d39c066718d42803e9fcb807a376f2e37863d3e601ab5226a74a7577;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7e342fec1ff38a99eef7b6610b62cc395fc5bd9fce1ab8a59821d31adcca5a7c2abc692007694e4d82c33f7bb8fbdb2471c6a1e21258b50a8c1b757d2b4c05a91b5f6334c8b233369b38e3f8f86f2a8a46883e9cef3421478e31d65ba244367da65d55acf048a9cb6d52ba8011820281bb181ef73184151;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d2c4b660015a0f804df4c48105662b345142dd20c610885b3edc0e95b3b15a394658f10674d6a171dc918ca2e867668e74dc561ca6276c01bb395e92a1c646c052d6fc32f8dc012f34592cd50d291878d1be9b330b8aafdee6697a8070b41ee8a86d7d5266007fe7f34c03862b1d79c62cb8899018b94ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32f538b12eac7f2ec1b4a71a8ae093d99fdbc6b18980245c255f5ebc88bd49d9d3408af962809aca472fcf640c11dddbf4e540cb37cc1225ac3856206dcbfff82766ac75613d1cf98ba34bce9ad6b6d11c01cae9607840133ea932e61ec302ba3e121ec0fdd349bfe2760f9441c85d459fdc33dd6ca481b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181fd45e480780e1a6377a1dd7a37d65f88b2c5dbb3a53925a9a892096729186e1c26e49627fa40af9b3fc1de34acfbf546840086fc7ed738c327c8dbdec616eec2198203e5c83aa85224494ed9cafc41a83da22b3772ac29a8541145898ed960206496531a2bc72b5da0dd206d8cd890669286ddb7f51e78;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31e6e63e21ff29f57edb0ac9eab8f58c0ad7ff56bfdd694794e327e4741c1f6ea5f3ba0f1184ed2deb4e1d9d6f888832c5af36864cf75d630b9846ba4e203d54d34ac0eda467781daf368bfd6b80af0ccd50014e2fe4bef63a8016fc45a224bde4a0e19a450018bad9eada694e666bc6e017ecc97b8c962b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c2ed09f12a7c046815705bad5675101af3a8d649d7c52c55d5809590776757bbd4981530cbec49ceb1d5c436e79a5195b5e074ccc2efbb32e16b98d2c245c49a42ee83cfcda3aa8ede39621f3e193913b90a9b5383904ccf2ff4e31df82b5435642a2f1620588de15b2c82feec9c2a9b99e4709780d372;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7413666dce785b32571e556b4337b892dd3c18072b9d04bec91f12e0b558ec36cd9474b807f46026da3d876a8fa5be64235807549b7165d259fc9b1660f4f2faf68ee4f9a58ed7d3d7b6b212590b239504cab1da425ef67426190566747d68845a0d9ea9c09249293e4ce2ace7606df47082a3ec2f7cc883;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa21c44b17ce41bf75406791844467affa445d8e629034e61ff53fbf8bb7784c25d62c03fa9eaa62db036843049f3a5932636cfb1f29849648280d0e5e428603bfadd52d7728bbfa06bba9fbe7467ed5ed05928f4e340c9bd258dee4a98ffb5e470d68064dd62876806f8a06f0d33b119ba163dd2a9ec961;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c45f27e48f0f6668077d7a29b1ab7f945fc816d0c1b77d130388385778d90c8097dc725ac053b241cb0b0aa048b48dcfe8980a8ced8f82b92f15ac68e8ebb5daf8a034c01c0e77cfd90d7e3b72a0c315c67b29b3be3937b092830927c40a9e7850990ee8f3b9a25c75118369ea49c25a7175fe987027fd7a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h577939954d9803a1d0a36139c1eac533b71d0cc78b52393dc2c50e8d1c0d0a6e355e5ef89474ec5254c12c7d1e351e66154f62ed55d20a09f4e68e48f54e5342f328374cccd5ef706ecd177dcb156660a1e44fe006719ee5f8f035178b17cf5cd65d0d8a0189d44baf7f0fadea0d8ef573099e77a0347ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee8f55ba685e805b74ef39700ef8a201a98ead807504dd8714f2e3c52f9a6d86abcafb0f959a863b1fde39d992cf56334ed5294f1de4f39fe39986929f800626910167da9f29b5d7e5ad784c24c90857ca9cb11270e44570a6a19fd88e054ed402487b509ce88aa3a09c9bfa92ca9331e419f59277f4060;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17479a3edda458bb0d6babc2da383a6deb8485dc9d2a9a19de0e5fe40dd8c96899adcfbb302a129499a697f3a0bb47f64cb58597303dcbbb243cf5e26a6a54e987dbc65aad804f5c64f79d0db49b11643923b22a972f8644eb0677916c5738fb3b624c02719bc3bb3cadcc9ed1c0396ee49ebfac34cb001a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a4b74e1ed93817933a662948de18658ee11ecfbd54f06dd418db310adfbbe90b27bab2d91c57445a60b2f6edcec8a73ff75076ad4a5dfc29e7124cb094b110bae3205eaae56474dd101a97a2b56d3fc9a272a8ca296a64cfcc8526b51ef6b6ae7b5f011da6bef9c5a9378cf0114a2515699ccdb753eb905;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1218b82428501897a65e03676c2b6cadc90a1b7961bbd25491483ae69306a36d54eff877bcd5cdaa63c04c8f6eb5fe0d0cb3be572f8a0f4f6d155d91d9cf9818d235c9f78b45630449e47c15f568435aa4dce75c5cd0195c850c6e30f43a1ec4898d9bb259ed053a8fcd91b649c57b8483ecc3e41cceb7295;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb891d4cc4d496f7e0ce5a4f02958814935440ff7007766945fd36624001e4a4a7c64635a9de6f51b7329d9dad52cc286691a219ae94f6c1a85e04b1e9fb691323741d4f2ec0c86c2aed02751d448bc56fd4e194504f26f6144f3acdf21063a510799bb4132b6d8864a3115997a43585b1e95b4687075890;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa643fcd8a4c1706524a797ca05676a96ed5e4e608b6c1fec04f38d8eee78f4ee16fea8c4d1f2e7548f170e6f11756b1c8745a1fdcf47943dbbd5b4e23c7c14dce6c1abc5c9e348d76b78009e31a53288e30a2912452126a3f68c7c42a9b522d81f443af3620b4ddac409a3a5477dece2791f7726c87af4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h164d0baccfa05e539c79ad51b02180fadcb4690394ea0c1e07eda959c25f55dd43c3e24ab97c7fb687f97ab6dee21745605487633e13bd17e7d19ce2307836024f09a31c3d9786f74a068fbe4e760e73609af65cd7d3c4ae993362ace1bb685d71eb4c6230a730716c1bfdb905add0fcaf201d6b3cf84c5c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1391188c90ba4204f905d5b6250039f6af9e3502bfa54b7c74ffcdfc372814ae5c4a2809ea1f88e0df18297cc720b4a9ffc56865a0db9d33fa39bcb5c5dd271be763333d93263e84809f36a9d2b2cf3360d05d09a77788e22dfc3c20c6b3efbd7ca803e8e5a7babc69aa1e4e98d20bcef19e1a0b41c1de846;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c673f20ada832494455c8c011cb7a04568327c5d9a633847bc543e093672dc60cae3c7d77034bd269720c3c83f2ac63c03bad2b9c52fc7bce98bd947f0a44a598c24d38abab7c219b903e4adb597d03fa9dd98026047c9bc77fe67bf3d0a458ae26463f1cabd2259b368a5a3b939b2e1ccedc08deab63a65;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1144760f51fd78ba57a761340fb42f052db02aa3991b37d845a5dbad6ed9fef57b01e35f132f3882956ef9753634f9b58019e86a74b0085e44358f723c1e8ef8d4981641ec5ed06995bde35eca574e14734deaf19bd6870d288a94e32ac1e7ae0189356001ef43ec3538117ce92e9d4af6c7e048558047834;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1800b897f061ae2bf6c5815e44f8ae1ba2dc36b4075fecd253d1b801794589e63992178cef9a3c56b6f1b446ea861f43026c7a4bbc7d0c509559dcd449e0f52fbb51c6a687d0cae440983756fdaeecfa5cfcb53a9ae306f6c8487f470ccc262d04c08028e7c86a6a9cf287944f14a613dc2e8c980d5be8df1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha616b68befa933d1a3f104400aba72457ff919359dd0f6eea6373fdee97db52029bf40cc4b8229b26fc63bdfd79c5852bb5979794faaa8a6f39a1b51004d652ee83713375479eac9dfc92d51b891d405ed0e74cc1812021def19a5cc75c5edd44471a95a6eb0316d72372a5ee06487d7c0509a121327e3f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa0c4cb716e2f678fe9c1acb8a15441bdfa9bb1e94fb640481311b7e0e2895eea246d166ef106930edb3eefdae1129560f718b190839df27c8c13d0fd825c57662bff18dd93e454ddc45f218e5f5f7ea930e722aa71a8e47d5a70bea8c8140a0a0eee349dc54a5fcf1d5ffa9672bbc82d2103f0351ad1d61;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c08a0543241d22aec39bfadad2e317c21170bbcf680956d2b0ac660c6708df5150199b4d26a54ccd43ef7ecb64ecf2ea257ee3d3cf7c32d66fdadfaa09126229a5cb08580bef951183523decbf9a4e91fe7db5ccd93b36e6ebea38056a37f75ed4cef3e8d137c8d12ec16b0af11a2301fdb10e233d0605e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h343db7cec6134175ca157fb81bed6b35a4e326b47e7822eb9ee193d66dc68df41c64e356b47d0794dc6d9414802c01b9742bee30dda7cac376a43f57edad62ad658fc39ce83e78d1a06b396196b228fdf3b2ab42d8a7e4df7975a97104b744b58612c1441f0983238972767c6041fc95ecc98a6b888eb8c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf33f9bf6e3d60242cf6bc9efaecfcb2e63a9d69ebeee900d92037d4a7671eafa33f3f3be941f6674b64d3bf4f32566204480e135cc0a3cb2731c1c19eed63e9785e740a9d06529a4952311c91878ab64d24366b390539a47156d5fc584c62720d27292b62a9ecbd4e3f44bb6694bec3b457e0c7f39c15f3c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab3ba7d9017ac2ed60ebb895a33dfaa685e45c832d6706816066991b4353919da3156f183337b53ed7b00eb8e2983eabc4a5202aa4db000f7177055e465f94922055623aaf516a55141d46e37b18759c1799f85ea931145bd975c6a5deeb94708eeb9030473e6ffc586da18c4bc156c4eecfa4c573e5a3ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13901cb1f3190ebe765ebba1b269dff1309968848731026d8655164eaa21c52a767abaff03b66391aa9434f7e9e407e43da9529d367d25ccbb1ea8d10be064423ffa2f1638098afc322a1b35c91685faaa1237662e928b3a4a5cc3e1ee66cf760fe1a9ec29872a9921d01325fa0abdc2e6a2c832541118c97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a155290b803ad734741f2d081412f86812a0c32bb6fdca4e55c921335e28e73c9386f3ebe5ce550cffad88f9b27f718ee6cea5408bed92c0f0b3e3f93fec9ea92cb6690b2628b191083cc151cfbc23f920e742e69bd1d92b5600fb32ca1914adb45eba3771dbdcbd305943a66778d23cc6dc206bff48478a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc85ca13459a6aaff0fc7e0f8876eaa72e4423413b12a846710e224836f5ce0c24f3d1ce5d925dd55d40002a11e0ac4b7a64dfa28eb5ead979c9314aabe1993bbd372bb8ccaaf75a0e2d92286f04e3bdce6ab4fd02ffde707eacd5cbd27dad48a96927331048ae2303bb82d18efd5de778421cef1d09c32c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10054aeeacc4dd68c69ec9ca223986b4ba6a7d19fb82267d7873d6460b636c3522d2281e3685e08621d6d1f6261f09905353385172d11671bd7f79932f9ffcad1e89588d1c15351439b34988ef55cf18b85ac8106943d0bf3cca07a2081f91276fc77cb099900865bc7e0d66d07128d1ee40a41aec17a6cdc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f99024771b71356fa6319567e51ca1ba8248a460abfc73ff67fb12e06e0af485dff892b18e3bdf2a3a73fa16308b42f1f5d59ed40cc73d036e9a5c08b24c9325c8ef2320777908e4863aeb5214b600f94787353fe56c15e9e0ffe6403acd6c8746910ef2124bc748990fe4d18f32712933c21a793b3ca85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebe67f6210431b2fe5392a7507822e7f00bcce73d4b42657453a43a5972566f219c71356812a6ce49cc2a0f5ea00ed758fefeb48812ee3e4a37123b334fc07201c63e7578b4865989f2e4d608c60a50737dbe9291e60472c199f14bdc81c1d010ec32af77ca73650a2866e6f2ec07510469aafb9fb465ee2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9f89d515f3813b935eb76d7f65258d91742c5221ecbd358c6e153b3f1378e1c3d3ce5ce8e6bc0ca07773a8db2517081f8d24f6d92795323ceb6564fccbc35260200c1dfcb6613ecf268e26068c244841978567922cbb0934fbb0c5ebbfff80e58489ba9a7fa56519ec568820ca9d26c286bab7492213a4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c5dae7a82883cba4849afd724bef831c87071537d534b420e9fdf3644364269342492cd5e02dab70483c81a7f190516acacd1f503582ed821e00e2432a8695076f07ae637852b32b0451d25d229e9bdb235483577812e41cba09cbe247f55b5348894ff5108a48e82abcadab69a8aeff4cf9cc742b91c3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf472f9c840ebb7388113837a50c49cfe427f24f3b814d2b04d648736a32c0839d54b8be02ff4d6c540ad5ab14f289a7253f9c7890431b44535853b72a27e80ed47f4ab81ac5aecba7b82c5f81f5b5098e8ded31c642a1875025caef1c56c5c186f4771b9769bec7f0f8533f4cfb26359f0823d7336a81c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d14a1605e960457e835d9e91f8577ef44534ef280be63e2a95deadf5b9ddb7aa26f457620b44c4c9014ad34f2d14a97b17934f56635de99777a2d28855a2e1a2f00386707d1eef9e0d6e1933e43a41bb0503fb323f9dbcefe8204579b34d97728a886fe2101fe0d5db58168f154391a7527bcc8534605a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd69c57b26dd5f57f18c65638cd8916581c3f4374fb0a9668c1243dbae6c818fe26a3f5e656bb9ca7c9e770d27c95e357828d2e5f003a1094d917fb05f0f119be30a8e8a682c78ebd18bafe9d550a6ac8c56468493c1a56c7c2b642da5b0a1262bbcdff1c215349bd655260bb211981d471b5aab67eca725f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13725638bbd43f2ca0538ab81247496d7251e3fddf2a1120cbb8d1a07af4390b2ae0ace2ec0d228f81402f3bd8c9b2ceabe33960e9563fed7f2a698ce81f9fd22c0a278881474641507532d24f9d3b0f4c82f403104ee373d48b4cc6acf5dbf2360fc5b391612699a7fd14be206a53f6885a5a43c770fecdb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a90b2e2addac0db726bca363bfa9fc14bb2b9bbf6e16c118194a32ac7ecde4b02bd4af327f2398e32b5bcea8ce441cc4f8e3ba5948625a39f6981816c544190d3e0620784b9933c040c9dae79c17fa79e10c9654cb11855273386e6d8e0f5a714daddb041b0d6c0ade98e75bb06d9f9ed46ea0ef85a16fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h431a71054b12806de434cdd24faa42453799675b432b2c6e4a0241b9f2fe23f101b4e60a2180bf9af0fee245adb961d2bf2f8878387fbd105c4edd80568f13eabe7b9cc2161d24b603cdeb2efbb44ee3746a4291341b22b716b4d085dff3c35c57b32786984523ce343575f4a6d75403fdd1a33b9e068c1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42e6324955c0dda250341a4bc9875aa26be854acb39cae50e67edabdaf336e19047a725e5b68f3a41a1d6269de9eefddf5decba642f7eb23a98192fb02d6735f89a406263075ddcac2b354bd9066d49909db56e926eb0855927b4de01553356129e891f4e26ad68b78d0521f6c9f466a5e586ed2b5aa0a51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5ffaa831409b5e8617fd555150a2cbe1301fba71f97332b5002221f03358311e0a445a47fb6d06e2d9d67304246055592ac0835ae84137cf61429fb680cebc7ff27e6f68612993d2d8401fec197c4067cb24366312ea128b9bbdb5b652aa587cefc455af763bcddb63b7236fbf9d5fe15586b93450b384e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50507438c923efe4c57d593865705d90db372c51f091b89d2c313b40a69172ed06a2634a41d43241dcf25c4f58f8d7103cfdec55d53d91f6fb5603494bf04d9d009d1a9aed85aeb8db3c97f6fdcc7f6af6712c394e53ab7c34dd7d040480c2e7d3be31687a1ed319e847426df03fedf7f815a4361e0e99e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc80394ecda8a58cc73561f00df906ffcfe1542f0684b848793c9a3d4f72269ec4e01c4a16bdb9a1570adc04f1e2bef9cf08a3add863be41d5dd7f054d7a55fd7a90bd49cdaa7f720e4f80f0f72db06e0bb9a598973819ae554b15f051511302be6adda79371cb3c63d2185692836fc725fac28ab73826921;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee07a6c8d8402ba11eff291ac01971546702c49e3e81432cd38197a9906a58699ddf03d6472cfb330b37aa003ff034342b914a3f3b4e5b03b01814da6ef9281ca1f6bfc961f21e0c013b7b43771e148edb6fde841609bffbab2a1a7430d6bebec6856c50560f258a9850d5c47c93632db3937915a550ad75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13335237c55235c750601ffeb04bca837f5ac1134821f710a6639b050b12f5d5a0f3457515c72af93762462144f0a2199a76a2ae2a5d0559f56d21e8b688e1d92ef62b3737104f692a5106698d368fe0e0ce264e68c8c0bce38c6b0f4c18f203573aacd0af0ab2e029f78ee83a6ce937bd2abc23b041b4550;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b62b800a3f7ba13ece9dc0d03706174eee7dc11420e556c55c44100f21175c5eedce656ef0eca484949057ad299b6daddc404fa17f324486c8627948d8373c1e9e541c552bcd695a1a114d3a14facaa58f74c8e67392d742b916ece5cb3b52ea568f6f88c54c1a00a5e24df541b344e3684b817cf9b91448;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156950dceea5cb3eb0032f7d6e88b8a92ba2d856d7045611a148a09d53532a4d1e84f4eaf3f2e678f463cac4a762dc07ecc7389b681d5e3093aa925c512e4f420f861f6ca2f363e7bac78799557d3b6c64764afcc864b436d4a3fb2a4a89cc0c97edda13eae39c311e30d4bff903b6fe32828f85bbe9f1237;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h749785a75703a7febd3862f98df7b5e311cbf191f8949a63d772b430eb2b9f3fd85155d0728a9d4baf4155a94c7fb997cd0a71bad3694ac6ff000762161ed2bed17bcfd911c94885d1f8c2d56ab170ab177052c90812b5d760d3698e23778bea34a69c2dbf2cf714801a73ea55183cfb666a2da0d9cf297a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ba1a8027b345c888cc6834a49ffbaa1d49f976380586e0679875a76d9ece81d07d2dbf0db42ec2918b3cc8c1aafee4d888fae82bf4ba5df21da73bf9e06220b77dc4cac28b5c3d6e9272b45851fa00e1307e1417979171bf4e153c2b005e6773af3dd57f438184e3f00c3ed68b90b6626ee91697aef798;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f580b884e7f40c22bb95efad62716849dae8dd4723cd8891e780f15d68e81973477b4d8239233f49ed8283e00b825996c2983f2b5d79c608cfd14b9229f136b7b39d86dd46de89aaf9b4d72e1eb436b02987d79c15ae3e2dce67211f3846b09b40fe1951a34c1486b6be3a50fbac9cbb34722bd0317eb90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f0d4b3635f23e6c1bca87b065073bed19d64a4f0d97adaaf6559d62138330eb5baf62eb096706ce15b8639fd62322f5d8a6e1ac68c644cd1ba71395ad4ddf907d2cb0dd450ee193907d2c88edfcbe1c77834c6ef806ab8c36d71c2a55cbaf28669c7bac4a42a29c7024d87aeab8bf4c94d71292d4e94529;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb311a694bd966b8b1269c124e50633f00c6cec09abceb29375e3af833b4e524b92ad6aadb40df3a9b17325a18221be35fddfbf9cd41990eba64c72e6c33234d5d40f120b43df2deca950ff12af30d453ea974179a35f1cb81ff7606c9e4ae599f7e368637babfd25f58bc29bc45bf2a457433afb4de32b66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12886cf44100f1f1cca10214275147c0d255f5b3f5e157d57067b66f5e42650f587e59da437ba90b4e9a7f729179e02f31e351ad6e072b8287dbada64667ab51c883c42560b94ca7e7b6027d02839628574662a43187e7e96be980bbdbfe20f7eeca043f869ceac1ded494b25166085b9779a06f7575f348b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29694abe298ad011af581c6546b420333a76b07ce20b7a9d03b97326c9464c3b909db9e7146cb6a548892ce34578302aae5818764edac6ebb82291b2784489f92812100c4fc1bf9a6f32a08a3b3c184be6ffba3e0753fff0bc260541f4b2b2fa07f05c6e967405cb60ed5e8409be1cb31487e7dab25e1016;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb0b794e7aba29352031aeb04fea940dc85b09c28b107443887483e942051f86035480ef333effc017e6fd6aa7a46e0fd1f34015075b9e38a6f75bf557fd350d0f6d73b8700e1f84361cdc09f842d3b758f407ecd45cacbb8bbd78fa178a0b84ab968e61ce13f1e57336cd0d5ff6d5c3b70ec0ad0eb22c48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113f6e6edf93d4d290b1f34ded02215ec69c5d664703fb7155610ac6c4743b4b1d9bff2127e49ce31669d3f485228899fdbdc7f9121ba64ea804dacadedf7ef4bb5d2c774afc232500b3194e4aa530af9e48889328c7cc3656095645330899f7b5863ebbeab7a78571e8d276f1dd58b9a3196a161d10b9c81;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha457cc57aee03537f059293005dc73a440675f239286ff4d0fae46b714356eb0dfea171080bd471ebe07e38c50df39fb1ce0598b9274c2e888eb7fc0f94bb2d08be01087de0dca81b2c9bd3b211d0dd498f50dd8e9f58477e3f5af7c40fd14bad373c644a3fc872780fe70a385c5230ed404b8556536d516;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10684826d8e763901a55af1d9f8c3449a1b0c06f7479de650bf65704d4ef23132732716444567d5d608e97ed7581b9251d1f26c81fa997e7c03e6f1029fb8214d06e6a1bd572aa2efd103359919892b93c3d9e42d88fccaeb1efa63b06ae217397ba3826195420fc60b02159f42f2bd86f25f8365e86ecb73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h550709c58a17b1dbf5170f8701ff4e3fb165bacc1ad86715cc2c89fd34b73065e80c28693440675525da3f2c92af0d349b5e8c5d3d00531e215428d3708970fce534c901116324b2f18f05cd38c97a0dfa55173615958d6470c10550b92e10d826736308eb68a9e0c1c8c53c7712afcc1fa7684e10cf9f1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc229e6196286db2af4a1167237fac33d4e73556f87366988dee460572ca988030f95a2c5c5c7ca136352f95ff9b84c6951ae005033fc910a8ad9ac3a84a58d5c07df0db8476fcbac3c1bd12f492a7404595e89b5abda01296196398bc573a18e002796df511b0684558001f3bf05f7d44ca61e0dd1fa9f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e3f83645d8c65262d655add9a5f602d60772fdc2f233cf2c1c01a2acd1520b533154bdbff8f44f75f33b347c4e57933aa1c74a5e7e470fba886d06e630a9795281dee52ed76a14b129e8156742ae8d5aabea2803745358ccceef79ec3d90f314634f4d4375eae223e2a54d65aa384b333628d3c5fe9d10b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25f7d3d51ccb04710784668c8b0bc4581aabd5de2bf41a1711131de2a50acfab81a096e9fd4bebf7f24233e531633307f5a4d4cbaf2ce129ebd3bc9de107cc634b1ebcdcc41d340c833bbff707bd46c5a7ab2f16dc4477162a7d22a18a97ae1c6abd2c571924984bb0b15b71595605377edc11ce8df253aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a47d28495211f80690736c6da309e065ccae965c402a8c632210528ed67d2b6b0ca2bb1ace8e957a3d31e28f550c4b8e7b9cdf69861cb85102b1a63ef9a408be8f32af6793b562c4a39316518cfc31b7ef373ae6d908e2e03d547075dff312a33f2566121e5c7729199b765c9f20293b570ca5518f475a83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f7e118426f9ef4b4b27bb3519d9caedb9ba8dea7d051f383227d29f59572b633c30b83963ebe5e31e2d011bbbb6cafd16cae3d2cf044378bd0ca3a58068069dbc5864169f9186cbfc5daf35c8a32209c95c0f90ff549ad4cab1ed6a5da3a826fa77f221c8b45b8a99ce6e10bcaf19685ef397ef5e448f3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa5803b6b8635224a0ac9c0a57f42d9c87613efae830463cfb5ef12fe2d23ee7564de4f48f2c8e2d402b5e373431cb01114329dd1e6fd786c36f55789446af25a19920d6dc871c6bca9719e0feb9744379eb7d7b488abd22bf2286d076f8ee13bfa96200e7c6c2f813b273212c492036d7f241c9ea8172c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec9c54de79e86bd32de57fd802cb644a29d716790c5b159577fc34a4fe5bdd0950ba1ee55d5360ff3d5fe4469831623c206c6047472faefd0dd2a62eb286535ab9d84a39a16a33a004c0704b0c384db56c152ea3ec5eeb4c71b511ce0324addc6e04ebf5a447328a7d87828c245fd09bd7f4ae14da606f26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b116b1aab4e6879f904a13a84376a74aa5ea7483e43e6e5c44843ff7c1c1a524d927a35dd8818bd616582376bdc7fdda37cd3319af540373fb4881e189e70f216301ae2bb6c3ef1bcc91ab104c2e16024e896228aca21545e5ded0390009548179576217f2f08141240007b34048494750f9e4d0adf9488a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he38dcab9f68846008b6d2594499c394822f3c2d4ba5f921421cbc8726d41c063b1c3882cea9fd1242d7e8079ba746895128a2e31bb88c5d83731acd40470ef6dec3d8f7d0d93915590b20f06e236eafd1751a7cf379ba34e03c235839b79db713ea5ed1b87af2c336b38010137eed92d3f9f02ab8675273c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca1ef2f879c0130a9b8fa62080e4f6bb82b6fe309beb3f1656eca7fe7b8fd361a2ce54a539a5abe93d21f4dc393879ca34462411632213b9c0414f55dd598c4ac04e289e92e399ee0799aa862093de6cc401ea07ceba1eb8dd383439ddec35a18046f6979adcf3035515e0c17e88ac2394136f5ae92383fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1315fe5ced093d42aef955f24297fa97d8e3d92fa54ffaeeacd55ce3b6ea9e32a6374be7ec948d394bccfa05f08e8aab6658650d7adc6e5ef80f34630e876f5ebc76c5f03fe53cce099bf8f8fc6f166beae63239e38ecdd3f5f555f1898c92a37c4a8f42a31a70d28631a8bc1b0185bc31ed759e1b5a1fecc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178587e46ced6cc4a83875279a13d7903622f224320cf9c8282eb19da988d211e7e42746328c41f69018ec61e8b42b945bd81e7f9204624dcc84df7b233826a00e64da327b26b7933cac4e9e35c2cb725e1247b724409005252d2e4cdcbf67da352291ed4116b554ae0a178286b7634e77df9256874c91409;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h233e28bed42d5eb9056a12a79e0d5e9b10f6be238f9bccb78691fd0e76c6df62cc40111d1bd1ec1de25ce6f416c5b72c01710e068b44ff488c81c04fb6d46943d0f512ab5f17cf8aa01de10fb46c3fd0b2609f366bb9c6a7af38da176e5fe881c3768fa1b51bed03a9c26ab845ed25da58de19e6fd8d9e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34a64f01fd739f366878b34150590a5a6561fab505ada791775f7de608337e814a8011f56a0ad1a892cbd1c495593b72d13ff15cb5953cfc28d0351d9907a2cabbe5adc3014c0a6e2298041961c721ff274147557e855ee4b536efe8238aee46af93adde10605c28735abc92802b0d6018911e09e2fc720c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1347338a89abc0e79df07fb74cc6d00c9af430e39f7c3110e239cc2b6751df0dc8b4a6a64a1b1e359608bb8d9ff624e78ab5dbbefa497c73fb75520c5ca408980a907c70f2b6775327186557002a3a8b67a5397b8df4fefa96a386d0f4fd14816b461f95fa236b1907121f37b8f436c9f4d98fc3aa7fc5961;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142e014aa32a030ce0dc2f55b767adaea2505d682685f131836f14ddcb16f6880c39b87d8bd42ec6302434e9ddd0caf3469ac7b372caa8b373268ed97704b19a70f1c606e24271e95b3bc52a685a5d4c2f301b0f3fedc3de9fcdfd8ad668092d561f2b75249647652480e67d9325c64514b55c3f31deaaf42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68b39845d2f251dcb98ac13b51ce3652ad8c0a43a6a3f98dd577ecc07bacb71dcfe188a5bd960fa8efae4fcdce37b679b3142c9cb0d21de83fc4412d4c6bd219afcb006721432ad5413b7d9cde7f7b373b6a4ca5c381e06b3ec3ef9489998f806e397e99c21595441f81bdd906808f56412d4236bc3ddf9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193a9e45016ff41dd5136b10b94d0b8f723cbe1fe4fa7d9f69840044f600c90453da80acc7a154feea03a1459acbc767aceed5f9d71c6443ae05759d2922298b60cc959efd9cde51c5e1cdba2215f5c0e26ba640e75efc41b3d68e3d25d4c1f8275a928f97c4dff9aa93ff3ee44457c9b3ed7d5fca1b8c279;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12237c68137dafaf3fda81060884b6a48dc57271a371c3950e034c2b30c60ffab47c1cb711f119fcb31793e970885385a072358b91863da67c3460e112e852b20d6b0905db1b5499f75ea64bbc67c51046fb794cbd7c61e7f642167bb41a60a2d8f339dfe40b42c6e96114d88720865ad0a09efc700bd8b43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1835c1aeaf094b2a4a85a13cdfdcb9247b74ef058b549e8b9461ce6c2bbff46c9b7ae999b5cd18318d1837b0e4c2f126ac3c4a30157f61057c283361d5a1a1866346964f7121d8012c6ea878d64ea5ca509cc2f4b69010d25ab540dac57b2c1c9d603b4cb0aceb45aa757a0d2bf0ef70b3749f57c238beb93;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d6ecb06e061ff448008aa0263a9da17e2d77bde37313d772a357d26705a7a444f4173c9e84f4261e7a5b1b2afd670e0c494da2af8668d909a9bba5c6ab06aa387b8a2609411ba5a1c4055307d48a20aa8cf360e77e25dc4eaabc35449ab7a2bc08a69622fbac87a7bff26a58a01e8fba084a481ed339e97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ffe22183a25e6385cc0efeadab393b65dfdde974702cc04df6b7abddef44066ed14f7ac0fd2b73294aec67be1e5eda663d2da2544124395ddd2a6ccb69d1f2f6579fb8113df3f8189a8319c4bc5f3124361350aa9c09723879dd08d6f798c7b728831f32730971ff4873f1fea1aefdfbb202d2a0e38c9d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca18f52a48bcc5199c8383990f858e956d2c37b349d2736ba5c861e29681f0826f3f10452acad5e3dc419d53867664a666ae3b29ac3505d8373ac5d270ba67689d2eb90d57dc0eb22506e9cfc932c0f13f6451cc4ddebf55b42bc95266ccafd675da261d5b1d61dad9a1748d4f6f585b72aecf005e92c78;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77137374b2ccfec3064c90455a077838945ec932a60661cf6a0a17b5b83e95b08798cb92455155c81a0860e92e6b03a044fabe69ea68cae02befea1e29529c42afadf72bee4ade23156b52b12dbfe0bd611b517d7b5f123f2d72e9722f06915a12cbe9beef27181c3f109ff358c15191a17d1f96bec91d55;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a66ffa34ec243a3fe4856ed3794bce37d92424062a5ae376cf5b3954a88245fd3133cfe42b71598c2c80f93a5db133e403e746fea105954d70ab0770860313f389bd43f4efe8049d7bd194c461e0da662db069c59b3c8c1fa056826e94a043021024529998fbb359bf4b4fec07ae3e5ef6b22e84d4e7c4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190de362987424302cb136381e75350b8b89711379b23846010a14e783270c5c0e486737909d9a797d90aed0434663304380a62a1ea9725cfcf93ea218b2ab52d4723c090ddf7ebfcc49918448f713decf25e9d505ec2ae799bbc0e00e8fc89fb2c0270e21f74f0f69de45fcfc654b4e902a058cce00980b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cb30cd803a930291b05e8f2c5e7ee1accf296c68a5bf08587b0e92efd73f97b86492d29d592c76a6a223687ba8733449f970de19c2e34e781c2de8dd4c21428ad984c55028edce415ba2cd12eae0af21d81b9f50e382c6b2e2f619a99362fcb44a4cec85ff99f21124025dd64b713619c801936e5f8d4ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h922615f424575cbb559e4df19780c7d5a2192126c7b97c6a424d28f2a3972ec0317f237dbc7a0f6b139d352ce2d81c357458664575f8e255adf661f61475c234fe8a66aea7f01266050eb845aaf9a0c58116cf2bf24e9d15742415c940a9c748d4cac7ab9718d1e444b3598aefcc83fd03cb5fcfa402d7c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc0d4866cbc4ed0a83c0ed38918156a9677d7e4f34a7e3cf4317834a1461dd342b43503a1a836c1f6916aa117c0ee517094aeb980e1d94157cd6f1ec120be051d895bd909f0f927e0199e71c128244c90dabbc14f207703bc320ffd8dc70449ffccd4923d654275a9c003e8249fa3bd6d04763cf70c05168;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h375523f0b4f02dcee25795896dcc1917a7446eda8df8dba7c68f404c0bee78d2a91df59869aaaa2fa8e7a63e838ae7f69963ea0887aa460f38ceb46cc0a45566ed976614306fddf73e8822bd1d570ebf38e618c23495ee5a6ae07351619f2ba7ff3e2b6434ffc47c742c849265dc4af2ee9931abf2a63472;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c97ea0ebbfe65b309a560a5ab524428eb5e00e32aa4b67e020fd2decc866c34fe1e5696aa5f33fa5a21d4b305c59a381c8eb525c19913b15c50a3ff0c02ae70db83cac38a6367f8f23fa1903a7197c3d21e4f6880052bf6054da3e91201c582d6373f5433f7c3726e5a4fbe3afe019a454e908b2cee6769;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfadcc435e83271e11376f2717a9ab6fcc9cddb84d3aa27e6af8f8074ac11dbf54bc9982483c4e0838a01ad83b6553e567d8bf7f202847aa355fea9809b15d4bc8994e050717541a6f0528275fca0420d2cbb39ddb606522ae6599ddeeff632ba6b8cb0d3d030aaed464ff17513fa49053899bd06e659690e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c50444c08ad08ad69330e635d4037d03ed6fca58e06a2907b5451868f753339741689ba2007b7824815973e82a20f30c49b0696aea6117d0cc136a3a890a8dd7dace58b502cf699e1c540f7c5b4a05118d9134d70171d589580d3e8b5ed6a4c6864b2ffe061b46fe1e1ad2d1c2c1e9afcd07c8c34e9a912;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7ec9a5749ad7a918f3b5ed6518e27826ca12a1737cc6da94e599a142fb4f8531ee27f0764d065ca9aa1472cb0a6095602f2d38fa462d263ec85b850d6501a9a5122b9cde908c43e6e2a192fb02b95fa353a2084a15e9f2071845ce75c4421a4b52795e6f67535d231ed3d2b2daf7ce99998e93d626a878e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cfa3856479509eb129871379c8c0b016fe4fa4f0ecec24d36ffd158b504d02654c5bf2a3e418ee09f17f8c8f159774108a72d54274a1f9af9bf67900859f750f9115ec6bbe9e97d211174885a77b8076233eeb2170dbfe6adb2336081f98a0cbdc2d34cadcb8c136a1361373fc81fb37f4f6a0e73239827;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feaaa9aa839881fe2a13c992817b7341e59783a44cc5bc9c37c5f557d594ca0772352fc8cd2f645e4508b310ab065af01a38d295611dd84ca126b6021913d37da3d2ee42b455e77b2a4c8aec1e2af581931775c5ad0bcaa1596d9232e02b45e787a3711f6c4953e6d1a2815c28ac271cda92226da467d056;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a5c4a59f863d9c739f362e6860e4de1fbe0b4891711eb13dbace801fd4940d034b80854b4477ae4e0c54675d6b27b058b422deebbf3a22c0a65c40762a506134b754adc3beb361607ea6ee81d232d7598dba572a8ae34df84d2d553d183c1a56fb82c5d4669c65d04c57f89a9cd9089c2dce05b68649c06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e2f2837b30327c2453b0fb42ef8a42414dd4c95d71a9055641acc04d4c2fc8bf15d3c0989fcdac4bf03a7b53328d9835af6d7fe0e5bbf33e88bdd6e7cd09b2df4b1add984f759fc913070ec29fb04229a28eda32aa146f3f02cd08a8f33a79d56348e08edcd2aea872fdffa49914aeb2c19f29a6baef804;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb20ea0b4a2808ff62d4394e1979798c0a36b097f766f2f6d19e7fdfb621dc21b6df3cc7f126d58b0b6ce88bbcba178473cb00c7d1981dc17cc0ed4cb1403160b0df77dfef6746fa86ee69239f8dad34bbcd6f09c77ccbb0ebd87c42062f2c10c909fa0f91b7d5297db995015b6178802d85a2f528b56d2cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113e0c5fcfdeff980575b046807ffeaa79d0b600e99f64a2384b1be576f1545262d45a054a7698f3ef439957ef5683289c25fc1774e7e23a0948f064840fc1cfa952f64a3fcacfa6b65a647afef88d8abd285b1fe3bcf42f521324b6ece035ee0eddec90cac42e998584d0757ef5c2bb5ec2a535956e772b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef35ecad9828bf6b13d2c5396cb11ffbc4661291d5716b5a305439c24ecd6675d9cdf42255dbee671216fdc1855b5c8e4d0b018cb35184c25cb2b701f1d9448cac9398a1f560d0d47e3945bf805d50c9cae7c2b5b547d1101c446be71369ab8db3a3d66a315968f8deb3eaade359987ac48d7ef6d4ffc52d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a3edc3ade1ddae504905e4de635ed3cbe1bf04291d9cad845f81c12f472713f4cb3964ed2d16b47808d799891427b35b9e171b27726bafe6c50b22d8a54da0c81fe44a6bd3589b5e050827d2dd82fb0dfe9921ebb68fc2c41a98693be40c5c18b94d8cb95c133e966d8477bd300116694ca1232a043cc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3612c95e31e1ca84d4b61b223ebcaa9c6deba8757ca6817b056cdabd01d267434997f389c290c5684d83254c9691e98024defcae8a16ff9842369184e68402fe4f39a30f72befb09e22cb49eaba20ee788231ea9ece479c241de2df7bb3a3caf3a40e367952dcd41cb618ddf4aa32ac8291b8069c95022be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e0b75fec8a6ea7671483bd682e27c53002956bd942fd7e6e79a30421ed7bb272c99e8467e01ca4b1102adc81d74db1cc769a8ce72380adb4969849450328f47a0b073fb9da0b51cfe8ae31162af23f6f485c08ad81e08e9df00bf5bd1a5cd3c8a14684041ffc0b1c35c75764b103ccfff78522d82f8059e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18041fec1df38b3be73f8844ea0b3fa46e112c3fcb373fd214588142417742a9c2addfb9beece1ebe9e7201b66343aa3721f0b9eb8672f5c6d7bc8f410809a408e3d5f8ef847e8600ca8dca2e67daa3d9386e87561eafa7fdc01fa6f2e9c64b336c61967482e71df78fc454f63321e491363afb596c218350;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5f1205d390acc9345d3ebf2c4c1b96db45506ceb49537ad49aa95f7d3458d6d4cac6f0b60b7a45299ed437d9ad65909eac6781b6acdec6c5cf2629ff66fdf4c83cbb7276e4d1d95a3d66123b91172024e23b8bba02e416dee58c54f69f36efae4cb645e3e33394cecb0d6cfd1720ffde0c3bf5e6e2c3600;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dcb2a3aa7a2057a8331d2e73068328a76c76a5edc47c28b88dfaecc3395892e477353c270355f8363ed0bc0cd55d5ac4a3a5107c525da44cd8763b7804a3d54c4b92d88a5a99a556491e750b50621665300b4c21a20a4634a00a77cb8bc621070851cc123a1ca9b018ab73d9b6302606648fd236d50024c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1878257b35cf06a79de610eb6925ece18e5667dd65a4d8f151f19395e489c1a0148024bfea67b3d4e7778c8897dd58ff16cc47dd80ffbf2980ee82815e7e21b90a0e991d7b15b2f25c54c714578fed7e6c735fc388a8984d00eb7e341a4665eef1a6ac3a68c08daa7b342ab80aaebcb39c956231732d3795e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e8ffc38bbfeb7bdd13d09ea321fb8f1dcef044f8d764096b1511366053b404491ba74d8d1a83fb9b9dda10c811c8b8a20ecc861a6dad288e373e07ca78323baab8c8caa705c1a1801d7a59cd3e2b4987ed5f5bf33a69717adab7a90231dff153b96379d62ae5752d2dd79bd6ffdf4e16f6f82492bd64150;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5295b0250b5687889639ee74dc5cd5c77de145d8141f3d9b6e854f030ca759235dfc59b04359024de21b8ab36efb92f085ad2cf46e820511715ccace4350699e0b626fb9eea1f22c2ac503cc7e0be5355a9517de494f6996f6274477d6d689649220584762df2a7c02b00f489bdbd3254f67acf3cf4b947a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9b4cd5d99bd0c7bad5cf3fd83d059880ae2ef107a8c5dd491e77944eeb8c55a62f3ad6f51d74d28bc1e122f1cd53d40170465835177fcf8e5273b3476ddda38cb5e3ae92a45f090ccb3a271c37b6f5dfe70b400195f072a8b0c344ac60c3e6c114a677b42d81c0f8b8c768c76fcd9fc8ee850e1f7a6d333;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c35c0d3724d2ca39b4ab8d084de886d566b54b43f6b61484b68958b5152ee5a2a46d9c9f2447c3b763fac228b04c6a5ccaf1a5daaa3459460f8f778132d1d7a36210046bcfdfee06095e0f86b05d5252eda92cefbc2ed4ef43b2219a188de983c4a0d2dfd6d8f14cf5001c3e46e8c8685350d87edb94831;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbafbc1dbdd04fe330321e896938b452152c54122a6c35af00003284146f4a6ce59935838594187716665d059722ba4429be257305a619745d0869d57303d2298bb982967919621a27adddcda1339a9a97f65757ba7862d9f2ef05560cee713bb40fe8d1b1905d85959e0addc3e8f6d877aee9ef9b8272f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3eeb769ae4f6d76048f7ff04d5ca1099c062d5f36e3d1f8d854ab523deea0c2dcb26e3fc3ff344e1e3d8a9260877ba7870a2d6ac7cf68bafe7a4cbbbdd81cb8a52b7cf70df2f9e0e62a5edaa9b3eb08c8b6296141b61a0a007a7bfaa54afd9f71878f293038215ef17025d3e15d436a2e42e5872e4b3e307;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58b0c83dd28879e22cd29ba8c82fbbb633958b5e6bce1bbfa56620f54d34c0f54184621084f4fe664bce59eb64d8ecc998152926b883fc0c4070ab813293bc6352edacfeb4e8c3765d942df36c6b61c024a407391fe7c3b9ee49baf086cf024f6506db8194b3aa348c90cc1143ab7920347269620b3cba82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47dfebc7c4072de55aead4ead6674706f10f5ee42bbb71bcdd4365b3a77dc36f4a22027e5ab1a086b043c1f90177f1368f2a8c470b0e97311df74902bc8dd62ec8a5aeff99008bc173277a9fbc31edc3c9526e7ce90502eebdecf44ecdc2b1f58c4aec9d7d29d942cffdfdaf60803e1e321a7a990521e3b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101bcd77de1ddde2fd1485c8441a43a7a5960fab9c407f6ba2e55d0d7630c367c67ab1e5a5551f15b88112a78494761ff7178199c9fa2a6145b069ac549ee30fe02345bfdf34438794e2d677fa4a667cc5c713bb31630a2f843f9ea88fbf4c311553089adb15a8404083caaa66634376a589771e120746856;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bb89d3c2aadc5d3b395c3196822d94c436af664015a1da4f23d3041a91a3f38cb14fa476dd29d71fa903f6b76a8d29e2469aecc17c810612d88f4bf02656b777bcff461292d102c8ca56f7a9f9d415232fe90869fce070787b4c5ac29ef21fce5d44e7f645ab190d6207267f0c29b9793f3a905dc1ad4b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc47642450a3dd89a0d96195a503cc846222df92b59b7544bdaf9ffb317e7385cb27636d966c4333b7f50c3a0ce0e15bed6eafe821a4dcf27bb2b44a9b7195a3131975012860736efe565fb492f676bbc9c97a91b1f37d944174f52e060dab2380ccbcb29d2bf46e44a851327e5e5f989752e73e0af1273b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa477882f19c05ec651b016d7c4508fdb621c359196a0e54264b5e31da3c7ee1c9f56485386a38637fd073dbd182fcf4380715ace861da9f72191501caabd211b782c8cce93a234a940856656b58d1f7a18dbbeef097410d460c75285cc507d80959e9a56fcdbf860f15306b7e437ca11a47431d2027734c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha358db6834adad9d8416148fb0c52344161936ed8965edbd627e3b9d34fec7c732746fba369e1f81f35022cc9547ae30e75d39679042f918534c3cb71f557bcb6efbcb07127237b307fa971fea89a5791dcbbda240f02822ddf02aa1655809aaf1fc73b772762d9742210eaa5dd41e0b1035b3dafc67a92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb4cdd8d86a83895620dd63a7855138881d5b9ce8f208132a63cd4dee759cd53e73465dc115e58681fa31db0876978fbe3f6b860e475ef9dde5d028ad4c2b9623c6314206e20786b7322fba2bce4a5437a9c4e29ebcaf044b66859ff93891c80a17cb6bf1a1f28441c440bdddec2482fa7bdd90b0a73cd5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3212930badf3cd8dc6d040e825c43357ed751f3745d153fbed08396092602043325e7dcc6d2c3e78bffd632f41100ae2e8f05b7ea2e87f0ea5f95fa4b5a7f5e2d2ca9b21905d0b11afc574a332e91e4fd08906ce35625651c109a2226b7578f3b0996de13eb7bbd29562d8a788be6abaad3964a86b6e072;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6ac7b24aae7fc85960f21f12fe265e72054ed9d1d9b5b052de0de642a5108fbca8427bd16bc60843764bd4127f5dbc579e0a3be505b145ff933c68aecaa2d22460841eaf00195de9b61f1557ba89c522d720a5204322d4dcdc582c5d23c54d98bf3a5bdfcc385bd9add08cc309369fd01b1f4c1b086aa95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed8fd243113e827dbb6ce9d05ab0a9a951b702eaa0eb02c2cdfa3344b64fd1fd1a2d1af72d6df427d69e05a4136601dcb20f88f630bd46366f0605972dd28d8cfc6b73d36c2609072eca88f44e6cedd2fa37ed6e75ad1e5aa8ed738c984b0ac47374d5315a547c3fbb93523e3fbb09421a27b9440ffdfc07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17098b9e06b6cae5db7646a6b4a8b73ba0dbddbbbda48d5c10353f00f281464818b4aabb4f9da86fcd78603e1ebe99740accccf0cb1a71a54109a36f926836e1c217979b3ba599eeb6ae7b6a08236f37455d81c56482d89a269cceb1fe17e39556c0d62c4e676505d4a998322b0ff9452ab5425d04c4d70a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha818f454c720b358e8fc81eda705f7f108d7d865f9c9427b11d39ff292dc2861d7bdd757d5969e755ad27e2fb3bc3f57647fdc711a34038934aca2eaae6baeb182d8eba69f3a64422a6722a98a87a912b935bfa93607b91a0814b3f9cc9646ae7ca6ea7041ccbb94b39a6b6035c41c313bb2f88879897df7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0a6e0a4ad9b55d7ee5936d59fc6e7de3ea47b67a096f9c9562c5b4a4afb569ea00ea7ad33c2ea35050d5309c378ba6ae7a5ceb1470044706ccbe221c3c3f4304de2f39a3a5ee9938f04bb29e92fb5709dc430a38f8ede75b0a663a43ca2d8accda7462970ebc7bb37249866f0e463317b36f0903ba1b2ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18357e4baca6951efb94b87760c4b098e5317ec97ee9212ed8b74e2661d2c809c2c00a52601473b156a1f2ee9691af81190d6a02dbd0975e0e1cc149c8bf7cf53a9a5b3ac0edd4c2b228999262edb5d40f53c90a0e86f6704ff9da8858c30c0179a477f3413fccfcfa7da25c101bdae2d85602bbd30527d2d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ff3e9cfa510dc714a68de842f8f22ab6cf57ddfd607371251165f79300db1b7db79a8a2f64c2cfbb9fc41fce238681cf700280bfbc9b7873c94e95fcc6091c5aae8f90b4d0dca2ba0e00c613158849b33aeab8b247f02c9c66de9103f469ae3807c1822d9903aa78adb285bbdda48a38104e9c6fc56bd1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb11c687ffbdab97ba875823904de80f73626a808ede2f240c712c36309951d00a9696b1cb095a7bdc2dda714d77c92e14be205c8211c07d07b842da41d1c0de70f22162e1abb3edeecaa25657f7de9f3baa647c8ec0b551cd9ca7be7405bc1706a4ea046dff9238da03bb7342f2ec04aa6a3566fbd05231;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148c1885d552530903a09ce6b057e3203fa7679a254b5077a8b71ceb0d00ebd110121693259b88c02afc39edec6f7956c669554c4e8ee7426d327595b071e3f1a998bb97d9503bc8684fcf48612ff5dbf857f3516436a1c258fbf781376087f2e5926aa897437061fb8d00185c039659578b287f0101bbb67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1446bbda2ad32f8aaca09cc25ffaf8d4396b739291619b596bd2c63b80eec3e0f815e642d6c755ce36ae5b4cabec257acb06e9636532d6b0a21657b4966a29c57bf7db5ce9b017f5e610ce6d744e97cd1a6f8e3d0fc102a28beb283fde917ffe66d9474de5d44deb683ea0c823b71d7aa6c3b90116c8670d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c6db1aa5910cf37ff87278a980749d8589174a4b7e5efea88e39841bad49ec689e56b7edafae64b7a14c3d83db138f7c7ae9287bb98143500cb6795c21287fbc20e709ecd73d317a284575e3aef88290a0e2bd6a36c4e8dab1b1b5b44c55a3a1bd57666bd5fc33eacbe40cf2c26c14a00ce1e99ac61df8f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b86d85a99923749abd2b4c38e85ffeb2edb43758c1c001e72a52c1d1e7d6a18e254823b6bfa4dbc71b08c0add14da86fea172c16ee6afc1524713249b254fc79e3ab3d6b67c22f6d6658f2ae6a9609abab8b4ffcbc969ca261f79f9b814f23eff0a65feebfd6ef734ecc1541877bbd43e28d0207cd64534;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dfa6db1d145080038fc55db0694437941590ebb870d4ece147b55d03c0ef90dd0c075f9e6fb8c04d98bd360e9d9746f0d1658d36d594c9cfac29fbca5e9dfb465662a8743f0b92ed87a82ff544dc074f31626060811bd3b909000f7e616d90f12903e75be93d441295a005831ef711cd1b7f3eb0fc6ada91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99bd3cb4d19b113992a9113736c2cda44ebaccfe4755e9244f87dce01edd9bb08dd56cdfdbd34a4cbdbbb65f9c3e8cba98c61ca8bcd95409918af59eb961bdfebce1fccdb5c9737f0745391b659e582a8b957505acba117bf4f3cad95e40a9f26f5eef24dbc9077065b920acd854cb6afaec3e526082ce10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169617eb215c531d837e145f8c40cbc9f4e66026e676b6de7d09209f0523f00e67750c873fea23947d669ccdcd461628fe26c4372e106d085b3139386bfaf5ce65b63ef0b0391f1bd93abab9d5496bbdb9007d1b46e862be4764f1c0b51e3ee667d911b4041000c733f07afa03df1a4b8f3160087850cbc5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19275d033d2ec8a7584a577086751f294c6c005e270e6d4112ea7d3088bf9c9797ea951c561e8a8fa15130d8407ac2a5c5403b8448ccbbafb817a9ae209ec06c473cd699f98ab53bbfea8a3887de14257452a26192d855e88b7a13df2687948f771e9b20805528b549c6a08df92df93107fbaa3e8a04fec28;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h336984067d2c3f0fe02187185f52d13cb19b4e4008fa43a6875077dc534d3ddf4ea2f2e2657e023773d927a5668c4c4bab514c5601b74ede8c75b6135cad00c5b31e40236023eec77eb33a6792e61e0cb7a567e4ce22882267aefe919f0315342d9b98cd2c926cd0b46e832b8ecd47b8e1a59af1b982a39f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1751a5117f8c4bc4ada07d49751b20d1c1a6d123c1822eeb358f327fb879dfcc778349edf1832cc6d0d2a8e7cd75bd9e3ff02f837b736c88484f8e99d7482c62c6bb93742432ecce1b3cc8a11460039453c48e2b9a538f01d1af86a433918e3a716e5676cd24a7244429f97cc6993a02ae4ded86d02274a70;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84391f2b9d5b48e88c954ba8e49b94da0f64dd9c57c201457cb2ca335c86795e591c5568ba9f7b3e3117e7f62f8e71500bcae1de23648a37d2b05a3b0df83e0844c1d93c3747db9c55ce5a974a670b2c350fba75a415ddd1246b41547e0c194b080566ab9e54aea8c49ef92bb089e24acdb92b6b30bfb97b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d2ae3b4fc7887320eac982b3ea0e56d79237f17f794865dd741c9d43a924a643138af6c5ff920c16014a75f2ebdf59490fd910139c06cf49e7852d4fae12a5012fa3e27e79362a4b630185d1416edda25a941ee52affe446f496bd1183c26067ea61df2b1738228620c7d0ee1f44fdce8c9ac684461b681;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb93b6686b9a2a4804693d6a7052f2f87ebd506fa2916b01a973d890a1dc7799604817fbe1d2db583df7c717a8f0ee9b19d5bab7c6bca9905e383d349a67ed71280fb246525f4e90d9c75b4e51aa1cfdb47d31638e0bfa0e099c3a65f619cc418d90ea01c1ad18634f8b9931197603c4d444a7e8ced47552d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156544e654df2872efe7e3c8bf405382ff33a68d302e727d349119d5dcc2c459edfc1b5c7cba2325139bbbc4e3bca3a91d882de3d24f66e06a87d15bae413c995364f413026f4c16c9c73177340c8d29dc5d289c5c6ce1329a87ecac019661eb45a1043886b8a4bac6f48d1121419dbcac5891ab1057f968b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ef95c59658e499b9fb70b2543050ba38f9da6882af0f960ec2e24e2abdf8a136415f1a571237309be4b5571edf7ca5064951ddeea5f88e0d7846a793b4ca2898111a9682869416a2eaa5cfbf1de661f8a639b675b32110af6cb377b1b12d8d357754dc5a008023dcb11da105326a2b9b1a10ef32e9b7aaf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h830f4b3f8f334b699766d7bce5be7644f601b7015dbd484bb3e3dc4d540ed31da8e8b33a1e394abc81fc38f726102e67eb94686355cc88f47a980f4faeeff4b3b510de2a3e96974291f209c584a1c0f6a8610ff574ad93a777db511b37c9a4d5c4e35cf002b2f50e8ba6d68b1560195e7e7b93f9ea778f9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14deef07e02b5113f2692e99a8294920bdd2468e305696120f817421eb6cf79a31f5b197c6f9c807fe934a1251602385821cf528a00f4eabdffe7572e9c7034441c9db8066db6b8d8fab0a38633dbee076e91723904e50586445e5cdd073442541c4816e341bdab5a4afb3ebb3e6cd451513df6c8b2d3d29d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179182d8c40ec76cb85a6d16b9b8b8ef060e03868b1beae368d4904a7dec74cdea9d0576fdb8e1ddf6469513881ade66b89ac6401432fca9e336eb9826d233a71cf34016e60fd676584366e5d7d8de4d9e0a116096396d59cd545d1f9d9f0db08401e7c0a08b7025f023d5870b506c00367104b7626568a80;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h788f0816ef1b53e93bafa35bca6f152488d99335474be2a1a9ef2ff032542b49c2e4f78aa074eddb7650339cdc28bdb0841de7b003cdd034e26c24f736283dd87f95c652cf2cca3eb95e9007fb074ab99864f6fcde5738b6d93b83d3e3b0a2dc540ac98d54a0adf5638ce3e50ac4e3fcdc32f7249e2da548;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbda5a25b18132e78ef5d09d4437bcc56234e124b8a0371cb64017bff5982632fafdc7f808ce20a9cf62ce0909e434b48150696577beb0c1bb8f39d81a95bb644ba462da1cce270d3d73076513d430655b0ca68d5b7ce152090351cd6118231d2964ce9c5f7d105f00e16f8459e6498d756e715509aa309a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169ee2aed2504bfb2f614b52f35d73df3046b6332ba28a0cce76e6876237cc73a1b167f3f2118076831721d365c5df46a77ed130aa16f8ec44942d9c76d662bd7c96fdfc489066f90bcadd78faa3561035912f5ed6a99a40b0802d5660aebf35f6ed88744b78c6d68721ca55121447674ec4a474934fb6277;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a5b8fa0eef4a73a1d6538df54fe51556d55a754860c7f41eea4544e00b382a6ef58152d43e2b51fa23ed1c7fe1d6920f7c35067f9a7269cd9aa57f0c84a73c1d254d9a9ce0d5dfd09142ef2a4e1b0a0efb85388f974622fd8f874b7668c68b39042d7984e54a0b65fe38145d1b79b4b1696961bd70ced42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h994523ee5afd46e14031f206001a8db22cbf64c7e58ed6e286c1fa5aa2707248ed87d875036cbb484e7f65d011ed702a723df612f65d3b119dc46565c90549b3e483239adf5751a5651ef4cf331a70fa145e59a333247114dfc68cf20ef38f68969e0293e06450cd04953d4815b2a61f0e21857705d74132;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a465d2619c25a33942404d714b4ba682197b9ed10ba2320efb577f358d6c950da95926c499be8637ab36790feb8a0fe47af3c6078b1939a80355db97f53ada8b0d7dbf017b6a8ffa66d4d7b56b2ce8b758e1d0e606aa589626390f7298c1c8ca0f8460be88c0c26f07f65520dd4780e0110819bdaa79036;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6939c033ccda0a4c3ec11f3d27d10ca72469fc8756f3c9e9fd12dec75b738a1d7398c6b398d33cf467a5a51d54847d1ef69f16c9c53e6e3be7b4d537ec6cda677db61b65cc231d3587d168628e8efc0c1405469125c30625399d69c798cc553a023073228b01cf095582b2be83536f6923a787d93cb68b1e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16da42c10d6768f44d4c217cc24115262a3e4e9ff46345c0093f6b40ab1c2937fd986f1538d7f28cace55e8b9a4eb0fec0e757cfff700ebf70d435b853acf35f205163845d8685fb5828a790a870afe0d13659ed123861202ff2744b1713c840307b1dedd06bc14274bc8e9aee94ab78a9370280ad3042d57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdba37afe81f6d569ab99faf509a54ca00b9a2b1b08d0c0b438bb7c3cbb66c01687d9879efcc7801cb924473f2849bc64dacd910a6a6142c908c89ea1c1cd61377dfa0de8943b7e71848a708a6f36338318f2b36bd2bdf9940545a492c8374676f737cbf62b1a2fcbf265c4064b169d3392964c87587a637a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h602d4e8c309d3e5df997287aa7d6e9122a1a46f83197d08612ea9e355429c61e4161d9a7df0011819667375e251c8bea3ab5f02e5f77a1b25e24f3eb6cf27e7b8ce7f94c23377a28f5bf7fc543e9e26ea6c9a362280f4169fad8b675ee5a27f47b741b6287afd145a16ddf7fcb68702ae27a9d11ea1409df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f10cfbed8ffa8a8493ce8547f80de9bb65413ae3ed93bae6865307aff42417bbac81ec7865910c2b14d9ab18db32eb922777f4c9636c993fea7146b08bd5c8fa0d7755586fe081cf0160acb4414971dab77db8cfede5d4d70f989b52100135f957162ab9738dd5c5cbae225d39caf0283c55553aa6354c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c673083bf8544e70c720b2a8f661287846035d9d6544bc758fc9d990b1d2f6b4759b4a91482dac800f2d1b53b262d5b6f868788268879db762e80552e9a959bc42b0270c7bab3a4eb5e6daa1c19bb784e4295573829f6731b43f6a43dd15c1f8f168e1467b557784dcb3a9524f8fa36469ba41b7cd66f33a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65149fcf3a4e93ec95a19d3045dff25c67d6b1eab00f76fa805decfb4a09b01038fdfd046f28c08fc411c020ad1b677967031d634c225cedf9f9b7b3cd68d8853a9c8bbd930e53cf207a528599a1a74143a2b488e00f0c08a64bf8640333a8e68f608bf441523ee988e5802c9e78ca3cbe21c68d9013f249;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef57ed1a75bbd992fbb1575f3d0b231e92072454989091b55d1a797ee1b6764d0544ff34ff0122d94bc71bc94204453b3dc9700e6a900201cca1bf5b8523d478e859b493a60206c2db367ac411ca4e3e74ef7db79574a8c27ccd10ba87f607a08dd955292a10447378526e748904182fc1a445bd32e0e553;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1408be3db0af058e3d26e127e30ba392da4439274e2e9efc37bb0e4c315e9b9c91eb3fddd07f9dcbfbe57ced80fae27d4d819ce13f546fc5516ddd51d8103cfc7747ab3f10407742fd586c3ca067863920d6af9fa70450f8c3e73b068793e0e37673d8b8f2c94212883893f1a3199a335c279f9dcd8dd972e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11fb41d2a673bfbcb7aba3412959e72ada4fd81c97da0f57b8fd00c21c6630e202057fe905c4df9581c0542bfd4c49f58a5a42b7b20895f755407de6a3e57454c4ef73216909e5fbf2b6b6a3038c6d3ae0c1bdc79cc006d346ae54473e42f761977a0343fd92baceb1500842c1f8eeb646e90511354f090d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5d4aa3f8a80dfc2bed2a2e1209757d6574fcec20df6cc83107dde0b2dab31543ea189ccf29d8f5e76f6c0b996a766dfa844ce8814e5bd19057e7501b0a5dc8ad7852967fb6b34fb45f1aa26fd606ae60202ea46c5cb1178e0c11aefcb53676f230586f3a18e3a026d92b74c1ee8b6f8c4f10375e09f9cec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f999b10e23320a1f211a494afb4a99c3bfa6281c890f82dd31b1d9c2209be68bf4e8708f79e0d817f65897217622567c524f794937810db0104d6855378cbd1220096b00c20a3e5cfcb6d6c8655a3d698bbcf9d39bbf0e7b2330a34cdb222702c3a21b1ac17e4a7779e96f76c2e57e2f00c773fd10b0fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1397d1de1a5d903c844f9d2665534b9132bfaeead6705aef1341d7f83d5643cb0223d22e2808f4b7fcd7bc77bd00884747a3ee2aec49b868bb03abbe6be32365565438086e31ea897975e5259a6c4756e2cf1e7493597fd2e595c27ae18e98c9fb2780fe0f025c09593982d41a9f637bf1c722f945bbee805;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9d5dd9a0bad0f47c1fb7e56aedef06955983a728142c963438050d9c1a8badfa8b6ff65458445cc5af390f97aa8f65c57ba037d8b92318a18ca1d72e3f8e2d11b5b82d83262575ba1b86ed0651d012c29709f84d6a847e9f02f0968e2e7255b955194eba53e8bc8e7c6c4b037c520a74d9a57ae98705114;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac1847531458a9a62204e463b958c4cd697a85e69147f4ba4185f36af82c3aab9947f15514f8deea9628f6197a5ae6df37393cf18237d58b2c05c7c831f6c37684c5c3919662ac43323cdaad2bc5e1826e94ffd8013f31060200f724609b356c2f9885af84012513d0fb86dc56b7c82741415a4546504291;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h158b20f3090cdd938a673ca2c6479cb49456198e74a89547de2aeda2e76adc2ba3aca32db8182a5de395391a3e33ae191615f4a2b15164fe1cb8afc5e3a8daf9aaf9a192d45aaf77ec4e1df93bb2863a86a16dbf48809e1731d2772bc2fc94b5e0c51b80802848058ba5ee8b3b167b69c0d83bec04166c522;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43694bf7f7820924666e7246e120db3233884993e2cde012f10aee3d5894079320c3952855ef90ee8d7c3be1ecb10bb20a995015e61ffd9548aac243d63eba862122e4a08e5ebe4c3eea3ef5dd8fbe3acf4168b9ef4f7f3c9172219826dbe7cbb741d69e09f1209a0cd3bf5834009177b752aa3d7615d0ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce99298cb443948d9309acbbb2d8356f7ff264727d5359d08a5e04412824e7dd2ee307a3241b8af1382c7a9eca0e68638d97226a21e4ebb9dc89b3193d0c95b03c3550377ef67d251b8f3b35eb7e6b4f3ee1c9b0f1e0046d5e90a77f047c364eb6247ce121b71d5f3cb186d84faf2cb16b79685c8ccb83f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119f24ce3458298fc3da49fe217b1823ee730111a680e464d8f72e032748948fc980025fc469ad195932dd9e32453a28c71506b69980ac7395a10fe1d549cc3c3ac8f81ec98612ae15fa02f2e28cd8f199d4680bb171636b03135360c99980c9b0534de62726ef6901509263716cb94cb1fe685422a76dcd2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f0ce9f02b2cad7e7642ff395383df09380a85406ea73d20dda1cb0bfa5af8af8eee7af85eda802c543a3ea637915ffc328684b472e4db0036a42420af4beca149366cc387ebd2d5d4d3499b0f1c840b6d8016011f423914921be9f14a4c4e4b22ee769bb7b0c20d4ccf1238244cbfd4f3bae4b2776085cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edcbb1ce28df269c490a0080d704542bd292cd01501fe1871c97712bc33964dbb43f60e258b4cde32a4c92515e9c2e0d86f757ca5eaa2abf004085fe0a59ed40ef7acdc8918083b197e9051044c714b2dd9151b735472a76ad57d3f01aecf03926b05174c5bf2d11b48a5a20a42d29f928e1b693517c74b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11840ce968b2d18dba74d30d7ff9739767ebe876e882c4728d5dde74730b6873132d4ea2b7ef63493ad0474555af1440c9e3a73afa8aa7359bf48efceb51ba24b962662f0b2ca42f18e98dbe42d704dff9227a878914f1ac749f4ff5bf9c2736972f0931df24fe12c6132a3f03c344bd103ecef61b7e282b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c85e17dd2593c45c6abaf394d9a683651dcfd7bece970b06dab29b6aa3c48e57c3f0728342870a536aa2b87ec5021815951a1e132e814347117fc9f9deb20703d45dce39bc229fe922dfb924fe56b75e15b9220832e3fafccc409fc182d2eb8a412a6d6682ba5fa63ac10e60c2becb091f2bbd09c864d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b0813cef9eca1c86a4989b46073d11e78f2d428b3c4f5edf875ee3eaf4fe82c9718facfcaf4d46f97b46c461bda726f426400e9658535f039888c9b64feb275c510a86d892ada45a2f4307e297c0d800f82e9685034ffdb66ad613904b79e045bb06a547592c4424f839caed35fe70fd59fa05f54bcb00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1401ac438b47ebbd1b4c5b8bda148165530dac32a11c4f6703082b3ef96365a903c439692e99e9049fb966fea4e79178c6a79a6b5b1b4434b1e59340c7a6747b0c977c8a1ab4406987476afc1d721151837019f0b3d72e9f842d5f8bcb33b2a1d8fbdb81a47bb920d9f466986ea7215803ba68ab0ec435f6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1068763ab3e4c9037978deafa7e07a492aacc43a2245925867577e51d25ec8663da2d11d6d251949d543f8b8eb6b53e9a012e2f583c2af6b52f30476b60f2c10bbd1babb9cb6fca25d8d533613bb890830b0d33de8b2ff493e34baa205ffff544f726f03cdc9bbfe356eff509fea4d027ff1fa936d6ca302d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f3c7b0388f0a8a66a9f6bf5617d007efa5426868b962899c88f289736725fee0d53e056c7e7800a5bd9b4b08c7675c9f83a4b18a9876cc43bc638267188bcde0162ab0f72fe584f81f7847abb7673cb6feadf37f6df3c229eccfe7bf8e42262b5e879b0a942d54af6d2f48b40747cc02c062d0550a8269c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c39e8a6341574e8771b0f081a85b54c04441ea39d5d7de1cc25182a0f8b7799883583769831dec73cd9bfcbe70fb4b2737bb85a406895957ffc9ff3ce364b1a7e5eb5aff7322c6a10a748cc499a1acefec8f40ecbb9c4d99618039b1859eb9bba51dbf7d2f8e19052010557377744664ca2b57a480ca9470;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be58a17ccd603f6b11f0fd07abfad28142ae4820cf1884bd225a3fb7a3326fa8bdceb41bd2d96b35956d193cda561d4fdcec3240a15c9b934cd640be88615fd1b698e2ffa06835cd41adcf694ca418245f9f5d4e46358efd626fc091bcee414c6c068fcd7e5c3d9f92d3e6b5d46aa425472e2dc295e6c241;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a66af25d3974b1489d2e4643b112b8db713df778355a646b9d63ffa4ad30167f3082f7659735a917fb68bf477214af466160af5d3e862d2003ee48974acd47317b17f6e1c327148e5a39bb598e35276932ad11345619d739b47facbf0186a0574f5777c5b4d496bdef3dab892f24491201e9b40f33af193;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5903eaceaaf0a2c6891203bdd58454f6730cf31262797c94b221feb61baf08a226dbd10045b9bce3893a2f118735b10b566fa47b6b1080f415fcbbf4a72b7d1722e1b59789aec434f89d63b003b4ffd2aa7d67715defd2caec0c16b0c33f8f8c270fdffc874a7287c79368919b711ef2a86d5bbcd5c3c7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1745fba327d83881198403d5ebd33b14841489fc032460cc76952569ca18d8fdec4a0127d465dfa5a1b7687c7a37bca6d9cc9999a2aee8ca04901142d9d1482342318b21eeaae1fe238a6902cf62012b1b5f0cc45a4d97aea4ead63c8be28be9d8c85a4eae3a18c9cdbcf810f7c505eccbfc0124b97409c8d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e394879288e2f51f9aff57c27f46c5695410a5d828b16d3f039754d08e2fcf21ca58810705200de4c0a062b3463f0d566c572a433c56e0cb45693db2298fd218c12ac08d9672d0229b4a92febf3730d37be839548d62baa62e467f2bb7b748f751db380cf1eab30b3f3ccffcf8dfae160c2dd152dcb0257;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48c31b15096cb5bcd9066ab8077aed710d30bdc97d97fcc290a842cf7fd1c018319fdaefd85dc4a2d3e8bae92a10bdd8d1b3bf5473cfe1328e394e6791c9d33f63e7e2b53a4ec9178564484df90a060d58ad5d2d612e8ecd9cef6dfe37658fa35c0786ceda94b8bbf78682eec2a81674475a7a72da5dd6d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac3dad5ee85d258a91cb9e337319fbb786659866f0018029b6bd02ba02f92e67216b4bd7730b33f1849ad423139715b253bf42e15573db1b612255cb64a517ee445ea83d7732070517709bff814f6e60e7bc1402474d478fe809edbabd1dfeeec83a40a0bd90c5909ac7a902d9b8ba7c7c84be5bbc9b9aaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d80cba9a86ed2a934af169692329241933c11784a3525bdc56daceeeb64896822e6502817b4d9a9f0602aac1b52c34e2ce4216226130f874665bc2af7a4a725428d3dd2778e57e1258beceb6c9221e615a9182170ae480fca31fb50d7c0d407bef21dcfff61f3d4e522ced68ff61a20b18112ca888a404d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5b78a0cd0044bdcb5f2e1a89a4b65274141e1415fa995dc1e53dda785ab77b5b85022b26f230d7ad33d44d8096156106e46aa80cab257fdaac6a9b678379875111f253ab9540d4a1463af6a4e642738d66f52422f6277d88fce9b820a093cb64513d5d7d7802c1bb0801696d17d6ce2d07d42b9f633cddf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e4073dcbd1131d924e3b21434028e7d43d9d01242f8b117a99f3388e5fed3d74ef888b218fc96da9628561613ebe54763277e20a3bc6245b7c7d3cbcc6239b0ac9e814a7a5206505b15c72d97fc5d27902dacbaa150cf8282359701e9b5ba4dd163ceb0af3b42738d8852837cc9f278ca298af9e77995b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58a99236007cecc865648220218b667f8a588fe574637797fef6d7e7f62032abcce6b370038731d934ce8acca5d4a4cbb14753fe34cc29b82ee1676e609a0111e3a3dc500f4329ad1cd1b68db468513bfb160d2400afc85666f5c5d718e42e177a14607c392692ad315b3447212276108893fb690683da5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61856b19721cde3acaaf4c0255fda8a2fc8831008abb19e7065d962aed562a9c365855f99419877a077e858491f8b80cf848928dd4c2462ede47e68dfe301510cd660b07566eb54cf874571a542ba2c4172b722f4b917b89addfe54105a1bee3caf3c3ec6380c428283569cf8e11a82d5cbce208e43d9a58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111b2a55c87c9d8ea0d533e0167ef757861a306f36a24ecdfaf82cb3fd4f47329d7c7384632cca732905d28b3efd115078fd52263391e8e11d2c505f144413dba4d1d4b5a645db8d0ec981f3ed3539665b2661781a2a33f91f781160d2c1e3680248733d0ffdec099b563bb70c0c1df8d801d586047ec2b83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edc230a43d25cd0790619ea240c5de5accf66e4dd8271ebc217e7b1358393596fd58411ed10f6cf596e5be374c46c6fcd74ff01a3d2f7bc88086e8e583307f16c4c5b10c4d00f2348d806d5bfc6540f333ae87d2a3ad3b17c023a53c177eb98a4e58c268af7486d89e69bea11077ae7d15c9a5f3458e8af5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h385a482e7f4cf3508aa52a572531d7088ff1cb1487771e8010fb940007ce7ec3e13f8a6e5f6eec41a08339db5f7579fcd993b4c537bed184635229524163327428826239ba6d81c037f864ed09e96783ddaf0dfb175da8beec923e55643dc7fe6b7f7b6e74b6e918cde7fdb01fe5082deb5c1e6e38800f91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107c4e17968190b015f89ca821b31b80012d5ae782d942ea88b4b90410aff9a5dbf49d9bdd82aebd33854a15a10cf77ef948de9dc1084249d57425062f466305352a3e963dda6ee3b12dea9474b1102153e00bb3575e75ac0a8f056508e642e179a66eb0452fc98f7bf46c027ec5bd53502b9efd7a1a9a04d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131d756fadb4ea2d4c0dda294af6f368bb3fc99aacd0a323faed6fba5c8b3e25eac11e8a6c829d8859d2e1c29c2c8f72f1577c3f57301c13658d94677eeb0004dcd1b5df843b88443563486453a7dffea378dc20d9bbbcec9d063e4a26b69bd595b769274d0e33fb40bd1dea7b70e083367ea915e59227e52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106dd17d1fdff935e52c813e44d424366400a79740b7d12ccae0f52e6f6bd75c684effdbb4ea7004903439d9a8e6ec3dffc41d48c65c8e7d76b794df439554d9fb851b8cb4003196f0e28d338cb77433d2d7d97e150b54861daf1a34f4a4c7f0c0dfa41c8f1b855f2f47ae8697bf1dfcaaf65113976e9a05f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c7537fc5a782226a6e00a5d188f3b499c25ca9e42ca703fb17bc3e7e29476031037fbdb64389aa5f75e6c5966d0d59f83c78e7379f18bb8eac144a97f60d5d77cee703c0e1794ec6e96eefaa706a9eaf969237282f58d893d7e0dcb45c1cc5b6f4c461835c5051bf4f44bcaeefe32dc349f9af77b10e873;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a030539384d08f3a012e4337eb735ea48523d3881c959472bf99ea84ae851f6ceafd1a3716278720f7a00424695d3c502470e731161aabb1341686a39d2c399debe9f3fa30d1d5a0e6d1cfff4aabd723ab6b66cf80920d0c846ac290b341aae531840c849a5bbc702f96f3d69d3a3ed13d733f604f914c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6c07e159d5a464a1c3d5a3973bec59567e82c7e316a448306361638066ceebf99f5c7e0a4ec8b95ce017b2d6eca271a5cfbae8fbdcd71028e76e49922d5dc935410710ad8abe76aff426051ad6cce8257fc16d331881f74c4a4078d9fcd74c28719430b23a43a49689617037864b77adf1d3531a25bda51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haaeb27f872212631bbf0ae315d3694b924c9bd0a7f9937e0350f85632bbbcb32a2b6dcfe3079ab884590f65e6ad79c5cdbb55bb574ab91b20ea5bca96a6bd76768079c490fe2d43873d2671f59a8810c30102036ca8511cfe484f3420f308547e0f27db15854655aa4f65962c40620d67f17a0763b471ec9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5be199f870acf327a8c9c3a9e5da127d39921470641d0d8f825967b895c3571c1079e287914484e80b7281e200885d6fb372e4b440797504b4088cca852cc72f467577ca4b627d78c5bb74cc64dc515db5a89f7ca75d3ea5eba36ce74628da5535ffe59247c814bd853e4eaaf7e7a4d0a55d37f8268d47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa53e7fc0fc590228ae24696e2d9172f217cefe2c387cbb21a5a13f2341975bb99f37b7636ded9d2bc2957e5362454a33d925e7ee997378e0afda6815e7cb23068143407d0abaa4461171600880c6edb59fa15c4c286c9fe45fcdb7ebb0134ecb192fc5c144f5d7c9035ee70cceb09b902e95284fde57823;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf9675f466275799d2d0c156737cff4161c9fff3dc63cc1a3c78eacb4e1dbbc99b679fa7c6c4b3854093a98979485826ad5a469f6d92a50b51ac5b1cf12205351d59184c0605813e4861315920e77d646326fe9bfcc11c4f0fd77b98a5b053b28a7ce5b7689ec718e931d572124022e88ee280e1ae26b31c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bdeb82e9101d311a6e235bd9992bba1eb7f8f1809e135cbcab5198ee458846eaace9b78a8b76f06bb134d73dd03f87b84b7fc2ad644b7e1c868a54dca349a6f86aef474adbf070c6be3ab6479b750cb0e6f8f4d0885e3935ec212320d5966c254f1499d3b003d0a06d9759a56b996175e1a572ee1b1e17fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae77993bc105d77784d9e0668a12f01ad68ea789f986365f11c1b73ad5a7bec2bd9ddec95f3642f2e3d0edafb1ff4ffd20014c1c7bff745fc171d1fb1077fbae5223d21166d3eac470927347822a6576f8ff5dd30e6eb314cd380a26a88fd4b6f4bc07d663c36ab9f2200a2ad2cc139e28faa1064b68ef4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9ecd3cdeb03aa1ce2a00d6d3b74b0dae728fa3f3e312ff417cc1bd847fa111d5b1b3a82c44dd171c9360cf55894932b849af5af616b3eb0fd7b1c3c29848d65b35df4e3b17ae85f9e643a27c285dc5b8f9b3c6eaebf77cc8bd988d3a7cf374b2f075a8356d8544c78b5f3c40d53e760eabfb0207b3394dce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac9950a847ab223f97f63459262377f7c3aa73860db0f95c665ea76dd270d2934cb56e5bbfaf52831550f55a170f64519fa1c24859bf12e631082a105468456ec80653c556b833805d8d39970e28f52f6a1ccfee9fb9b36c0ee54e8b8fb79143a39ea889ae78afe0664fd1320470a9209cb4aebd5681543;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1086668b878c6588cdc23e09fb772ec96c4114af05e35f040e6ec66a36bca9fe5e58e9d7c7db4782b3588b735b01b41e4dab52ee8d3d9bec5b4914b77abfadf78f7e388e8e08fa52626c4d94ce16826f28c0cd6b0816fa47099fec4886868955f8245ae4c051f67cba69cfad49ac46f2cb454e2aeeb9aaa43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a48db35aee1bd20629623fea29c04e782ef7bbeae7e7c1da386adc6af1a94a788f82f853fe782eacb0b309230712dc19f8bf550c4d62622c533420f3b25a8130c158b60ddf8f8250b27f8c1574abd19648eae4fae59a94c47a51db3378b6cf91a8a5577e0955fb5554aa8beac72a64dc226fb17d68143e82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3e6d8e4f4c4f1fcb701c407a01a0173c3686964a0edff9a3e86a1bfb16286d1575e3aadec0b7f0751ea2a00ab908d400e20749eba800b0d94d82748b126a5b71bb58d6cfa0e0991036eda07f5d6be3dd530052f1fae7793647eda7eaf146479f4c0ffdb4c4a43bb0cef5c8032e517cd7e35e62c26a7f384;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h578b0d401ea800ead05d89dcbe5d82736864efe9f0cdce99b504f67b11490f96821978e5810cd192d81f367548cc2f2256264e896e2877ce66dfb7faa8e2432d39b3c07813ecae2fdaa9365a4b6546a1167907e96527fea34047aadb7f2fe176510922f4c49dddd4a29385c819cd81f1a736f44e8eda2c0b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c90d999da6f888a9a9e1724915f19b0c3fd9d76f6d2b868dae66992d8f1caa7f60784546cbcaadb9581cb8b8332e9f3c23649ce6b800da990a5c4b7bd8ade922656900fd3163f830971b213243d6470e77e48462fdbf9d549056616bf57f4572f64b712fcceead99969a721a51029001cf511ba4f0e94d3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b70be15c5e1c850f818b2cc2bcd8ae71140d9d7de4ccb9b09a322f63cf376d24c4bcf33f09d74b421365c20f15310824c1b797f75080f3ad1d091822b574313d99b2b239af0eeda93900f9abe8cca34c92b5ae28b7aec6527e3be1e6a93048f6720b9f7272734bd9154b01717ee25a466680575ee040c04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc916192994918b4677bf521979316fec2e47a122dba7ac5e1326c6494fbc52ada7ad1d7ae67fd4d32b89db6cd70aff5f3f9705d7f57f1e5b7a969926945515f8f494dada1c2d6d2a948ad9d5a0995dfceecda223f2a4a7924307adb9c8500e8c462095f17282a5d6fd7bebcd219afc604eda3bfafa113034;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he64ca067616364dcd5bdb2b9ab371ae54151e645e2fa15b5da726a9e4f68a7633db6dedc0870f16a89bb680001598be676a2147bd5aa2cdbfe4379d78f16804732b42b7655135a30d65f64da34d393740790855a120138e886ad640228f60562316d5ff869bb5a4c84893881946504b80377c1f3c16b36ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ee4fb30d1d486bc09d1ea90de5ed653af6be75931895c7eb3bfe6160b9ac486256d11838f70d1a5d0eba0f08785752fcef1bbd13db3a077274aaebaa791b6f7f6369588c67609174dae5aca05d4feabeb3c0f3f72a770e3469a985e33a91354175e64ad6724cbc650177f4b8d46293b8babd9fddbeed083;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b425d65ad4ab16685e4a6c7eeb9dbe0e064df06388ad453e97ce194bf5594ce2611aba807e6ff4441c8181fc1e904bef356448115774295ef48647e293444d3823aa0d71df0b3df5bf509e22dc1a35d2ac484d5d0e73db73378e912bd558f12c166520f1fe1c3538ac0785fa21dfe9b75de5edc7f51138bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2d05abba0cb5ec3fedc221de9608f5ecf8ec094c5bbdd737d9e484f19cbc338fbb7459c0cba879e268ed724a49c076f07062bd4dee83a9609b176640496aa6dd2e88fdb6ff059d7a176d9a9805701ac5688c11d6d4a91b27542dc5a42ce1749525b3afde3911f71efc1740760eef6908c387868967e4b4a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d8827b914510f8d916b2b03958fa62d02f91bf996755fe1c6d1bcf83539f9d60d865ae358d398a5723adbcff477ec9ada73c65e6a723f7a9b55dd652aae4c36eb5e92a11d5b33ecd8ab86ee048a0698690b2aacc561f0bacdce97409661b0b6dba7a31d4b96d99963334f0daaa1e555c96ee73e4046e177;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd265ded48f279d212a2455330e81bc6e514b70d7c57dbbb7d89aca2e0689863f631ad33a8f69b70d0c28425ecdb683affb0701f47e2c886b7ebcec69a058a370fc6bfa552b22deec1a54d06bf1e66017010ed7c3d46d24bc037c134d65b3988d28abe73db25c1233e634a57024ad507737c73fbf31eb72cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100d2e88a597747f5ab0e5cb96697ed644a7d278dcaedcc3165e97cfbd827a37670f06fac69f5bef1dbe0827fa87427c1b4bad8c2983af138e200c579d3074e2960d63e305603db820a8f70698a08278723c49c6c5982c51395f5a31c1146834d0db698214985971a6e0cede929ee6091bd5e1f1b1d74bb9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea94fc0674182a0051a249a482ac293806208108c9b119d42bcae7f878f6d062ab97d48f875e0e52592495ea99f33963fb7831a421c9e81e0df17f04736c6e7eaa09a265549469699b7880575995dfff1ea0800d8ac767a202cad78fb40d88f0197ed33d17bcc6cc5cde505a62e220dad96e44668e3a77f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbd528bded698d3eb2d6372ad905a870c52e81961bf9c5c723718743ef886ad23c70b28d6d6c481948d51db26e723963440ea4beba2a65e7435b19294f58ceaed3c39596bade79d47416998ef9fef15ea56034b3e39544c9cf74e6b6fce601071277c13fa49d1c53046364ac14ae782602cc596699f3e393;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d22c7f9d4ec5f1b973f6dd622c6bf62dfeb4d16d986b51f7f8fba4d31400763a8ee1c664bd2a6047ced11e82395dd7b6c6995c2b8e450ce7b8547bde950be423d019e6309df035ea7543a6d4ffdeb4df0cf35082257f7a3e9fd7b80f3bb096354e762c0a00eca8e0090654466f37ca46ba57b3fd173c2e20;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61acd7f7901d5cf0e4d127eca4a9bcac1f49b293b42ffd0dccbece5cd5db06a18a200cba0de9aea0809012c0098529c8086d6dc2f3c2792445eea3c3f673639f07b972917df96bd22b1387a9137a647aa8de10eeb99c04b4b6d2df7e673b0d138f37835e60302d9ebf1e8f3617b6d0c182339443773a6164;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3f71ea45a99b5a669d1276c432da173dc0264096d8e925c0e03f4aac9aa137a5e6f615084d79413ce806f72684784fd33aef99f31082b323414e5dbdb7de9bf0b83857241a3555502f046dd33c8a2894c58c0f8a08393445e9005c3972c9d1a677247a01e94544370b845c00de8b914002009572c940c38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e8cd6f8459d686e6eb60e7df4197abe7d9029a5ea5305d9bfe9731cfac4c379557bfa799315d40f56583aa9e390a9a3dc2912de5a386b920c91fa9f39aaf32d541c438adb24e755607ef7ef102fb95789362d9b652d95bca2095099ee47eb0981ff7d7b826ddc9c3088da6658ec71f8536f3e002a90d5ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haaaaa3e0a53a86cee789c4b71b106191d0cab384efc74e043f461209f9e7ca79ed65088afc645d8c4e858505215316703d6a632284f7dee798ff8cd1b347b85b344b6759d470fa611cac9b39537e2460007178e82bef3974f946d78554b85a603125a97b3cbdf0955117fa7fc51f57fa0667f3c07466415a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heaaef65eeaf78d7b3b835baaee4b8b441b13e51f3b549df460645c833c898cb6f185064a483174965f98af7be9b8c59b4f7a27b77064ed73202be0ab9ccf48febb9ecd1dd40bfbd21cd0961a558f6ca7db145e0e6b105b1367f9bfdc664477ee03ad13beeaf39d01cae30f15ce167799fa11e2cef4033c0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ba90202b464d0c57cf234256105f46fdd29b71241e16ef35348dfebe8e9d7b67bc3755604a256fb1761b34406a68613ada9ba5136e3302603f17e4851304050ff9b920d636f221492f4a7e21a4890e332d9ba6e4da68137134ddf3b5bb5b910f39963abbf24081603cb2d902dfd58de0a023f5269e35d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167b8e6dbf36345607345213807d4590651bd583a7d5bcc06347e8cdd3a7bf9ce317cfa6dc1a4c0dd13cd77544b9f96101d8cd7dbaf39fb8ac72a327d49204c2f488313776894160a11e6cf9922891bc74e74e4391e2282f64afc5504c9b78b059cb510a758363f3185488d3a1c2c0a3595a55c4538492fc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde143505c7a897794d73d5d76f1ebc31f7df4f1a6353ef3446d8c47879a9aed1c937ec20015e4b4b311c83441d9d609fb6986c52a4fe4f1f6083a1b359c5ea75956265450929803a95636831ad9c9edc3066f5530bf7f1fe038c2433e8a126c9302aa8a3cf549721d62b490a3659f8f251085a4b2c79f28e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88475415e6e20980e1a4f37a4b8514264cefe40819c7ef4c94ce6a1dcd12e5df3e68cb3b23f05080624859a22aa1c19ac3e67722e7afdfc56aa632b7eeb9ca33bfe843c3b16b031283a04c33ebd0bc4117c5f7667e6ccc3ede01440edca7ff921876c8704586a2c85bcfa9d74331547a6bb1953df001aae5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6b8280b766378fb2ec2baacf008023abc56b15baa772b2f645ad83a4bdaf490fed198e885c7e3873bfc02eddec8e9a5747f90eee9fdcf6728f3c69ef883e4fd6d4872e06bf62bcefdb879b6e1d99b9f85cf521191d5a3d99d0347f9e42b591a6ef931c06d8480db91118351506bf08d6baaef74439a9226;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2b727ebcb2fd8995c1948a23e47fda42446163976a3bae53399a376d815d7b59c6cb1839c1780ffe376a8a7937ef4438a0cef9b1adcd3698589454c63cb527b5a51c2d0e9bafe87277e4fd1409a198006ddf9ccceb3c66b38eb6e846268ca64de8b2ebfdaefe492928b56c79b0285bb266558c68a019035;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc94245925c2bfe8e86b55b71c9b091c97295f6ee5f426bdecb9fb319bde55388901901b2e92506e916de6a16ef5d6d14e24324a30d19fafe40f387fa6b0981a5d46ec480c18c004eef18c73856f2e3a8a358ef9775f33dfa8d25e19bfcd650e04423205c0204670e800f3e98434178350c9fac7b3739841;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ab903cf57551850bb578b6def61327d07c56212004bf1fa43f74be26c524d7304dad504d22945019f251f1dd76a10aaaba011d86961742c7224de6737a669b830402a6c835b502c746712aa33b4993c92f01dfb1cf7fdf03d6f0d6b90074efc758f2cc89823fab6ecac9025122273ed2ff4148068a3ad2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1953df0d383c9230eba4b3bc0503ca128858040297d3288f4c67323cd28aebac47413c10b087837c36d9d2ad3221af69225d529463024c7e1c83d220359eb21560e28ce46fb6a16f2c41925528dc156d88250807a4073f00ed7a67409294ab5f35fadac6282130752ec79010578de89b5dd899fb4d6fb3717;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157fe36918172cf94f75ae6915ab1434518ea9cd5a676d0d7818e84ae9de73d45e5661c77b4f4a89619b9d63cc352e0459bfb8c52789ab3b6b407a23cb012362751c0ce38a3f6a1fa1065415f5b591851edeec03cce5313deaef5f2456575c64a1e65f92432601776b616c16e0cefd192b9d91b30ea2b2eed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ee680081470f550cebe8cada17f72e2a12fcba015c2c7cd76d0954527320fe43c9acfecf9f2b7a94ce53e7f22eeb6a902788ae2825310289279c1575b2b12b0cedc54743de3bfdc6c2be3dab3217aab6bf527027ea98c1ec7138c8edd88208d15b2694f7222cb31318f577cf06ba1c33b41755a76c47248;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0012d0d56cb78cc4b535a06c1cbcbfbcd2359a576b688515b685b05736211aafa1bf5697d9cfbda89f57bb195038949ae757c8ed949a9d12cb49f738af5cdd269b305cce2edbdebbb7599343f6eb7264ac8a3f21816bd9f0a76e292d93302230d38b982d92274a9981574f10cf547cf7146078ead61bb9e;
        #1
        $finish();
    end
endmodule
