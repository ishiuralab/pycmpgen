module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    compressor_CLA486_12 compressor_CLA486_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA486_12(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [1:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[1], 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [1:0] dst20);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [85:0] stage1_0;
   wire [154:0] stage1_1;
   wire [197:0] stage1_2;
   wire [195:0] stage1_3;
   wire [240:0] stage1_4;
   wire [229:0] stage1_5;
   wire [169:0] stage1_6;
   wire [161:0] stage1_7;
   wire [238:0] stage1_8;
   wire [240:0] stage1_9;
   wire [179:0] stage1_10;
   wire [170:0] stage1_11;
   wire [156:0] stage1_12;
   wire [78:0] stage1_13;
   wire [30:0] stage2_0;
   wire [57:0] stage2_1;
   wire [53:0] stage2_2;
   wire [83:0] stage2_3;
   wire [88:0] stage2_4;
   wire [74:0] stage2_5;
   wire [97:0] stage2_6;
   wire [88:0] stage2_7;
   wire [70:0] stage2_8;
   wire [91:0] stage2_9;
   wire [98:0] stage2_10;
   wire [81:0] stage2_11;
   wire [111:0] stage2_12;
   wire [51:0] stage2_13;
   wire [26:0] stage2_14;
   wire [11:0] stage2_15;
   wire [13:0] stage3_0;
   wire [25:0] stage3_1;
   wire [16:0] stage3_2;
   wire [24:0] stage3_3;
   wire [33:0] stage3_4;
   wire [31:0] stage3_5;
   wire [44:0] stage3_6;
   wire [37:0] stage3_7;
   wire [30:0] stage3_8;
   wire [42:0] stage3_9;
   wire [37:0] stage3_10;
   wire [53:0] stage3_11;
   wire [46:0] stage3_12;
   wire [33:0] stage3_13;
   wire [25:0] stage3_14;
   wire [17:0] stage3_15;
   wire [4:0] stage3_16;
   wire [0:0] stage3_17;
   wire [8:0] stage4_0;
   wire [11:0] stage4_1;
   wire [6:0] stage4_2;
   wire [6:0] stage4_3;
   wire [12:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [18:0] stage4_7;
   wire [12:0] stage4_8;
   wire [16:0] stage4_9;
   wire [18:0] stage4_10;
   wire [15:0] stage4_11;
   wire [17:0] stage4_12;
   wire [22:0] stage4_13;
   wire [16:0] stage4_14;
   wire [7:0] stage4_15;
   wire [11:0] stage4_16;
   wire [3:0] stage4_17;
   wire [6:0] stage5_0;
   wire [6:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [3:0] stage5_4;
   wire [4:0] stage5_5;
   wire [6:0] stage5_6;
   wire [5:0] stage5_7;
   wire [11:0] stage5_8;
   wire [6:0] stage5_9;
   wire [7:0] stage5_10;
   wire [7:0] stage5_11;
   wire [6:0] stage5_12;
   wire [10:0] stage5_13;
   wire [7:0] stage5_14;
   wire [6:0] stage5_15;
   wire [3:0] stage5_16;
   wire [6:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage6_0;
   wire [6:0] stage6_1;
   wire [4:0] stage6_2;
   wire [6:0] stage6_3;
   wire [3:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [6:0] stage6_8;
   wire [2:0] stage6_9;
   wire [3:0] stage6_10;
   wire [3:0] stage6_11;
   wire [1:0] stage6_12;
   wire [5:0] stage6_13;
   wire [4:0] stage6_14;
   wire [1:0] stage6_15;
   wire [2:0] stage6_16;
   wire [3:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;
   wire [0:0] stage6_20;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [0:0] stage7_19;
   wire [1:0] stage7_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[10]},
      {stage0_3[20]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[11]},
      {stage0_3[21]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[12]},
      {stage0_3[22]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[13]},
      {stage0_3[23]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[14]},
      {stage0_3[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[15]},
      {stage0_3[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[16]},
      {stage0_3[26]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc207_4 gpc17 (
      {stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_2[17], stage0_2[18]},
      {stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[46],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[47],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[48],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[49],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[50],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[51],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[52],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[53],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[54],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[55],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[56],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[57],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[58],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[59],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[60],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[61],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[62],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[63],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[64],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[65],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[66],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[67],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389]},
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage1_4[68],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395]},
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage1_4[69],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401]},
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage1_4[70],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage1_4[71],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413]},
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354]},
      {stage1_4[72],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419]},
      {stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360]},
      {stage1_4[73],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425]},
      {stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366]},
      {stage1_4[74],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431]},
      {stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372]},
      {stage1_4[75],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage1_4[76],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384]},
      {stage1_4[77],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448], stage0_0[449]},
      {stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390]},
      {stage1_4[78],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454], stage0_0[455]},
      {stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396]},
      {stage1_4[79],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461]},
      {stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage1_4[80],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage1_4[81],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472], stage0_0[473]},
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage1_4[82],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478], stage0_0[479]},
      {stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage1_4[83],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484], stage0_0[485]},
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426]},
      {stage1_4[84],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[0],stage1_4[85],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[1],stage1_4[86],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[2],stage1_4[87],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[3],stage1_4[88],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[4],stage1_4[89],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[5],stage1_4[90],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[6],stage1_4[91],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[7],stage1_4[92],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[8],stage1_4[93],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[9],stage1_4[94],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[10],stage1_4[95],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[11],stage1_4[96],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[12],stage1_4[97],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[13],stage1_4[98],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[14],stage1_4[99],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[15],stage1_4[100],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[16],stage1_4[101],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[17],stage1_4[102],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[18],stage1_4[103],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[19],stage1_4[104],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[20],stage1_4[105],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[21],stage1_4[106],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[22],stage1_4[107],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[23],stage1_4[108],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[24],stage1_4[109],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[25],stage1_4[110],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[26],stage1_4[111],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[27],stage1_4[112],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[28],stage1_4[113],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[29],stage1_4[114],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[30],stage1_4[115],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[31],stage1_4[116],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224]},
      {stage1_5[32],stage1_4[117],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage1_5[33],stage1_4[118],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage1_5[34],stage1_4[119],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage1_5[35],stage1_4[120],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248]},
      {stage1_5[36],stage1_4[121],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254]},
      {stage1_5[37],stage1_4[122],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260]},
      {stage1_5[38],stage1_4[123],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage1_5[39],stage1_4[124],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272]},
      {stage1_5[40],stage1_4[125],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278]},
      {stage1_5[41],stage1_4[126],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284]},
      {stage1_5[42],stage1_4[127],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage1_5[43],stage1_4[128],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage1_5[44],stage1_4[129],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302]},
      {stage1_5[45],stage1_4[130],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage1_5[46],stage1_4[131],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314]},
      {stage1_5[47],stage1_4[132],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage1_5[48],stage1_4[133],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage1_5[49],stage1_4[134],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332]},
      {stage1_5[50],stage1_4[135],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage1_5[51],stage1_4[136],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344]},
      {stage1_5[52],stage1_4[137],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage1_5[53],stage1_4[138],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage1_5[54],stage1_4[139],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362]},
      {stage1_5[55],stage1_4[140],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage1_5[56],stage1_4[141],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374]},
      {stage1_5[57],stage1_4[142],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage1_5[58],stage1_4[143],stage1_3[144],stage1_2[144],stage1_1[144]}
   );
   gpc606_5 gpc145 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385], stage0_3[386]},
      {stage1_5[59],stage1_4[144],stage1_3[145],stage1_2[145],stage1_1[145]}
   );
   gpc606_5 gpc146 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392]},
      {stage1_5[60],stage1_4[145],stage1_3[146],stage1_2[146],stage1_1[146]}
   );
   gpc606_5 gpc147 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[393], stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage1_5[61],stage1_4[146],stage1_3[147],stage1_2[147],stage1_1[147]}
   );
   gpc606_5 gpc148 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404]},
      {stage1_5[62],stage1_4[147],stage1_3[148],stage1_2[148],stage1_1[148]}
   );
   gpc606_5 gpc149 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage1_5[63],stage1_4[148],stage1_3[149],stage1_2[149],stage1_1[149]}
   );
   gpc606_5 gpc150 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415], stage0_3[416]},
      {stage1_5[64],stage1_4[149],stage1_3[150],stage1_2[150],stage1_1[150]}
   );
   gpc606_5 gpc151 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422]},
      {stage1_5[65],stage1_4[150],stage1_3[151],stage1_2[151],stage1_1[151]}
   );
   gpc606_5 gpc152 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[423], stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage1_5[66],stage1_4[151],stage1_3[152],stage1_2[152],stage1_1[152]}
   );
   gpc606_5 gpc153 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434]},
      {stage1_5[67],stage1_4[152],stage1_3[153],stage1_2[153],stage1_1[153]}
   );
   gpc606_5 gpc154 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage1_5[68],stage1_4[153],stage1_3[154],stage1_2[154],stage1_1[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_3[441]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[69],stage1_4[154],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436]},
      {stage0_3[442]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[70],stage1_4[155],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441]},
      {stage0_3[443]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[71],stage1_4[156],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446]},
      {stage0_3[444]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[72],stage1_4[157],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[73],stage1_4[158],stage1_3[159]}
   );
   gpc606_5 gpc160 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[74],stage1_4[159]}
   );
   gpc606_5 gpc161 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[75],stage1_4[160]}
   );
   gpc606_5 gpc162 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[76],stage1_4[161]}
   );
   gpc606_5 gpc163 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[77],stage1_4[162]}
   );
   gpc606_5 gpc164 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[78],stage1_4[163]}
   );
   gpc606_5 gpc165 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[79],stage1_4[164]}
   );
   gpc606_5 gpc166 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[80],stage1_4[165]}
   );
   gpc606_5 gpc167 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[81],stage1_4[166]}
   );
   gpc606_5 gpc168 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[82],stage1_4[167]}
   );
   gpc606_5 gpc169 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[83],stage1_4[168]}
   );
   gpc606_5 gpc170 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[84],stage1_4[169]}
   );
   gpc606_5 gpc171 (
      {stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[85],stage1_4[170]}
   );
   gpc606_5 gpc172 (
      {stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[86],stage1_4[171]}
   );
   gpc606_5 gpc173 (
      {stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[87],stage1_4[172]}
   );
   gpc606_5 gpc174 (
      {stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[88],stage1_4[173]}
   );
   gpc606_5 gpc175 (
      {stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc176 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc177 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[18],stage1_6[22],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc178 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[19],stage1_6[23],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc179 (
      {stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[20],stage1_6[24],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc180 (
      {stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[21],stage1_6[25],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc181 (
      {stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[22],stage1_6[26],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc182 (
      {stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[23],stage1_6[27],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc183 (
      {stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[24],stage1_6[28],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc184 (
      {stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[25],stage1_6[29],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc185 (
      {stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[26],stage1_6[30],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc186 (
      {stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[27],stage1_6[31],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc187 (
      {stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[28],stage1_6[32],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc188 (
      {stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[29],stage1_6[33],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc189 (
      {stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[30],stage1_6[34],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc190 (
      {stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[31],stage1_6[35],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc191 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[32],stage1_6[36],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc192 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[33],stage1_6[37],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc193 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[34],stage1_6[38],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc194 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[35],stage1_6[39],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc195 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[36],stage1_6[40],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc196 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[37],stage1_6[41],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc197 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[38],stage1_6[42],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc198 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[39],stage1_6[43],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc199 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[40],stage1_6[44],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc200 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[41],stage1_6[45],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc201 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[42],stage1_6[46],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc202 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[43],stage1_6[47],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc203 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[44],stage1_6[48],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc204 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[45],stage1_6[49],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc205 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[46],stage1_6[50],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc206 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[47],stage1_6[51],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc207 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[48],stage1_6[52],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc208 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[49],stage1_6[53],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc209 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[50],stage1_6[54],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc210 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[51],stage1_6[55],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc211 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[52],stage1_6[56],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc212 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[53],stage1_6[57],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc213 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[54],stage1_6[58],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc214 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[55],stage1_6[59],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc215 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[56],stage1_6[60],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc216 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[57],stage1_6[61],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc217 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[58],stage1_6[62],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc218 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[59],stage1_6[63],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc219 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[60],stage1_6[64],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc220 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[61],stage1_6[65],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc221 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[62],stage1_6[66],stage1_5[135],stage1_4[220]}
   );
   gpc606_5 gpc222 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[63],stage1_6[67],stage1_5[136],stage1_4[221]}
   );
   gpc606_5 gpc223 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[64],stage1_6[68],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc224 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[65],stage1_6[69],stage1_5[138],stage1_4[223]}
   );
   gpc606_5 gpc225 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[66],stage1_6[70],stage1_5[139],stage1_4[224]}
   );
   gpc606_5 gpc226 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[67],stage1_6[71],stage1_5[140],stage1_4[225]}
   );
   gpc606_5 gpc227 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[68],stage1_6[72],stage1_5[141],stage1_4[226]}
   );
   gpc606_5 gpc228 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[69],stage1_6[73],stage1_5[142],stage1_4[227]}
   );
   gpc606_5 gpc229 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[70],stage1_6[74],stage1_5[143],stage1_4[228]}
   );
   gpc606_5 gpc230 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[71],stage1_6[75],stage1_5[144],stage1_4[229]}
   );
   gpc615_5 gpc231 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455]},
      {stage0_5[6]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[72],stage1_6[76],stage1_5[145],stage1_4[230]}
   );
   gpc615_5 gpc232 (
      {stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_5[7]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[73],stage1_6[77],stage1_5[146],stage1_4[231]}
   );
   gpc615_5 gpc233 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_5[8]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[74],stage1_6[78],stage1_5[147],stage1_4[232]}
   );
   gpc615_5 gpc234 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470]},
      {stage0_5[9]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[75],stage1_6[79],stage1_5[148],stage1_4[233]}
   );
   gpc615_5 gpc235 (
      {stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_5[10]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[76],stage1_6[80],stage1_5[149],stage1_4[234]}
   );
   gpc615_5 gpc236 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[11]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[77],stage1_6[81],stage1_5[150],stage1_4[235]}
   );
   gpc606_5 gpc237 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[77],stage1_7[78],stage1_6[82],stage1_5[151]}
   );
   gpc606_5 gpc238 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[78],stage1_7[79],stage1_6[83],stage1_5[152]}
   );
   gpc606_5 gpc239 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[79],stage1_7[80],stage1_6[84],stage1_5[153]}
   );
   gpc606_5 gpc240 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[80],stage1_7[81],stage1_6[85],stage1_5[154]}
   );
   gpc606_5 gpc241 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[81],stage1_7[82],stage1_6[86],stage1_5[155]}
   );
   gpc606_5 gpc242 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[82],stage1_7[83],stage1_6[87],stage1_5[156]}
   );
   gpc606_5 gpc243 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[83],stage1_7[84],stage1_6[88],stage1_5[157]}
   );
   gpc606_5 gpc244 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[84],stage1_7[85],stage1_6[89],stage1_5[158]}
   );
   gpc606_5 gpc245 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[85],stage1_7[86],stage1_6[90],stage1_5[159]}
   );
   gpc606_5 gpc246 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[86],stage1_7[87],stage1_6[91],stage1_5[160]}
   );
   gpc606_5 gpc247 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[87],stage1_7[88],stage1_6[92],stage1_5[161]}
   );
   gpc606_5 gpc248 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[88],stage1_7[89],stage1_6[93],stage1_5[162]}
   );
   gpc606_5 gpc249 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[89],stage1_7[90],stage1_6[94],stage1_5[163]}
   );
   gpc606_5 gpc250 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[90],stage1_7[91],stage1_6[95],stage1_5[164]}
   );
   gpc606_5 gpc251 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[91],stage1_7[92],stage1_6[96],stage1_5[165]}
   );
   gpc606_5 gpc252 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[92],stage1_7[93],stage1_6[97],stage1_5[166]}
   );
   gpc606_5 gpc253 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[93],stage1_7[94],stage1_6[98],stage1_5[167]}
   );
   gpc606_5 gpc254 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[94],stage1_7[95],stage1_6[99],stage1_5[168]}
   );
   gpc606_5 gpc255 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[95],stage1_7[96],stage1_6[100],stage1_5[169]}
   );
   gpc606_5 gpc256 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[96],stage1_7[97],stage1_6[101],stage1_5[170]}
   );
   gpc606_5 gpc257 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[97],stage1_7[98],stage1_6[102],stage1_5[171]}
   );
   gpc606_5 gpc258 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[98],stage1_7[99],stage1_6[103],stage1_5[172]}
   );
   gpc606_5 gpc259 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[99],stage1_7[100],stage1_6[104],stage1_5[173]}
   );
   gpc606_5 gpc260 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[100],stage1_7[101],stage1_6[105],stage1_5[174]}
   );
   gpc606_5 gpc261 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[101],stage1_7[102],stage1_6[106],stage1_5[175]}
   );
   gpc606_5 gpc262 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[102],stage1_7[103],stage1_6[107],stage1_5[176]}
   );
   gpc606_5 gpc263 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[103],stage1_7[104],stage1_6[108],stage1_5[177]}
   );
   gpc606_5 gpc264 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[104],stage1_7[105],stage1_6[109],stage1_5[178]}
   );
   gpc606_5 gpc265 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[105],stage1_7[106],stage1_6[110],stage1_5[179]}
   );
   gpc606_5 gpc266 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[106],stage1_7[107],stage1_6[111],stage1_5[180]}
   );
   gpc606_5 gpc267 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[107],stage1_7[108],stage1_6[112],stage1_5[181]}
   );
   gpc606_5 gpc268 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[108],stage1_7[109],stage1_6[113],stage1_5[182]}
   );
   gpc606_5 gpc269 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[109],stage1_7[110],stage1_6[114],stage1_5[183]}
   );
   gpc606_5 gpc270 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[110],stage1_7[111],stage1_6[115],stage1_5[184]}
   );
   gpc606_5 gpc271 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[111],stage1_7[112],stage1_6[116],stage1_5[185]}
   );
   gpc606_5 gpc272 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[112],stage1_7[113],stage1_6[117],stage1_5[186]}
   );
   gpc606_5 gpc273 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[113],stage1_7[114],stage1_6[118],stage1_5[187]}
   );
   gpc606_5 gpc274 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[114],stage1_7[115],stage1_6[119],stage1_5[188]}
   );
   gpc606_5 gpc275 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[115],stage1_7[116],stage1_6[120],stage1_5[189]}
   );
   gpc606_5 gpc276 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[116],stage1_7[117],stage1_6[121],stage1_5[190]}
   );
   gpc606_5 gpc277 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[117],stage1_7[118],stage1_6[122],stage1_5[191]}
   );
   gpc606_5 gpc278 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[118],stage1_7[119],stage1_6[123],stage1_5[192]}
   );
   gpc606_5 gpc279 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[119],stage1_7[120],stage1_6[124],stage1_5[193]}
   );
   gpc606_5 gpc280 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[120],stage1_7[121],stage1_6[125],stage1_5[194]}
   );
   gpc606_5 gpc281 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[121],stage1_7[122],stage1_6[126],stage1_5[195]}
   );
   gpc606_5 gpc282 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[122],stage1_7[123],stage1_6[127],stage1_5[196]}
   );
   gpc606_5 gpc283 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[123],stage1_7[124],stage1_6[128],stage1_5[197]}
   );
   gpc606_5 gpc284 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[124],stage1_7[125],stage1_6[129],stage1_5[198]}
   );
   gpc606_5 gpc285 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[125],stage1_7[126],stage1_6[130],stage1_5[199]}
   );
   gpc606_5 gpc286 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[126],stage1_7[127],stage1_6[131],stage1_5[200]}
   );
   gpc606_5 gpc287 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[127],stage1_7[128],stage1_6[132],stage1_5[201]}
   );
   gpc606_5 gpc288 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[128],stage1_7[129],stage1_6[133],stage1_5[202]}
   );
   gpc606_5 gpc289 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[129],stage1_7[130],stage1_6[134],stage1_5[203]}
   );
   gpc606_5 gpc290 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[130],stage1_7[131],stage1_6[135],stage1_5[204]}
   );
   gpc606_5 gpc291 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[131],stage1_7[132],stage1_6[136],stage1_5[205]}
   );
   gpc606_5 gpc292 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[132],stage1_7[133],stage1_6[137],stage1_5[206]}
   );
   gpc606_5 gpc293 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[133],stage1_7[134],stage1_6[138],stage1_5[207]}
   );
   gpc606_5 gpc294 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[134],stage1_7[135],stage1_6[139],stage1_5[208]}
   );
   gpc606_5 gpc295 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[135],stage1_7[136],stage1_6[140],stage1_5[209]}
   );
   gpc606_5 gpc296 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[136],stage1_7[137],stage1_6[141],stage1_5[210]}
   );
   gpc606_5 gpc297 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[137],stage1_7[138],stage1_6[142],stage1_5[211]}
   );
   gpc606_5 gpc298 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[138],stage1_7[139],stage1_6[143],stage1_5[212]}
   );
   gpc606_5 gpc299 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376], stage0_7[377]},
      {stage1_9[62],stage1_8[139],stage1_7[140],stage1_6[144],stage1_5[213]}
   );
   gpc606_5 gpc300 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383]},
      {stage1_9[63],stage1_8[140],stage1_7[141],stage1_6[145],stage1_5[214]}
   );
   gpc606_5 gpc301 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage1_9[64],stage1_8[141],stage1_7[142],stage1_6[146],stage1_5[215]}
   );
   gpc606_5 gpc302 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage1_9[65],stage1_8[142],stage1_7[143],stage1_6[147],stage1_5[216]}
   );
   gpc606_5 gpc303 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage1_9[66],stage1_8[143],stage1_7[144],stage1_6[148],stage1_5[217]}
   );
   gpc606_5 gpc304 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406], stage0_7[407]},
      {stage1_9[67],stage1_8[144],stage1_7[145],stage1_6[149],stage1_5[218]}
   );
   gpc606_5 gpc305 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413]},
      {stage1_9[68],stage1_8[145],stage1_7[146],stage1_6[150],stage1_5[219]}
   );
   gpc606_5 gpc306 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage1_9[69],stage1_8[146],stage1_7[147],stage1_6[151],stage1_5[220]}
   );
   gpc606_5 gpc307 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage1_9[70],stage1_8[147],stage1_7[148],stage1_6[152],stage1_5[221]}
   );
   gpc606_5 gpc308 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage1_9[71],stage1_8[148],stage1_7[149],stage1_6[153],stage1_5[222]}
   );
   gpc606_5 gpc309 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436], stage0_7[437]},
      {stage1_9[72],stage1_8[149],stage1_7[150],stage1_6[154],stage1_5[223]}
   );
   gpc606_5 gpc310 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442], stage0_7[443]},
      {stage1_9[73],stage1_8[150],stage1_7[151],stage1_6[155],stage1_5[224]}
   );
   gpc606_5 gpc311 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448], stage0_7[449]},
      {stage1_9[74],stage1_8[151],stage1_7[152],stage1_6[156],stage1_5[225]}
   );
   gpc606_5 gpc312 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455]},
      {stage1_9[75],stage1_8[152],stage1_7[153],stage1_6[157],stage1_5[226]}
   );
   gpc606_5 gpc313 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage1_9[76],stage1_8[153],stage1_7[154],stage1_6[158],stage1_5[227]}
   );
   gpc606_5 gpc314 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466], stage0_7[467]},
      {stage1_9[77],stage1_8[154],stage1_7[155],stage1_6[159],stage1_5[228]}
   );
   gpc606_5 gpc315 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471], stage0_7[472], stage0_7[473]},
      {stage1_9[78],stage1_8[155],stage1_7[156],stage1_6[160],stage1_5[229]}
   );
   gpc606_5 gpc316 (
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[79],stage1_8[156],stage1_7[157],stage1_6[161]}
   );
   gpc606_5 gpc317 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[80],stage1_8[157],stage1_7[158],stage1_6[162]}
   );
   gpc606_5 gpc318 (
      {stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[81],stage1_8[158],stage1_7[159],stage1_6[163]}
   );
   gpc606_5 gpc319 (
      {stage0_7[474], stage0_7[475], stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[82],stage1_8[159],stage1_7[160]}
   );
   gpc606_5 gpc320 (
      {stage0_7[480], stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[83],stage1_8[160],stage1_7[161]}
   );
   gpc606_5 gpc321 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[84],stage1_8[161]}
   );
   gpc606_5 gpc322 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[85],stage1_8[162]}
   );
   gpc606_5 gpc323 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[86],stage1_8[163]}
   );
   gpc606_5 gpc324 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[87],stage1_8[164]}
   );
   gpc606_5 gpc325 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[88],stage1_8[165]}
   );
   gpc606_5 gpc326 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[89],stage1_8[166]}
   );
   gpc606_5 gpc327 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[90],stage1_8[167]}
   );
   gpc606_5 gpc328 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[91],stage1_8[168]}
   );
   gpc606_5 gpc329 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[92],stage1_8[169]}
   );
   gpc606_5 gpc330 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[14],stage1_9[93],stage1_8[170]}
   );
   gpc606_5 gpc331 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[15],stage1_9[94],stage1_8[171]}
   );
   gpc606_5 gpc332 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[16],stage1_9[95],stage1_8[172]}
   );
   gpc606_5 gpc333 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[17],stage1_9[96],stage1_8[173]}
   );
   gpc606_5 gpc334 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[18],stage1_9[97],stage1_8[174]}
   );
   gpc606_5 gpc335 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[19],stage1_9[98],stage1_8[175]}
   );
   gpc606_5 gpc336 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[17],stage1_10[20],stage1_9[99],stage1_8[176]}
   );
   gpc606_5 gpc337 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[18],stage1_10[21],stage1_9[100],stage1_8[177]}
   );
   gpc606_5 gpc338 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[19],stage1_10[22],stage1_9[101],stage1_8[178]}
   );
   gpc606_5 gpc339 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[20],stage1_10[23],stage1_9[102],stage1_8[179]}
   );
   gpc606_5 gpc340 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[21],stage1_10[24],stage1_9[103],stage1_8[180]}
   );
   gpc606_5 gpc341 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[22],stage1_10[25],stage1_9[104],stage1_8[181]}
   );
   gpc606_5 gpc342 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[23],stage1_10[26],stage1_9[105],stage1_8[182]}
   );
   gpc606_5 gpc343 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[24],stage1_10[27],stage1_9[106],stage1_8[183]}
   );
   gpc606_5 gpc344 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[25],stage1_10[28],stage1_9[107],stage1_8[184]}
   );
   gpc606_5 gpc345 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[26],stage1_10[29],stage1_9[108],stage1_8[185]}
   );
   gpc606_5 gpc346 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[27],stage1_10[30],stage1_9[109],stage1_8[186]}
   );
   gpc606_5 gpc347 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[28],stage1_10[31],stage1_9[110],stage1_8[187]}
   );
   gpc606_5 gpc348 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[29],stage1_10[32],stage1_9[111],stage1_8[188]}
   );
   gpc606_5 gpc349 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[30],stage1_10[33],stage1_9[112],stage1_8[189]}
   );
   gpc606_5 gpc350 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[31],stage1_10[34],stage1_9[113],stage1_8[190]}
   );
   gpc606_5 gpc351 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[32],stage1_10[35],stage1_9[114],stage1_8[191]}
   );
   gpc606_5 gpc352 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[33],stage1_10[36],stage1_9[115],stage1_8[192]}
   );
   gpc606_5 gpc353 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[34],stage1_10[37],stage1_9[116],stage1_8[193]}
   );
   gpc606_5 gpc354 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[35],stage1_10[38],stage1_9[117],stage1_8[194]}
   );
   gpc606_5 gpc355 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[36],stage1_10[39],stage1_9[118],stage1_8[195]}
   );
   gpc606_5 gpc356 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[37],stage1_10[40],stage1_9[119],stage1_8[196]}
   );
   gpc606_5 gpc357 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[38],stage1_10[41],stage1_9[120],stage1_8[197]}
   );
   gpc606_5 gpc358 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[39],stage1_10[42],stage1_9[121],stage1_8[198]}
   );
   gpc606_5 gpc359 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[40],stage1_10[43],stage1_9[122],stage1_8[199]}
   );
   gpc606_5 gpc360 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[41],stage1_10[44],stage1_9[123],stage1_8[200]}
   );
   gpc606_5 gpc361 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[42],stage1_10[45],stage1_9[124],stage1_8[201]}
   );
   gpc606_5 gpc362 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[43],stage1_10[46],stage1_9[125],stage1_8[202]}
   );
   gpc606_5 gpc363 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[44],stage1_10[47],stage1_9[126],stage1_8[203]}
   );
   gpc606_5 gpc364 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[45],stage1_10[48],stage1_9[127],stage1_8[204]}
   );
   gpc606_5 gpc365 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[46],stage1_10[49],stage1_9[128],stage1_8[205]}
   );
   gpc606_5 gpc366 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[47],stage1_10[50],stage1_9[129],stage1_8[206]}
   );
   gpc606_5 gpc367 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[48],stage1_10[51],stage1_9[130],stage1_8[207]}
   );
   gpc606_5 gpc368 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[49],stage1_10[52],stage1_9[131],stage1_8[208]}
   );
   gpc606_5 gpc369 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[50],stage1_10[53],stage1_9[132],stage1_8[209]}
   );
   gpc606_5 gpc370 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[51],stage1_10[54],stage1_9[133],stage1_8[210]}
   );
   gpc606_5 gpc371 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[52],stage1_10[55],stage1_9[134],stage1_8[211]}
   );
   gpc606_5 gpc372 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[53],stage1_10[56],stage1_9[135],stage1_8[212]}
   );
   gpc606_5 gpc373 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[54],stage1_10[57],stage1_9[136],stage1_8[213]}
   );
   gpc606_5 gpc374 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[55],stage1_10[58],stage1_9[137],stage1_8[214]}
   );
   gpc606_5 gpc375 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[56],stage1_10[59],stage1_9[138],stage1_8[215]}
   );
   gpc606_5 gpc376 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[57],stage1_10[60],stage1_9[139],stage1_8[216]}
   );
   gpc606_5 gpc377 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[58],stage1_10[61],stage1_9[140],stage1_8[217]}
   );
   gpc606_5 gpc378 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[59],stage1_10[62],stage1_9[141],stage1_8[218]}
   );
   gpc606_5 gpc379 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[60],stage1_10[63],stage1_9[142],stage1_8[219]}
   );
   gpc606_5 gpc380 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[61],stage1_10[64],stage1_9[143],stage1_8[220]}
   );
   gpc606_5 gpc381 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[62],stage1_10[65],stage1_9[144],stage1_8[221]}
   );
   gpc606_5 gpc382 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[63],stage1_10[66],stage1_9[145],stage1_8[222]}
   );
   gpc606_5 gpc383 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[64],stage1_10[67],stage1_9[146],stage1_8[223]}
   );
   gpc606_5 gpc384 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[65],stage1_10[68],stage1_9[147],stage1_8[224]}
   );
   gpc606_5 gpc385 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[66],stage1_10[69],stage1_9[148],stage1_8[225]}
   );
   gpc606_5 gpc386 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[67],stage1_10[70],stage1_9[149],stage1_8[226]}
   );
   gpc606_5 gpc387 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[68],stage1_10[71],stage1_9[150],stage1_8[227]}
   );
   gpc606_5 gpc388 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[69],stage1_10[72],stage1_9[151],stage1_8[228]}
   );
   gpc606_5 gpc389 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[70],stage1_10[73],stage1_9[152],stage1_8[229]}
   );
   gpc606_5 gpc390 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[71],stage1_10[74],stage1_9[153],stage1_8[230]}
   );
   gpc606_5 gpc391 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[72],stage1_10[75],stage1_9[154],stage1_8[231]}
   );
   gpc606_5 gpc392 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[73],stage1_10[76],stage1_9[155],stage1_8[232]}
   );
   gpc606_5 gpc393 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437]},
      {stage1_12[72],stage1_11[74],stage1_10[77],stage1_9[156],stage1_8[233]}
   );
   gpc606_5 gpc394 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage1_12[73],stage1_11[75],stage1_10[78],stage1_9[157],stage1_8[234]}
   );
   gpc606_5 gpc395 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage1_12[74],stage1_11[76],stage1_10[79],stage1_9[158],stage1_8[235]}
   );
   gpc606_5 gpc396 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455]},
      {stage1_12[75],stage1_11[77],stage1_10[80],stage1_9[159],stage1_8[236]}
   );
   gpc606_5 gpc397 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage1_12[76],stage1_11[78],stage1_10[81],stage1_9[160],stage1_8[237]}
   );
   gpc606_5 gpc398 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467]},
      {stage1_12[77],stage1_11[79],stage1_10[82],stage1_9[161],stage1_8[238]}
   );
   gpc606_5 gpc399 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[78],stage1_11[80],stage1_10[83],stage1_9[162]}
   );
   gpc606_5 gpc400 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[79],stage1_11[81],stage1_10[84],stage1_9[163]}
   );
   gpc606_5 gpc401 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[80],stage1_11[82],stage1_10[85],stage1_9[164]}
   );
   gpc606_5 gpc402 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[81],stage1_11[83],stage1_10[86],stage1_9[165]}
   );
   gpc606_5 gpc403 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[82],stage1_11[84],stage1_10[87],stage1_9[166]}
   );
   gpc606_5 gpc404 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[83],stage1_11[85],stage1_10[88],stage1_9[167]}
   );
   gpc606_5 gpc405 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[84],stage1_11[86],stage1_10[89],stage1_9[168]}
   );
   gpc606_5 gpc406 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[85],stage1_11[87],stage1_10[90],stage1_9[169]}
   );
   gpc606_5 gpc407 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[86],stage1_11[88],stage1_10[91],stage1_9[170]}
   );
   gpc606_5 gpc408 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[87],stage1_11[89],stage1_10[92],stage1_9[171]}
   );
   gpc606_5 gpc409 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[88],stage1_11[90],stage1_10[93],stage1_9[172]}
   );
   gpc606_5 gpc410 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[89],stage1_11[91],stage1_10[94],stage1_9[173]}
   );
   gpc606_5 gpc411 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[90],stage1_11[92],stage1_10[95],stage1_9[174]}
   );
   gpc606_5 gpc412 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[91],stage1_11[93],stage1_10[96],stage1_9[175]}
   );
   gpc606_5 gpc413 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[92],stage1_11[94],stage1_10[97],stage1_9[176]}
   );
   gpc606_5 gpc414 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[93],stage1_11[95],stage1_10[98],stage1_9[177]}
   );
   gpc606_5 gpc415 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[94],stage1_11[96],stage1_10[99],stage1_9[178]}
   );
   gpc606_5 gpc416 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[95],stage1_11[97],stage1_10[100],stage1_9[179]}
   );
   gpc606_5 gpc417 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[96],stage1_11[98],stage1_10[101],stage1_9[180]}
   );
   gpc606_5 gpc418 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[97],stage1_11[99],stage1_10[102],stage1_9[181]}
   );
   gpc606_5 gpc419 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[98],stage1_11[100],stage1_10[103],stage1_9[182]}
   );
   gpc606_5 gpc420 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[99],stage1_11[101],stage1_10[104],stage1_9[183]}
   );
   gpc606_5 gpc421 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[100],stage1_11[102],stage1_10[105],stage1_9[184]}
   );
   gpc606_5 gpc422 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[101],stage1_11[103],stage1_10[106],stage1_9[185]}
   );
   gpc606_5 gpc423 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[102],stage1_11[104],stage1_10[107],stage1_9[186]}
   );
   gpc606_5 gpc424 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[103],stage1_11[105],stage1_10[108],stage1_9[187]}
   );
   gpc606_5 gpc425 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[104],stage1_11[106],stage1_10[109],stage1_9[188]}
   );
   gpc606_5 gpc426 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[105],stage1_11[107],stage1_10[110],stage1_9[189]}
   );
   gpc606_5 gpc427 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[106],stage1_11[108],stage1_10[111],stage1_9[190]}
   );
   gpc606_5 gpc428 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[107],stage1_11[109],stage1_10[112],stage1_9[191]}
   );
   gpc606_5 gpc429 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[108],stage1_11[110],stage1_10[113],stage1_9[192]}
   );
   gpc606_5 gpc430 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[109],stage1_11[111],stage1_10[114],stage1_9[193]}
   );
   gpc606_5 gpc431 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[110],stage1_11[112],stage1_10[115],stage1_9[194]}
   );
   gpc606_5 gpc432 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[111],stage1_11[113],stage1_10[116],stage1_9[195]}
   );
   gpc606_5 gpc433 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[112],stage1_11[114],stage1_10[117],stage1_9[196]}
   );
   gpc606_5 gpc434 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[113],stage1_11[115],stage1_10[118],stage1_9[197]}
   );
   gpc606_5 gpc435 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[114],stage1_11[116],stage1_10[119],stage1_9[198]}
   );
   gpc606_5 gpc436 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[115],stage1_11[117],stage1_10[120],stage1_9[199]}
   );
   gpc606_5 gpc437 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[116],stage1_11[118],stage1_10[121],stage1_9[200]}
   );
   gpc606_5 gpc438 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[117],stage1_11[119],stage1_10[122],stage1_9[201]}
   );
   gpc606_5 gpc439 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[118],stage1_11[120],stage1_10[123],stage1_9[202]}
   );
   gpc606_5 gpc440 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[119],stage1_11[121],stage1_10[124],stage1_9[203]}
   );
   gpc606_5 gpc441 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[120],stage1_11[122],stage1_10[125],stage1_9[204]}
   );
   gpc606_5 gpc442 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[121],stage1_11[123],stage1_10[126],stage1_9[205]}
   );
   gpc606_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[122],stage1_11[124],stage1_10[127],stage1_9[206]}
   );
   gpc606_5 gpc444 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[123],stage1_11[125],stage1_10[128],stage1_9[207]}
   );
   gpc606_5 gpc445 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[124],stage1_11[126],stage1_10[129],stage1_9[208]}
   );
   gpc606_5 gpc446 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[125],stage1_11[127],stage1_10[130],stage1_9[209]}
   );
   gpc606_5 gpc447 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[126],stage1_11[128],stage1_10[131],stage1_9[210]}
   );
   gpc606_5 gpc448 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[127],stage1_11[129],stage1_10[132],stage1_9[211]}
   );
   gpc606_5 gpc449 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[128],stage1_11[130],stage1_10[133],stage1_9[212]}
   );
   gpc606_5 gpc450 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[129],stage1_11[131],stage1_10[134],stage1_9[213]}
   );
   gpc606_5 gpc451 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[130],stage1_11[132],stage1_10[135],stage1_9[214]}
   );
   gpc606_5 gpc452 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[131],stage1_11[133],stage1_10[136],stage1_9[215]}
   );
   gpc606_5 gpc453 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[132],stage1_11[134],stage1_10[137],stage1_9[216]}
   );
   gpc606_5 gpc454 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[133],stage1_11[135],stage1_10[138],stage1_9[217]}
   );
   gpc606_5 gpc455 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[134],stage1_11[136],stage1_10[139],stage1_9[218]}
   );
   gpc606_5 gpc456 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[135],stage1_11[137],stage1_10[140],stage1_9[219]}
   );
   gpc606_5 gpc457 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[136],stage1_11[138],stage1_10[141],stage1_9[220]}
   );
   gpc606_5 gpc458 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[137],stage1_11[139],stage1_10[142],stage1_9[221]}
   );
   gpc606_5 gpc459 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[138],stage1_11[140],stage1_10[143],stage1_9[222]}
   );
   gpc606_5 gpc460 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[139],stage1_11[141],stage1_10[144],stage1_9[223]}
   );
   gpc606_5 gpc461 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[140],stage1_11[142],stage1_10[145],stage1_9[224]}
   );
   gpc606_5 gpc462 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[141],stage1_11[143],stage1_10[146],stage1_9[225]}
   );
   gpc606_5 gpc463 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[142],stage1_11[144],stage1_10[147],stage1_9[226]}
   );
   gpc606_5 gpc464 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[390], stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage1_13[65],stage1_12[143],stage1_11[145],stage1_10[148],stage1_9[227]}
   );
   gpc606_5 gpc465 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400], stage0_11[401]},
      {stage1_13[66],stage1_12[144],stage1_11[146],stage1_10[149],stage1_9[228]}
   );
   gpc606_5 gpc466 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405], stage0_11[406], stage0_11[407]},
      {stage1_13[67],stage1_12[145],stage1_11[147],stage1_10[150],stage1_9[229]}
   );
   gpc606_5 gpc467 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[408], stage0_11[409], stage0_11[410], stage0_11[411], stage0_11[412], stage0_11[413]},
      {stage1_13[68],stage1_12[146],stage1_11[148],stage1_10[151],stage1_9[230]}
   );
   gpc606_5 gpc468 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419]},
      {stage1_13[69],stage1_12[147],stage1_11[149],stage1_10[152],stage1_9[231]}
   );
   gpc606_5 gpc469 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage1_13[70],stage1_12[148],stage1_11[150],stage1_10[153],stage1_9[232]}
   );
   gpc606_5 gpc470 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430], stage0_11[431]},
      {stage1_13[71],stage1_12[149],stage1_11[151],stage1_10[154],stage1_9[233]}
   );
   gpc606_5 gpc471 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435], stage0_11[436], stage0_11[437]},
      {stage1_13[72],stage1_12[150],stage1_11[152],stage1_10[155],stage1_9[234]}
   );
   gpc606_5 gpc472 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441], stage0_11[442], stage0_11[443]},
      {stage1_13[73],stage1_12[151],stage1_11[153],stage1_10[156],stage1_9[235]}
   );
   gpc606_5 gpc473 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449]},
      {stage1_13[74],stage1_12[152],stage1_11[154],stage1_10[157],stage1_9[236]}
   );
   gpc606_5 gpc474 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage1_13[75],stage1_12[153],stage1_11[155],stage1_10[158],stage1_9[237]}
   );
   gpc606_5 gpc475 (
      {stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460], stage0_11[461]},
      {stage1_13[76],stage1_12[154],stage1_11[156],stage1_10[159],stage1_9[238]}
   );
   gpc606_5 gpc476 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479]},
      {stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465], stage0_11[466], stage0_11[467]},
      {stage1_13[77],stage1_12[155],stage1_11[157],stage1_10[160],stage1_9[239]}
   );
   gpc606_5 gpc477 (
      {stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_11[468], stage0_11[469], stage0_11[470], stage0_11[471], stage0_11[472], stage0_11[473]},
      {stage1_13[78],stage1_12[156],stage1_11[158],stage1_10[161],stage1_9[240]}
   );
   gpc1_1 gpc478 (
      {stage0_2[447]},
      {stage1_2[159]}
   );
   gpc1_1 gpc479 (
      {stage0_2[448]},
      {stage1_2[160]}
   );
   gpc1_1 gpc480 (
      {stage0_2[449]},
      {stage1_2[161]}
   );
   gpc1_1 gpc481 (
      {stage0_2[450]},
      {stage1_2[162]}
   );
   gpc1_1 gpc482 (
      {stage0_2[451]},
      {stage1_2[163]}
   );
   gpc1_1 gpc483 (
      {stage0_2[452]},
      {stage1_2[164]}
   );
   gpc1_1 gpc484 (
      {stage0_2[453]},
      {stage1_2[165]}
   );
   gpc1_1 gpc485 (
      {stage0_2[454]},
      {stage1_2[166]}
   );
   gpc1_1 gpc486 (
      {stage0_2[455]},
      {stage1_2[167]}
   );
   gpc1_1 gpc487 (
      {stage0_2[456]},
      {stage1_2[168]}
   );
   gpc1_1 gpc488 (
      {stage0_2[457]},
      {stage1_2[169]}
   );
   gpc1_1 gpc489 (
      {stage0_2[458]},
      {stage1_2[170]}
   );
   gpc1_1 gpc490 (
      {stage0_2[459]},
      {stage1_2[171]}
   );
   gpc1_1 gpc491 (
      {stage0_2[460]},
      {stage1_2[172]}
   );
   gpc1_1 gpc492 (
      {stage0_2[461]},
      {stage1_2[173]}
   );
   gpc1_1 gpc493 (
      {stage0_2[462]},
      {stage1_2[174]}
   );
   gpc1_1 gpc494 (
      {stage0_2[463]},
      {stage1_2[175]}
   );
   gpc1_1 gpc495 (
      {stage0_2[464]},
      {stage1_2[176]}
   );
   gpc1_1 gpc496 (
      {stage0_2[465]},
      {stage1_2[177]}
   );
   gpc1_1 gpc497 (
      {stage0_2[466]},
      {stage1_2[178]}
   );
   gpc1_1 gpc498 (
      {stage0_2[467]},
      {stage1_2[179]}
   );
   gpc1_1 gpc499 (
      {stage0_2[468]},
      {stage1_2[180]}
   );
   gpc1_1 gpc500 (
      {stage0_2[469]},
      {stage1_2[181]}
   );
   gpc1_1 gpc501 (
      {stage0_2[470]},
      {stage1_2[182]}
   );
   gpc1_1 gpc502 (
      {stage0_2[471]},
      {stage1_2[183]}
   );
   gpc1_1 gpc503 (
      {stage0_2[472]},
      {stage1_2[184]}
   );
   gpc1_1 gpc504 (
      {stage0_2[473]},
      {stage1_2[185]}
   );
   gpc1_1 gpc505 (
      {stage0_2[474]},
      {stage1_2[186]}
   );
   gpc1_1 gpc506 (
      {stage0_2[475]},
      {stage1_2[187]}
   );
   gpc1_1 gpc507 (
      {stage0_2[476]},
      {stage1_2[188]}
   );
   gpc1_1 gpc508 (
      {stage0_2[477]},
      {stage1_2[189]}
   );
   gpc1_1 gpc509 (
      {stage0_2[478]},
      {stage1_2[190]}
   );
   gpc1_1 gpc510 (
      {stage0_2[479]},
      {stage1_2[191]}
   );
   gpc1_1 gpc511 (
      {stage0_2[480]},
      {stage1_2[192]}
   );
   gpc1_1 gpc512 (
      {stage0_2[481]},
      {stage1_2[193]}
   );
   gpc1_1 gpc513 (
      {stage0_2[482]},
      {stage1_2[194]}
   );
   gpc1_1 gpc514 (
      {stage0_2[483]},
      {stage1_2[195]}
   );
   gpc1_1 gpc515 (
      {stage0_2[484]},
      {stage1_2[196]}
   );
   gpc1_1 gpc516 (
      {stage0_2[485]},
      {stage1_2[197]}
   );
   gpc1_1 gpc517 (
      {stage0_3[450]},
      {stage1_3[160]}
   );
   gpc1_1 gpc518 (
      {stage0_3[451]},
      {stage1_3[161]}
   );
   gpc1_1 gpc519 (
      {stage0_3[452]},
      {stage1_3[162]}
   );
   gpc1_1 gpc520 (
      {stage0_3[453]},
      {stage1_3[163]}
   );
   gpc1_1 gpc521 (
      {stage0_3[454]},
      {stage1_3[164]}
   );
   gpc1_1 gpc522 (
      {stage0_3[455]},
      {stage1_3[165]}
   );
   gpc1_1 gpc523 (
      {stage0_3[456]},
      {stage1_3[166]}
   );
   gpc1_1 gpc524 (
      {stage0_3[457]},
      {stage1_3[167]}
   );
   gpc1_1 gpc525 (
      {stage0_3[458]},
      {stage1_3[168]}
   );
   gpc1_1 gpc526 (
      {stage0_3[459]},
      {stage1_3[169]}
   );
   gpc1_1 gpc527 (
      {stage0_3[460]},
      {stage1_3[170]}
   );
   gpc1_1 gpc528 (
      {stage0_3[461]},
      {stage1_3[171]}
   );
   gpc1_1 gpc529 (
      {stage0_3[462]},
      {stage1_3[172]}
   );
   gpc1_1 gpc530 (
      {stage0_3[463]},
      {stage1_3[173]}
   );
   gpc1_1 gpc531 (
      {stage0_3[464]},
      {stage1_3[174]}
   );
   gpc1_1 gpc532 (
      {stage0_3[465]},
      {stage1_3[175]}
   );
   gpc1_1 gpc533 (
      {stage0_3[466]},
      {stage1_3[176]}
   );
   gpc1_1 gpc534 (
      {stage0_3[467]},
      {stage1_3[177]}
   );
   gpc1_1 gpc535 (
      {stage0_3[468]},
      {stage1_3[178]}
   );
   gpc1_1 gpc536 (
      {stage0_3[469]},
      {stage1_3[179]}
   );
   gpc1_1 gpc537 (
      {stage0_3[470]},
      {stage1_3[180]}
   );
   gpc1_1 gpc538 (
      {stage0_3[471]},
      {stage1_3[181]}
   );
   gpc1_1 gpc539 (
      {stage0_3[472]},
      {stage1_3[182]}
   );
   gpc1_1 gpc540 (
      {stage0_3[473]},
      {stage1_3[183]}
   );
   gpc1_1 gpc541 (
      {stage0_3[474]},
      {stage1_3[184]}
   );
   gpc1_1 gpc542 (
      {stage0_3[475]},
      {stage1_3[185]}
   );
   gpc1_1 gpc543 (
      {stage0_3[476]},
      {stage1_3[186]}
   );
   gpc1_1 gpc544 (
      {stage0_3[477]},
      {stage1_3[187]}
   );
   gpc1_1 gpc545 (
      {stage0_3[478]},
      {stage1_3[188]}
   );
   gpc1_1 gpc546 (
      {stage0_3[479]},
      {stage1_3[189]}
   );
   gpc1_1 gpc547 (
      {stage0_3[480]},
      {stage1_3[190]}
   );
   gpc1_1 gpc548 (
      {stage0_3[481]},
      {stage1_3[191]}
   );
   gpc1_1 gpc549 (
      {stage0_3[482]},
      {stage1_3[192]}
   );
   gpc1_1 gpc550 (
      {stage0_3[483]},
      {stage1_3[193]}
   );
   gpc1_1 gpc551 (
      {stage0_3[484]},
      {stage1_3[194]}
   );
   gpc1_1 gpc552 (
      {stage0_3[485]},
      {stage1_3[195]}
   );
   gpc1_1 gpc553 (
      {stage0_4[481]},
      {stage1_4[236]}
   );
   gpc1_1 gpc554 (
      {stage0_4[482]},
      {stage1_4[237]}
   );
   gpc1_1 gpc555 (
      {stage0_4[483]},
      {stage1_4[238]}
   );
   gpc1_1 gpc556 (
      {stage0_4[484]},
      {stage1_4[239]}
   );
   gpc1_1 gpc557 (
      {stage0_4[485]},
      {stage1_4[240]}
   );
   gpc1_1 gpc558 (
      {stage0_6[480]},
      {stage1_6[164]}
   );
   gpc1_1 gpc559 (
      {stage0_6[481]},
      {stage1_6[165]}
   );
   gpc1_1 gpc560 (
      {stage0_6[482]},
      {stage1_6[166]}
   );
   gpc1_1 gpc561 (
      {stage0_6[483]},
      {stage1_6[167]}
   );
   gpc1_1 gpc562 (
      {stage0_6[484]},
      {stage1_6[168]}
   );
   gpc1_1 gpc563 (
      {stage0_6[485]},
      {stage1_6[169]}
   );
   gpc1_1 gpc564 (
      {stage0_10[468]},
      {stage1_10[162]}
   );
   gpc1_1 gpc565 (
      {stage0_10[469]},
      {stage1_10[163]}
   );
   gpc1_1 gpc566 (
      {stage0_10[470]},
      {stage1_10[164]}
   );
   gpc1_1 gpc567 (
      {stage0_10[471]},
      {stage1_10[165]}
   );
   gpc1_1 gpc568 (
      {stage0_10[472]},
      {stage1_10[166]}
   );
   gpc1_1 gpc569 (
      {stage0_10[473]},
      {stage1_10[167]}
   );
   gpc1_1 gpc570 (
      {stage0_10[474]},
      {stage1_10[168]}
   );
   gpc1_1 gpc571 (
      {stage0_10[475]},
      {stage1_10[169]}
   );
   gpc1_1 gpc572 (
      {stage0_10[476]},
      {stage1_10[170]}
   );
   gpc1_1 gpc573 (
      {stage0_10[477]},
      {stage1_10[171]}
   );
   gpc1_1 gpc574 (
      {stage0_10[478]},
      {stage1_10[172]}
   );
   gpc1_1 gpc575 (
      {stage0_10[479]},
      {stage1_10[173]}
   );
   gpc1_1 gpc576 (
      {stage0_10[480]},
      {stage1_10[174]}
   );
   gpc1_1 gpc577 (
      {stage0_10[481]},
      {stage1_10[175]}
   );
   gpc1_1 gpc578 (
      {stage0_10[482]},
      {stage1_10[176]}
   );
   gpc1_1 gpc579 (
      {stage0_10[483]},
      {stage1_10[177]}
   );
   gpc1_1 gpc580 (
      {stage0_10[484]},
      {stage1_10[178]}
   );
   gpc1_1 gpc581 (
      {stage0_10[485]},
      {stage1_10[179]}
   );
   gpc1_1 gpc582 (
      {stage0_11[474]},
      {stage1_11[159]}
   );
   gpc1_1 gpc583 (
      {stage0_11[475]},
      {stage1_11[160]}
   );
   gpc1_1 gpc584 (
      {stage0_11[476]},
      {stage1_11[161]}
   );
   gpc1_1 gpc585 (
      {stage0_11[477]},
      {stage1_11[162]}
   );
   gpc1_1 gpc586 (
      {stage0_11[478]},
      {stage1_11[163]}
   );
   gpc1_1 gpc587 (
      {stage0_11[479]},
      {stage1_11[164]}
   );
   gpc1_1 gpc588 (
      {stage0_11[480]},
      {stage1_11[165]}
   );
   gpc1_1 gpc589 (
      {stage0_11[481]},
      {stage1_11[166]}
   );
   gpc1_1 gpc590 (
      {stage0_11[482]},
      {stage1_11[167]}
   );
   gpc1_1 gpc591 (
      {stage0_11[483]},
      {stage1_11[168]}
   );
   gpc1_1 gpc592 (
      {stage0_11[484]},
      {stage1_11[169]}
   );
   gpc1_1 gpc593 (
      {stage0_11[485]},
      {stage1_11[170]}
   );
   gpc1163_5 gpc594 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc595 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc596 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc597 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc598 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc599 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc600 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc601 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc602 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc603 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc604 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc605 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc606 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc607 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc608 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc609 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc1163_5 gpc610 (
      {stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_2[16]},
      {stage1_3[16]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc1163_5 gpc611 (
      {stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_2[17]},
      {stage1_3[17]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc1163_5 gpc612 (
      {stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_2[18]},
      {stage1_3[18]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc1163_5 gpc613 (
      {stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_2[19]},
      {stage1_3[19]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc614 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc615 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc616 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc617 (
      {stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc618 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc606_5 gpc619 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc606_5 gpc620 (
      {stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc621 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc622 (
      {stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage1_3[20]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc623 (
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_3[21]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc624 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[22]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30]}
   );
   gpc615_5 gpc625 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[23]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc615_5 gpc626 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[24]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc615_5 gpc627 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[25]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc615_5 gpc628 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[26]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc615_5 gpc629 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[27]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc615_5 gpc630 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[28]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc631 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[29]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc632 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[30]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc633 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[31]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc634 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[32]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc635 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[33]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc636 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[34]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc637 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[35]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc638 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[36]},
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage2_6[21],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc639 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[37]},
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136], stage1_4[137]},
      {stage2_6[22],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc640 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[38]},
      {stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143]},
      {stage2_6[23],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc641 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[39]},
      {stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149]},
      {stage2_6[24],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc642 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[40]},
      {stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage2_6[25],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc643 (
      {stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_3[41]},
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage2_6[26],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc644 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182]},
      {stage1_3[42]},
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167]},
      {stage2_6[27],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc645 (
      {stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187]},
      {stage1_3[43]},
      {stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173]},
      {stage2_6[28],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc646 (
      {stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_3[44]},
      {stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179]},
      {stage2_6[29],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc647 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197]},
      {stage1_3[45]},
      {stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage2_6[30],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc648 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[186]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[31],stage2_5[31],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc649 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[187]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[32],stage2_5[32],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc650 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[188]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[33],stage2_5[33],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc651 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[189]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[34],stage2_5[34],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc652 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[190]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[35],stage2_5[35],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc653 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[191]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[36],stage2_5[36],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc654 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[192]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[37],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc655 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[193]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[38],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc656 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[194]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[39],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc657 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[195]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[40],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc658 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[196]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[41],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc659 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[197]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[42],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc660 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[198]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[43],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc661 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[199]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[44],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc662 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[200]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[45],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc663 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[201]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[46],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc664 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[202]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[47],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc665 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[203]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[48],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc666 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[204]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[49],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc667 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[205]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[50],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc668 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[206]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[51],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc669 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[207]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[52],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc670 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[208]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[53],stage2_5[53],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc671 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[209]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[54],stage2_5[54],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc672 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[210]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[55],stage2_5[55],stage2_4[78],stage2_3[78]}
   );
   gpc615_5 gpc673 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[211]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[56],stage2_5[56],stage2_4[79],stage2_3[79]}
   );
   gpc615_5 gpc674 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[212]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[57],stage2_5[57],stage2_4[80],stage2_3[80]}
   );
   gpc615_5 gpc675 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[213]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[58],stage2_5[58],stage2_4[81],stage2_3[81]}
   );
   gpc615_5 gpc676 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[214]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[59],stage2_5[59],stage2_4[82],stage2_3[82]}
   );
   gpc615_5 gpc677 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[215]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[60],stage2_5[60],stage2_4[83],stage2_3[83]}
   );
   gpc606_5 gpc678 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[30],stage2_6[61],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc679 (
      {stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[31],stage2_6[62],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc680 (
      {stage1_4[228], stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[32],stage2_6[63],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc681 (
      {stage1_4[234], stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[33],stage2_6[64],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc682 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[34],stage2_6[65],stage2_5[65]}
   );
   gpc606_5 gpc683 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[5],stage2_7[35],stage2_6[66],stage2_5[66]}
   );
   gpc606_5 gpc684 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[6],stage2_7[36],stage2_6[67],stage2_5[67]}
   );
   gpc606_5 gpc685 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[7],stage2_7[37],stage2_6[68],stage2_5[68]}
   );
   gpc606_5 gpc686 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[8],stage2_7[38],stage2_6[69],stage2_5[69]}
   );
   gpc606_5 gpc687 (
      {stage1_5[210], stage1_5[211], stage1_5[212], stage1_5[213], stage1_5[214], stage1_5[215]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[9],stage2_7[39],stage2_6[70],stage2_5[70]}
   );
   gpc606_5 gpc688 (
      {stage1_5[216], stage1_5[217], stage1_5[218], stage1_5[219], stage1_5[220], stage1_5[221]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[10],stage2_7[40],stage2_6[71],stage2_5[71]}
   );
   gpc606_5 gpc689 (
      {stage1_5[222], stage1_5[223], stage1_5[224], stage1_5[225], stage1_5[226], stage1_5[227]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[11],stage2_7[41],stage2_6[72],stage2_5[72]}
   );
   gpc606_5 gpc690 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[12],stage2_7[42],stage2_6[73]}
   );
   gpc606_5 gpc691 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[13],stage2_7[43],stage2_6[74]}
   );
   gpc606_5 gpc692 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[14],stage2_7[44],stage2_6[75]}
   );
   gpc606_5 gpc693 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[15],stage2_7[45],stage2_6[76]}
   );
   gpc606_5 gpc694 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[16],stage2_7[46],stage2_6[77]}
   );
   gpc606_5 gpc695 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[17],stage2_7[47],stage2_6[78]}
   );
   gpc606_5 gpc696 (
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[18],stage2_7[48],stage2_6[79]}
   );
   gpc606_5 gpc697 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[19],stage2_7[49],stage2_6[80]}
   );
   gpc606_5 gpc698 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[20],stage2_7[50],stage2_6[81]}
   );
   gpc606_5 gpc699 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[21],stage2_7[51],stage2_6[82]}
   );
   gpc606_5 gpc700 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[22],stage2_7[52],stage2_6[83]}
   );
   gpc606_5 gpc701 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[23],stage2_7[53],stage2_6[84]}
   );
   gpc606_5 gpc702 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[24],stage2_7[54],stage2_6[85]}
   );
   gpc606_5 gpc703 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[25],stage2_7[55],stage2_6[86]}
   );
   gpc606_5 gpc704 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[26],stage2_7[56],stage2_6[87]}
   );
   gpc606_5 gpc705 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[23],stage2_8[27],stage2_7[57],stage2_6[88]}
   );
   gpc606_5 gpc706 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[24],stage2_8[28],stage2_7[58],stage2_6[89]}
   );
   gpc606_5 gpc707 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[25],stage2_8[29],stage2_7[59],stage2_6[90]}
   );
   gpc606_5 gpc708 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[26],stage2_8[30],stage2_7[60],stage2_6[91]}
   );
   gpc606_5 gpc709 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[27],stage2_8[31],stage2_7[61],stage2_6[92]}
   );
   gpc606_5 gpc710 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[28],stage2_8[32],stage2_7[62],stage2_6[93]}
   );
   gpc615_5 gpc711 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154]},
      {stage1_7[48]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[29],stage2_8[33],stage2_7[63],stage2_6[94]}
   );
   gpc615_5 gpc712 (
      {stage1_6[155], stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159]},
      {stage1_7[49]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[30],stage2_8[34],stage2_7[64],stage2_6[95]}
   );
   gpc615_5 gpc713 (
      {stage1_6[160], stage1_6[161], stage1_6[162], stage1_6[163], stage1_6[164]},
      {stage1_7[50]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[31],stage2_8[35],stage2_7[65],stage2_6[96]}
   );
   gpc615_5 gpc714 (
      {stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168], stage1_6[169]},
      {stage1_7[51]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[32],stage2_8[36],stage2_7[66],stage2_6[97]}
   );
   gpc615_5 gpc715 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[150]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[25],stage2_9[33],stage2_8[37],stage2_7[67]}
   );
   gpc615_5 gpc716 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[151]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[26],stage2_9[34],stage2_8[38],stage2_7[68]}
   );
   gpc615_5 gpc717 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[152]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[27],stage2_9[35],stage2_8[39],stage2_7[69]}
   );
   gpc615_5 gpc718 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[153]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[28],stage2_9[36],stage2_8[40],stage2_7[70]}
   );
   gpc615_5 gpc719 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[154]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[29],stage2_9[37],stage2_8[41],stage2_7[71]}
   );
   gpc615_5 gpc720 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[155]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[30],stage2_9[38],stage2_8[42],stage2_7[72]}
   );
   gpc615_5 gpc721 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[156]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[31],stage2_9[39],stage2_8[43],stage2_7[73]}
   );
   gpc615_5 gpc722 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[157]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[32],stage2_9[40],stage2_8[44],stage2_7[74]}
   );
   gpc615_5 gpc723 (
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_8[158]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[33],stage2_9[41],stage2_8[45],stage2_7[75]}
   );
   gpc615_5 gpc724 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage1_8[159]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[34],stage2_9[42],stage2_8[46],stage2_7[76]}
   );
   gpc615_5 gpc725 (
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106]},
      {stage1_8[160]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[35],stage2_9[43],stage2_8[47],stage2_7[77]}
   );
   gpc615_5 gpc726 (
      {stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111]},
      {stage1_8[161]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[36],stage2_9[44],stage2_8[48],stage2_7[78]}
   );
   gpc615_5 gpc727 (
      {stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115], stage1_7[116]},
      {stage1_8[162]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[37],stage2_9[45],stage2_8[49],stage2_7[79]}
   );
   gpc615_5 gpc728 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[163]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[38],stage2_9[46],stage2_8[50],stage2_7[80]}
   );
   gpc615_5 gpc729 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[164]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[39],stage2_9[47],stage2_8[51],stage2_7[81]}
   );
   gpc615_5 gpc730 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[165]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[40],stage2_9[48],stage2_8[52],stage2_7[82]}
   );
   gpc615_5 gpc731 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[166]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[41],stage2_9[49],stage2_8[53],stage2_7[83]}
   );
   gpc615_5 gpc732 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[167]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[42],stage2_9[50],stage2_8[54],stage2_7[84]}
   );
   gpc615_5 gpc733 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[168]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[43],stage2_9[51],stage2_8[55],stage2_7[85]}
   );
   gpc615_5 gpc734 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[169]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[44],stage2_9[52],stage2_8[56],stage2_7[86]}
   );
   gpc615_5 gpc735 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[170]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[45],stage2_9[53],stage2_8[57],stage2_7[87]}
   );
   gpc615_5 gpc736 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[171]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[46],stage2_9[54],stage2_8[58],stage2_7[88]}
   );
   gpc606_5 gpc737 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[22],stage2_10[47],stage2_9[55],stage2_8[59]}
   );
   gpc606_5 gpc738 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[23],stage2_10[48],stage2_9[56],stage2_8[60]}
   );
   gpc606_5 gpc739 (
      {stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187], stage1_8[188], stage1_8[189]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[24],stage2_10[49],stage2_9[57],stage2_8[61]}
   );
   gpc606_5 gpc740 (
      {stage1_8[190], stage1_8[191], stage1_8[192], stage1_8[193], stage1_8[194], stage1_8[195]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[25],stage2_10[50],stage2_9[58],stage2_8[62]}
   );
   gpc606_5 gpc741 (
      {stage1_8[196], stage1_8[197], stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[26],stage2_10[51],stage2_9[59],stage2_8[63]}
   );
   gpc606_5 gpc742 (
      {stage1_8[202], stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[27],stage2_10[52],stage2_9[60],stage2_8[64]}
   );
   gpc606_5 gpc743 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212], stage1_8[213]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[28],stage2_10[53],stage2_9[61],stage2_8[65]}
   );
   gpc615_5 gpc744 (
      {stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217], stage1_8[218]},
      {stage1_9[132]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[29],stage2_10[54],stage2_9[62],stage2_8[66]}
   );
   gpc615_5 gpc745 (
      {stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222], stage1_8[223]},
      {stage1_9[133]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[30],stage2_10[55],stage2_9[63],stage2_8[67]}
   );
   gpc615_5 gpc746 (
      {stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_9[134]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[31],stage2_10[56],stage2_9[64],stage2_8[68]}
   );
   gpc615_5 gpc747 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233]},
      {stage1_9[135]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[32],stage2_10[57],stage2_9[65],stage2_8[69]}
   );
   gpc615_5 gpc748 (
      {stage1_8[234], stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238]},
      {stage1_9[136]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[33],stage2_10[58],stage2_9[66],stage2_8[70]}
   );
   gpc606_5 gpc749 (
      {stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[12],stage2_11[34],stage2_10[59],stage2_9[67]}
   );
   gpc606_5 gpc750 (
      {stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[13],stage2_11[35],stage2_10[60],stage2_9[68]}
   );
   gpc606_5 gpc751 (
      {stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[14],stage2_11[36],stage2_10[61],stage2_9[69]}
   );
   gpc606_5 gpc752 (
      {stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[15],stage2_11[37],stage2_10[62],stage2_9[70]}
   );
   gpc606_5 gpc753 (
      {stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[16],stage2_11[38],stage2_10[63],stage2_9[71]}
   );
   gpc606_5 gpc754 (
      {stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[17],stage2_11[39],stage2_10[64],stage2_9[72]}
   );
   gpc606_5 gpc755 (
      {stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[18],stage2_11[40],stage2_10[65],stage2_9[73]}
   );
   gpc615_5 gpc756 (
      {stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_10[72]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[19],stage2_11[41],stage2_10[66],stage2_9[74]}
   );
   gpc615_5 gpc757 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188]},
      {stage1_10[73]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[20],stage2_11[42],stage2_10[67],stage2_9[75]}
   );
   gpc615_5 gpc758 (
      {stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193]},
      {stage1_10[74]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[21],stage2_11[43],stage2_10[68],stage2_9[76]}
   );
   gpc615_5 gpc759 (
      {stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_10[75]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[22],stage2_11[44],stage2_10[69],stage2_9[77]}
   );
   gpc615_5 gpc760 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_10[76]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[23],stage2_11[45],stage2_10[70],stage2_9[78]}
   );
   gpc615_5 gpc761 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208]},
      {stage1_10[77]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[24],stage2_11[46],stage2_10[71],stage2_9[79]}
   );
   gpc615_5 gpc762 (
      {stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_10[78]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[25],stage2_11[47],stage2_10[72],stage2_9[80]}
   );
   gpc615_5 gpc763 (
      {stage1_9[214], stage1_9[215], stage1_9[216], stage1_9[217], stage1_9[218]},
      {stage1_10[79]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[26],stage2_11[48],stage2_10[73],stage2_9[81]}
   );
   gpc615_5 gpc764 (
      {stage1_9[219], stage1_9[220], stage1_9[221], stage1_9[222], stage1_9[223]},
      {stage1_10[80]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[27],stage2_11[49],stage2_10[74],stage2_9[82]}
   );
   gpc615_5 gpc765 (
      {stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227], stage1_9[228]},
      {stage1_10[81]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[28],stage2_11[50],stage2_10[75],stage2_9[83]}
   );
   gpc615_5 gpc766 (
      {stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage1_10[82]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[29],stage2_11[51],stage2_10[76],stage2_9[84]}
   );
   gpc606_5 gpc767 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[30],stage2_11[52],stage2_10[77]}
   );
   gpc606_5 gpc768 (
      {stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[19],stage2_12[31],stage2_11[53],stage2_10[78]}
   );
   gpc606_5 gpc769 (
      {stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[20],stage2_12[32],stage2_11[54],stage2_10[79]}
   );
   gpc606_5 gpc770 (
      {stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[21],stage2_12[33],stage2_11[55],stage2_10[80]}
   );
   gpc606_5 gpc771 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[22],stage2_12[34],stage2_11[56],stage2_10[81]}
   );
   gpc606_5 gpc772 (
      {stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[23],stage2_12[35],stage2_11[57],stage2_10[82]}
   );
   gpc606_5 gpc773 (
      {stage1_10[119], stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[24],stage2_12[36],stage2_11[58],stage2_10[83]}
   );
   gpc606_5 gpc774 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[25],stage2_12[37],stage2_11[59],stage2_10[84]}
   );
   gpc606_5 gpc775 (
      {stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[26],stage2_12[38],stage2_11[60],stage2_10[85]}
   );
   gpc606_5 gpc776 (
      {stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[27],stage2_12[39],stage2_11[61],stage2_10[86]}
   );
   gpc606_5 gpc777 (
      {stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[28],stage2_12[40],stage2_11[62],stage2_10[87]}
   );
   gpc606_5 gpc778 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[29],stage2_12[41],stage2_11[63],stage2_10[88]}
   );
   gpc606_5 gpc779 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[30],stage2_12[42],stage2_11[64],stage2_10[89]}
   );
   gpc606_5 gpc780 (
      {stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[31],stage2_12[43],stage2_11[65],stage2_10[90]}
   );
   gpc606_5 gpc781 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[32],stage2_12[44],stage2_11[66],stage2_10[91]}
   );
   gpc615_5 gpc782 (
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112]},
      {stage1_12[90]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[15],stage2_13[33],stage2_12[45],stage2_11[67]}
   );
   gpc615_5 gpc783 (
      {stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[91]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[16],stage2_13[34],stage2_12[46],stage2_11[68]}
   );
   gpc615_5 gpc784 (
      {stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122]},
      {stage1_12[92]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[17],stage2_13[35],stage2_12[47],stage2_11[69]}
   );
   gpc615_5 gpc785 (
      {stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127]},
      {stage1_12[93]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[18],stage2_13[36],stage2_12[48],stage2_11[70]}
   );
   gpc615_5 gpc786 (
      {stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[94]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[19],stage2_13[37],stage2_12[49],stage2_11[71]}
   );
   gpc615_5 gpc787 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[95]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[20],stage2_13[38],stage2_12[50],stage2_11[72]}
   );
   gpc615_5 gpc788 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[96]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[21],stage2_13[39],stage2_12[51],stage2_11[73]}
   );
   gpc615_5 gpc789 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[97]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[22],stage2_13[40],stage2_12[52],stage2_11[74]}
   );
   gpc615_5 gpc790 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[98]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[23],stage2_13[41],stage2_12[53],stage2_11[75]}
   );
   gpc615_5 gpc791 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[99]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[24],stage2_13[42],stage2_12[54],stage2_11[76]}
   );
   gpc615_5 gpc792 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[100]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[25],stage2_13[43],stage2_12[55],stage2_11[77]}
   );
   gpc615_5 gpc793 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[101]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[26],stage2_13[44],stage2_12[56],stage2_11[78]}
   );
   gpc1_1 gpc794 (
      {stage1_0[78]},
      {stage2_0[23]}
   );
   gpc1_1 gpc795 (
      {stage1_0[79]},
      {stage2_0[24]}
   );
   gpc1_1 gpc796 (
      {stage1_0[80]},
      {stage2_0[25]}
   );
   gpc1_1 gpc797 (
      {stage1_0[81]},
      {stage2_0[26]}
   );
   gpc1_1 gpc798 (
      {stage1_0[82]},
      {stage2_0[27]}
   );
   gpc1_1 gpc799 (
      {stage1_0[83]},
      {stage2_0[28]}
   );
   gpc1_1 gpc800 (
      {stage1_0[84]},
      {stage2_0[29]}
   );
   gpc1_1 gpc801 (
      {stage1_0[85]},
      {stage2_0[30]}
   );
   gpc1_1 gpc802 (
      {stage1_1[120]},
      {stage2_1[23]}
   );
   gpc1_1 gpc803 (
      {stage1_1[121]},
      {stage2_1[24]}
   );
   gpc1_1 gpc804 (
      {stage1_1[122]},
      {stage2_1[25]}
   );
   gpc1_1 gpc805 (
      {stage1_1[123]},
      {stage2_1[26]}
   );
   gpc1_1 gpc806 (
      {stage1_1[124]},
      {stage2_1[27]}
   );
   gpc1_1 gpc807 (
      {stage1_1[125]},
      {stage2_1[28]}
   );
   gpc1_1 gpc808 (
      {stage1_1[126]},
      {stage2_1[29]}
   );
   gpc1_1 gpc809 (
      {stage1_1[127]},
      {stage2_1[30]}
   );
   gpc1_1 gpc810 (
      {stage1_1[128]},
      {stage2_1[31]}
   );
   gpc1_1 gpc811 (
      {stage1_1[129]},
      {stage2_1[32]}
   );
   gpc1_1 gpc812 (
      {stage1_1[130]},
      {stage2_1[33]}
   );
   gpc1_1 gpc813 (
      {stage1_1[131]},
      {stage2_1[34]}
   );
   gpc1_1 gpc814 (
      {stage1_1[132]},
      {stage2_1[35]}
   );
   gpc1_1 gpc815 (
      {stage1_1[133]},
      {stage2_1[36]}
   );
   gpc1_1 gpc816 (
      {stage1_1[134]},
      {stage2_1[37]}
   );
   gpc1_1 gpc817 (
      {stage1_1[135]},
      {stage2_1[38]}
   );
   gpc1_1 gpc818 (
      {stage1_1[136]},
      {stage2_1[39]}
   );
   gpc1_1 gpc819 (
      {stage1_1[137]},
      {stage2_1[40]}
   );
   gpc1_1 gpc820 (
      {stage1_1[138]},
      {stage2_1[41]}
   );
   gpc1_1 gpc821 (
      {stage1_1[139]},
      {stage2_1[42]}
   );
   gpc1_1 gpc822 (
      {stage1_1[140]},
      {stage2_1[43]}
   );
   gpc1_1 gpc823 (
      {stage1_1[141]},
      {stage2_1[44]}
   );
   gpc1_1 gpc824 (
      {stage1_1[142]},
      {stage2_1[45]}
   );
   gpc1_1 gpc825 (
      {stage1_1[143]},
      {stage2_1[46]}
   );
   gpc1_1 gpc826 (
      {stage1_1[144]},
      {stage2_1[47]}
   );
   gpc1_1 gpc827 (
      {stage1_1[145]},
      {stage2_1[48]}
   );
   gpc1_1 gpc828 (
      {stage1_1[146]},
      {stage2_1[49]}
   );
   gpc1_1 gpc829 (
      {stage1_1[147]},
      {stage2_1[50]}
   );
   gpc1_1 gpc830 (
      {stage1_1[148]},
      {stage2_1[51]}
   );
   gpc1_1 gpc831 (
      {stage1_1[149]},
      {stage2_1[52]}
   );
   gpc1_1 gpc832 (
      {stage1_1[150]},
      {stage2_1[53]}
   );
   gpc1_1 gpc833 (
      {stage1_1[151]},
      {stage2_1[54]}
   );
   gpc1_1 gpc834 (
      {stage1_1[152]},
      {stage2_1[55]}
   );
   gpc1_1 gpc835 (
      {stage1_1[153]},
      {stage2_1[56]}
   );
   gpc1_1 gpc836 (
      {stage1_1[154]},
      {stage2_1[57]}
   );
   gpc1_1 gpc837 (
      {stage1_4[240]},
      {stage2_4[88]}
   );
   gpc1_1 gpc838 (
      {stage1_5[228]},
      {stage2_5[73]}
   );
   gpc1_1 gpc839 (
      {stage1_5[229]},
      {stage2_5[74]}
   );
   gpc1_1 gpc840 (
      {stage1_9[234]},
      {stage2_9[85]}
   );
   gpc1_1 gpc841 (
      {stage1_9[235]},
      {stage2_9[86]}
   );
   gpc1_1 gpc842 (
      {stage1_9[236]},
      {stage2_9[87]}
   );
   gpc1_1 gpc843 (
      {stage1_9[237]},
      {stage2_9[88]}
   );
   gpc1_1 gpc844 (
      {stage1_9[238]},
      {stage2_9[89]}
   );
   gpc1_1 gpc845 (
      {stage1_9[239]},
      {stage2_9[90]}
   );
   gpc1_1 gpc846 (
      {stage1_9[240]},
      {stage2_9[91]}
   );
   gpc1_1 gpc847 (
      {stage1_10[173]},
      {stage2_10[92]}
   );
   gpc1_1 gpc848 (
      {stage1_10[174]},
      {stage2_10[93]}
   );
   gpc1_1 gpc849 (
      {stage1_10[175]},
      {stage2_10[94]}
   );
   gpc1_1 gpc850 (
      {stage1_10[176]},
      {stage2_10[95]}
   );
   gpc1_1 gpc851 (
      {stage1_10[177]},
      {stage2_10[96]}
   );
   gpc1_1 gpc852 (
      {stage1_10[178]},
      {stage2_10[97]}
   );
   gpc1_1 gpc853 (
      {stage1_10[179]},
      {stage2_10[98]}
   );
   gpc1_1 gpc854 (
      {stage1_11[168]},
      {stage2_11[79]}
   );
   gpc1_1 gpc855 (
      {stage1_11[169]},
      {stage2_11[80]}
   );
   gpc1_1 gpc856 (
      {stage1_11[170]},
      {stage2_11[81]}
   );
   gpc1_1 gpc857 (
      {stage1_12[102]},
      {stage2_12[57]}
   );
   gpc1_1 gpc858 (
      {stage1_12[103]},
      {stage2_12[58]}
   );
   gpc1_1 gpc859 (
      {stage1_12[104]},
      {stage2_12[59]}
   );
   gpc1_1 gpc860 (
      {stage1_12[105]},
      {stage2_12[60]}
   );
   gpc1_1 gpc861 (
      {stage1_12[106]},
      {stage2_12[61]}
   );
   gpc1_1 gpc862 (
      {stage1_12[107]},
      {stage2_12[62]}
   );
   gpc1_1 gpc863 (
      {stage1_12[108]},
      {stage2_12[63]}
   );
   gpc1_1 gpc864 (
      {stage1_12[109]},
      {stage2_12[64]}
   );
   gpc1_1 gpc865 (
      {stage1_12[110]},
      {stage2_12[65]}
   );
   gpc1_1 gpc866 (
      {stage1_12[111]},
      {stage2_12[66]}
   );
   gpc1_1 gpc867 (
      {stage1_12[112]},
      {stage2_12[67]}
   );
   gpc1_1 gpc868 (
      {stage1_12[113]},
      {stage2_12[68]}
   );
   gpc1_1 gpc869 (
      {stage1_12[114]},
      {stage2_12[69]}
   );
   gpc1_1 gpc870 (
      {stage1_12[115]},
      {stage2_12[70]}
   );
   gpc1_1 gpc871 (
      {stage1_12[116]},
      {stage2_12[71]}
   );
   gpc1_1 gpc872 (
      {stage1_12[117]},
      {stage2_12[72]}
   );
   gpc1_1 gpc873 (
      {stage1_12[118]},
      {stage2_12[73]}
   );
   gpc1_1 gpc874 (
      {stage1_12[119]},
      {stage2_12[74]}
   );
   gpc1_1 gpc875 (
      {stage1_12[120]},
      {stage2_12[75]}
   );
   gpc1_1 gpc876 (
      {stage1_12[121]},
      {stage2_12[76]}
   );
   gpc1_1 gpc877 (
      {stage1_12[122]},
      {stage2_12[77]}
   );
   gpc1_1 gpc878 (
      {stage1_12[123]},
      {stage2_12[78]}
   );
   gpc1_1 gpc879 (
      {stage1_12[124]},
      {stage2_12[79]}
   );
   gpc1_1 gpc880 (
      {stage1_12[125]},
      {stage2_12[80]}
   );
   gpc1_1 gpc881 (
      {stage1_12[126]},
      {stage2_12[81]}
   );
   gpc1_1 gpc882 (
      {stage1_12[127]},
      {stage2_12[82]}
   );
   gpc1_1 gpc883 (
      {stage1_12[128]},
      {stage2_12[83]}
   );
   gpc1_1 gpc884 (
      {stage1_12[129]},
      {stage2_12[84]}
   );
   gpc1_1 gpc885 (
      {stage1_12[130]},
      {stage2_12[85]}
   );
   gpc1_1 gpc886 (
      {stage1_12[131]},
      {stage2_12[86]}
   );
   gpc1_1 gpc887 (
      {stage1_12[132]},
      {stage2_12[87]}
   );
   gpc1_1 gpc888 (
      {stage1_12[133]},
      {stage2_12[88]}
   );
   gpc1_1 gpc889 (
      {stage1_12[134]},
      {stage2_12[89]}
   );
   gpc1_1 gpc890 (
      {stage1_12[135]},
      {stage2_12[90]}
   );
   gpc1_1 gpc891 (
      {stage1_12[136]},
      {stage2_12[91]}
   );
   gpc1_1 gpc892 (
      {stage1_12[137]},
      {stage2_12[92]}
   );
   gpc1_1 gpc893 (
      {stage1_12[138]},
      {stage2_12[93]}
   );
   gpc1_1 gpc894 (
      {stage1_12[139]},
      {stage2_12[94]}
   );
   gpc1_1 gpc895 (
      {stage1_12[140]},
      {stage2_12[95]}
   );
   gpc1_1 gpc896 (
      {stage1_12[141]},
      {stage2_12[96]}
   );
   gpc1_1 gpc897 (
      {stage1_12[142]},
      {stage2_12[97]}
   );
   gpc1_1 gpc898 (
      {stage1_12[143]},
      {stage2_12[98]}
   );
   gpc1_1 gpc899 (
      {stage1_12[144]},
      {stage2_12[99]}
   );
   gpc1_1 gpc900 (
      {stage1_12[145]},
      {stage2_12[100]}
   );
   gpc1_1 gpc901 (
      {stage1_12[146]},
      {stage2_12[101]}
   );
   gpc1_1 gpc902 (
      {stage1_12[147]},
      {stage2_12[102]}
   );
   gpc1_1 gpc903 (
      {stage1_12[148]},
      {stage2_12[103]}
   );
   gpc1_1 gpc904 (
      {stage1_12[149]},
      {stage2_12[104]}
   );
   gpc1_1 gpc905 (
      {stage1_12[150]},
      {stage2_12[105]}
   );
   gpc1_1 gpc906 (
      {stage1_12[151]},
      {stage2_12[106]}
   );
   gpc1_1 gpc907 (
      {stage1_12[152]},
      {stage2_12[107]}
   );
   gpc1_1 gpc908 (
      {stage1_12[153]},
      {stage2_12[108]}
   );
   gpc1_1 gpc909 (
      {stage1_12[154]},
      {stage2_12[109]}
   );
   gpc1_1 gpc910 (
      {stage1_12[155]},
      {stage2_12[110]}
   );
   gpc1_1 gpc911 (
      {stage1_12[156]},
      {stage2_12[111]}
   );
   gpc1_1 gpc912 (
      {stage1_13[72]},
      {stage2_13[45]}
   );
   gpc1_1 gpc913 (
      {stage1_13[73]},
      {stage2_13[46]}
   );
   gpc1_1 gpc914 (
      {stage1_13[74]},
      {stage2_13[47]}
   );
   gpc1_1 gpc915 (
      {stage1_13[75]},
      {stage2_13[48]}
   );
   gpc1_1 gpc916 (
      {stage1_13[76]},
      {stage2_13[49]}
   );
   gpc1_1 gpc917 (
      {stage1_13[77]},
      {stage2_13[50]}
   );
   gpc1_1 gpc918 (
      {stage1_13[78]},
      {stage2_13[51]}
   );
   gpc1163_5 gpc919 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc920 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc921 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc922 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc923 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc924 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc925 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc926 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc927 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc928 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc615_5 gpc929 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[37]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc930 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[38]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc931 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[39]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc932 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc933 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc934 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc935 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc936 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc937 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc938 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc939 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc940 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc941 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73]},
      {stage2_4[47]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc942 (
      {stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78]},
      {stage2_4[48]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc943 (
      {stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83]},
      {stage2_4[49]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc606_5 gpc944 (
      {stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25]}
   );
   gpc606_5 gpc945 (
      {stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26]}
   );
   gpc606_5 gpc946 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27]}
   );
   gpc606_5 gpc947 (
      {stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28]}
   );
   gpc606_5 gpc948 (
      {stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc949 (
      {stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc950 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[6],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc951 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[7],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc615_5 gpc952 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_6[36]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[8],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc615_5 gpc953 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage2_6[37]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[9],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc615_5 gpc954 (
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74]},
      {stage2_6[38]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[10],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc615_5 gpc955 (
      {stage2_6[39], stage2_6[40], stage2_6[41], stage2_6[42], stage2_6[43]},
      {stage2_7[30]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[11],stage3_7[19],stage3_6[26]}
   );
   gpc615_5 gpc956 (
      {stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47], stage2_6[48]},
      {stage2_7[31]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[12],stage3_7[20],stage3_6[27]}
   );
   gpc615_5 gpc957 (
      {stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage2_7[32]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[7],stage3_8[13],stage3_7[21],stage3_6[28]}
   );
   gpc615_5 gpc958 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[33]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[8],stage3_8[14],stage3_7[22],stage3_6[29]}
   );
   gpc615_5 gpc959 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[34]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[9],stage3_8[15],stage3_7[23],stage3_6[30]}
   );
   gpc615_5 gpc960 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[35]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[10],stage3_8[16],stage3_7[24],stage3_6[31]}
   );
   gpc615_5 gpc961 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[36]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[11],stage3_8[17],stage3_7[25],stage3_6[32]}
   );
   gpc615_5 gpc962 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[37]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[12],stage3_8[18],stage3_7[26],stage3_6[33]}
   );
   gpc615_5 gpc963 (
      {stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage2_7[38]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[13],stage3_8[19],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc964 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[39]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[14],stage3_8[20],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc965 (
      {stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[10],stage3_9[15],stage3_8[21],stage3_7[29]}
   );
   gpc606_5 gpc966 (
      {stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[11],stage3_9[16],stage3_8[22],stage3_7[30]}
   );
   gpc606_5 gpc967 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[12],stage3_9[17],stage3_8[23],stage3_7[31]}
   );
   gpc606_5 gpc968 (
      {stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[13],stage3_9[18],stage3_8[24],stage3_7[32]}
   );
   gpc615_5 gpc969 (
      {stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[60]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[14],stage3_9[19],stage3_8[25],stage3_7[33]}
   );
   gpc615_5 gpc970 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73]},
      {stage2_8[61]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[15],stage3_9[20],stage3_8[26],stage3_7[34]}
   );
   gpc615_5 gpc971 (
      {stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78]},
      {stage2_8[62]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[16],stage3_9[21],stage3_8[27],stage3_7[35]}
   );
   gpc615_5 gpc972 (
      {stage2_7[79], stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83]},
      {stage2_8[63]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[17],stage3_9[22],stage3_8[28],stage3_7[36]}
   );
   gpc615_5 gpc973 (
      {stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87], stage2_7[88]},
      {stage2_8[64]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[18],stage3_9[23],stage3_8[29],stage3_7[37]}
   );
   gpc606_5 gpc974 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[9],stage3_10[19],stage3_9[24],stage3_8[30]}
   );
   gpc1163_5 gpc975 (
      {stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[1],stage3_11[10],stage3_10[20],stage3_9[25]}
   );
   gpc1163_5 gpc976 (
      {stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[1]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[2],stage3_11[11],stage3_10[21],stage3_9[26]}
   );
   gpc1163_5 gpc977 (
      {stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[2]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[3],stage3_11[12],stage3_10[22],stage3_9[27]}
   );
   gpc1163_5 gpc978 (
      {stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[3]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[4],stage3_11[13],stage3_10[23],stage3_9[28]}
   );
   gpc615_5 gpc979 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70]},
      {stage2_10[30]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[4],stage3_12[5],stage3_11[14],stage3_10[24],stage3_9[29]}
   );
   gpc615_5 gpc980 (
      {stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75]},
      {stage2_10[31]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[5],stage3_12[6],stage3_11[15],stage3_10[25],stage3_9[30]}
   );
   gpc615_5 gpc981 (
      {stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_10[32]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[6],stage3_12[7],stage3_11[16],stage3_10[26],stage3_9[31]}
   );
   gpc606_5 gpc982 (
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage3_14[0],stage3_13[7],stage3_12[8],stage3_11[17],stage3_10[27]}
   );
   gpc606_5 gpc983 (
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15]},
      {stage3_14[1],stage3_13[8],stage3_12[9],stage3_11[18],stage3_10[28]}
   );
   gpc606_5 gpc984 (
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21]},
      {stage3_14[2],stage3_13[9],stage3_12[10],stage3_11[19],stage3_10[29]}
   );
   gpc606_5 gpc985 (
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage3_14[3],stage3_13[10],stage3_12[11],stage3_11[20],stage3_10[30]}
   );
   gpc606_5 gpc986 (
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33]},
      {stage3_14[4],stage3_13[11],stage3_12[12],stage3_11[21],stage3_10[31]}
   );
   gpc606_5 gpc987 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67], stage2_10[68]},
      {stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39]},
      {stage3_14[5],stage3_13[12],stage3_12[13],stage3_11[22],stage3_10[32]}
   );
   gpc606_5 gpc988 (
      {stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72], stage2_10[73], stage2_10[74]},
      {stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45]},
      {stage3_14[6],stage3_13[13],stage3_12[14],stage3_11[23],stage3_10[33]}
   );
   gpc606_5 gpc989 (
      {stage2_10[75], stage2_10[76], stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80]},
      {stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51]},
      {stage3_14[7],stage3_13[14],stage3_12[15],stage3_11[24],stage3_10[34]}
   );
   gpc606_5 gpc990 (
      {stage2_10[81], stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57]},
      {stage3_14[8],stage3_13[15],stage3_12[16],stage3_11[25],stage3_10[35]}
   );
   gpc606_5 gpc991 (
      {stage2_10[87], stage2_10[88], stage2_10[89], stage2_10[90], stage2_10[91], stage2_10[92]},
      {stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage3_14[9],stage3_13[16],stage3_12[17],stage3_11[26],stage3_10[36]}
   );
   gpc606_5 gpc992 (
      {stage2_10[93], stage2_10[94], stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98]},
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69]},
      {stage3_14[10],stage3_13[17],stage3_12[18],stage3_11[27],stage3_10[37]}
   );
   gpc606_5 gpc993 (
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[18],stage3_12[19],stage3_11[28]}
   );
   gpc606_5 gpc994 (
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[19],stage3_12[20],stage3_11[29]}
   );
   gpc606_5 gpc995 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[20],stage3_12[21],stage3_11[30]}
   );
   gpc606_5 gpc996 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[21],stage3_12[22],stage3_11[31]}
   );
   gpc606_5 gpc997 (
      {stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[22],stage3_12[23],stage3_11[32]}
   );
   gpc606_5 gpc998 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[23],stage3_12[24],stage3_11[33]}
   );
   gpc615_5 gpc999 (
      {stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_12[70]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[24],stage3_12[25],stage3_11[34]}
   );
   gpc606_5 gpc1000 (
      {stage2_12[71], stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[18],stage3_13[25],stage3_12[26]}
   );
   gpc606_5 gpc1001 (
      {stage2_12[77], stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[19],stage3_13[26],stage3_12[27]}
   );
   gpc606_5 gpc1002 (
      {stage2_12[83], stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[20],stage3_13[27],stage3_12[28]}
   );
   gpc606_5 gpc1003 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[21],stage3_13[28],stage3_12[29]}
   );
   gpc606_5 gpc1004 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[11],stage3_14[22],stage3_13[29]}
   );
   gpc1_1 gpc1005 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1006 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1007 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1008 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1009 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1010 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1011 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1012 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1013 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1014 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1015 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1016 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1017 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1018 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1019 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1020 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc1021 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc1022 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc1023 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc1024 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc1025 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc1026 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc1027 (
      {stage2_1[54]},
      {stage3_1[22]}
   );
   gpc1_1 gpc1028 (
      {stage2_1[55]},
      {stage3_1[23]}
   );
   gpc1_1 gpc1029 (
      {stage2_1[56]},
      {stage3_1[24]}
   );
   gpc1_1 gpc1030 (
      {stage2_1[57]},
      {stage3_1[25]}
   );
   gpc1_1 gpc1031 (
      {stage2_4[86]},
      {stage3_4[31]}
   );
   gpc1_1 gpc1032 (
      {stage2_4[87]},
      {stage3_4[32]}
   );
   gpc1_1 gpc1033 (
      {stage2_4[88]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1034 (
      {stage2_6[89]},
      {stage3_6[36]}
   );
   gpc1_1 gpc1035 (
      {stage2_6[90]},
      {stage3_6[37]}
   );
   gpc1_1 gpc1036 (
      {stage2_6[91]},
      {stage3_6[38]}
   );
   gpc1_1 gpc1037 (
      {stage2_6[92]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1038 (
      {stage2_6[93]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1039 (
      {stage2_6[94]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1040 (
      {stage2_6[95]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1041 (
      {stage2_6[96]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1042 (
      {stage2_6[97]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1043 (
      {stage2_9[81]},
      {stage3_9[32]}
   );
   gpc1_1 gpc1044 (
      {stage2_9[82]},
      {stage3_9[33]}
   );
   gpc1_1 gpc1045 (
      {stage2_9[83]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1046 (
      {stage2_9[84]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1047 (
      {stage2_9[85]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1048 (
      {stage2_9[86]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1049 (
      {stage2_9[87]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1050 (
      {stage2_9[88]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1051 (
      {stage2_9[89]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1052 (
      {stage2_9[90]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1053 (
      {stage2_9[91]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1054 (
      {stage2_11[63]},
      {stage3_11[35]}
   );
   gpc1_1 gpc1055 (
      {stage2_11[64]},
      {stage3_11[36]}
   );
   gpc1_1 gpc1056 (
      {stage2_11[65]},
      {stage3_11[37]}
   );
   gpc1_1 gpc1057 (
      {stage2_11[66]},
      {stage3_11[38]}
   );
   gpc1_1 gpc1058 (
      {stage2_11[67]},
      {stage3_11[39]}
   );
   gpc1_1 gpc1059 (
      {stage2_11[68]},
      {stage3_11[40]}
   );
   gpc1_1 gpc1060 (
      {stage2_11[69]},
      {stage3_11[41]}
   );
   gpc1_1 gpc1061 (
      {stage2_11[70]},
      {stage3_11[42]}
   );
   gpc1_1 gpc1062 (
      {stage2_11[71]},
      {stage3_11[43]}
   );
   gpc1_1 gpc1063 (
      {stage2_11[72]},
      {stage3_11[44]}
   );
   gpc1_1 gpc1064 (
      {stage2_11[73]},
      {stage3_11[45]}
   );
   gpc1_1 gpc1065 (
      {stage2_11[74]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1066 (
      {stage2_11[75]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1067 (
      {stage2_11[76]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1068 (
      {stage2_11[77]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1069 (
      {stage2_11[78]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1070 (
      {stage2_11[79]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1071 (
      {stage2_11[80]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1072 (
      {stage2_11[81]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1073 (
      {stage2_12[95]},
      {stage3_12[30]}
   );
   gpc1_1 gpc1074 (
      {stage2_12[96]},
      {stage3_12[31]}
   );
   gpc1_1 gpc1075 (
      {stage2_12[97]},
      {stage3_12[32]}
   );
   gpc1_1 gpc1076 (
      {stage2_12[98]},
      {stage3_12[33]}
   );
   gpc1_1 gpc1077 (
      {stage2_12[99]},
      {stage3_12[34]}
   );
   gpc1_1 gpc1078 (
      {stage2_12[100]},
      {stage3_12[35]}
   );
   gpc1_1 gpc1079 (
      {stage2_12[101]},
      {stage3_12[36]}
   );
   gpc1_1 gpc1080 (
      {stage2_12[102]},
      {stage3_12[37]}
   );
   gpc1_1 gpc1081 (
      {stage2_12[103]},
      {stage3_12[38]}
   );
   gpc1_1 gpc1082 (
      {stage2_12[104]},
      {stage3_12[39]}
   );
   gpc1_1 gpc1083 (
      {stage2_12[105]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1084 (
      {stage2_12[106]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1085 (
      {stage2_12[107]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1086 (
      {stage2_12[108]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1087 (
      {stage2_12[109]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1088 (
      {stage2_12[110]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1089 (
      {stage2_12[111]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1090 (
      {stage2_13[48]},
      {stage3_13[30]}
   );
   gpc1_1 gpc1091 (
      {stage2_13[49]},
      {stage3_13[31]}
   );
   gpc1_1 gpc1092 (
      {stage2_13[50]},
      {stage3_13[32]}
   );
   gpc1_1 gpc1093 (
      {stage2_13[51]},
      {stage3_13[33]}
   );
   gpc1_1 gpc1094 (
      {stage2_14[24]},
      {stage3_14[23]}
   );
   gpc1_1 gpc1095 (
      {stage2_14[25]},
      {stage3_14[24]}
   );
   gpc1_1 gpc1096 (
      {stage2_14[26]},
      {stage3_14[25]}
   );
   gpc1_1 gpc1097 (
      {stage2_15[6]},
      {stage3_15[12]}
   );
   gpc1_1 gpc1098 (
      {stage2_15[7]},
      {stage3_15[13]}
   );
   gpc1_1 gpc1099 (
      {stage2_15[8]},
      {stage3_15[14]}
   );
   gpc1_1 gpc1100 (
      {stage2_15[9]},
      {stage3_15[15]}
   );
   gpc1_1 gpc1101 (
      {stage2_15[10]},
      {stage3_15[16]}
   );
   gpc1_1 gpc1102 (
      {stage2_15[11]},
      {stage3_15[17]}
   );
   gpc606_5 gpc1103 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1104 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc1105 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1106 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1107 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[18]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc615_5 gpc1108 (
      {stage3_2[11], stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15]},
      {stage3_3[19]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc1109 (
      {stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc606_5 gpc1110 (
      {stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[3],stage4_5[6],stage4_4[7]}
   );
   gpc606_5 gpc1111 (
      {stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[4],stage4_5[7],stage4_4[8]}
   );
   gpc606_5 gpc1112 (
      {stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[3],stage4_6[5],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc1113 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[4],stage4_6[6],stage4_5[9]}
   );
   gpc606_5 gpc1114 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[5],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc1115 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[6],stage4_6[8],stage4_5[11]}
   );
   gpc606_5 gpc1116 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[6],stage4_7[7],stage4_6[9],stage4_5[12]}
   );
   gpc606_5 gpc1117 (
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[7],stage4_7[8],stage4_6[10]}
   );
   gpc615_5 gpc1118 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[8],stage4_7[9],stage4_6[11]}
   );
   gpc615_5 gpc1119 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[25]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[9],stage4_7[10],stage4_6[12]}
   );
   gpc615_5 gpc1120 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[26]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[10],stage4_7[11],stage4_6[13]}
   );
   gpc615_5 gpc1121 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[27]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[11],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1122 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[30]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[5],stage4_9[9],stage4_8[12],stage4_7[13]}
   );
   gpc606_5 gpc1123 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[6],stage4_9[10]}
   );
   gpc606_5 gpc1124 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[2],stage4_10[7],stage4_9[11]}
   );
   gpc606_5 gpc1125 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[3],stage4_10[8],stage4_9[12]}
   );
   gpc606_5 gpc1126 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[4],stage4_10[9],stage4_9[13]}
   );
   gpc606_5 gpc1127 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[4],stage4_11[5],stage4_10[10],stage4_9[14]}
   );
   gpc606_5 gpc1128 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[5],stage4_11[6],stage4_10[11],stage4_9[15]}
   );
   gpc2135_5 gpc1129 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[6],stage4_12[6],stage4_11[7],stage4_10[12]}
   );
   gpc2135_5 gpc1130 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[1]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[1],stage4_13[7],stage4_12[7],stage4_11[8],stage4_10[13]}
   );
   gpc2135_5 gpc1131 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[42], stage3_11[43], stage3_11[44]},
      {stage3_12[2]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[2],stage4_13[8],stage4_12[8],stage4_11[9],stage4_10[14]}
   );
   gpc2135_5 gpc1132 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage3_12[3]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[3],stage4_13[9],stage4_12[9],stage4_11[10],stage4_10[15]}
   );
   gpc606_5 gpc1133 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage4_14[4],stage4_13[10],stage4_12[10],stage4_11[11],stage4_10[16]}
   );
   gpc606_5 gpc1134 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage4_14[5],stage4_13[11],stage4_12[11],stage4_11[12],stage4_10[17]}
   );
   gpc606_5 gpc1135 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[16], stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21]},
      {stage4_14[6],stage4_13[12],stage4_12[12],stage4_11[13],stage4_10[18]}
   );
   gpc615_5 gpc1136 (
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_12[22]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[7],stage4_13[13],stage4_12[13],stage4_11[14]}
   );
   gpc606_5 gpc1137 (
      {stage3_12[23], stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[8],stage4_13[14],stage4_12[14]}
   );
   gpc606_5 gpc1138 (
      {stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[2],stage4_14[9],stage4_13[15],stage4_12[15]}
   );
   gpc606_5 gpc1139 (
      {stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[3],stage4_14[10],stage4_13[16],stage4_12[16]}
   );
   gpc606_5 gpc1140 (
      {stage3_12[41], stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[4],stage4_14[11],stage4_13[17],stage4_12[17]}
   );
   gpc606_5 gpc1141 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[4],stage4_15[5],stage4_14[12],stage4_13[18]}
   );
   gpc606_5 gpc1142 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[5],stage4_15[6],stage4_14[13],stage4_13[19]}
   );
   gpc606_5 gpc1143 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[6],stage4_15[7],stage4_14[14],stage4_13[20]}
   );
   gpc1_1 gpc1144 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1145 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1146 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1147 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1148 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1149 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1150 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1151 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1152 (
      {stage3_1[18]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1153 (
      {stage3_1[19]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1154 (
      {stage3_1[20]},
      {stage4_1[6]}
   );
   gpc1_1 gpc1155 (
      {stage3_1[21]},
      {stage4_1[7]}
   );
   gpc1_1 gpc1156 (
      {stage3_1[22]},
      {stage4_1[8]}
   );
   gpc1_1 gpc1157 (
      {stage3_1[23]},
      {stage4_1[9]}
   );
   gpc1_1 gpc1158 (
      {stage3_1[24]},
      {stage4_1[10]}
   );
   gpc1_1 gpc1159 (
      {stage3_1[25]},
      {stage4_1[11]}
   );
   gpc1_1 gpc1160 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1161 (
      {stage3_4[31]},
      {stage4_4[10]}
   );
   gpc1_1 gpc1162 (
      {stage3_4[32]},
      {stage4_4[11]}
   );
   gpc1_1 gpc1163 (
      {stage3_4[33]},
      {stage4_4[12]}
   );
   gpc1_1 gpc1164 (
      {stage3_5[30]},
      {stage4_5[13]}
   );
   gpc1_1 gpc1165 (
      {stage3_5[31]},
      {stage4_5[14]}
   );
   gpc1_1 gpc1166 (
      {stage3_6[44]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1167 (
      {stage3_7[33]},
      {stage4_7[14]}
   );
   gpc1_1 gpc1168 (
      {stage3_7[34]},
      {stage4_7[15]}
   );
   gpc1_1 gpc1169 (
      {stage3_7[35]},
      {stage4_7[16]}
   );
   gpc1_1 gpc1170 (
      {stage3_7[36]},
      {stage4_7[17]}
   );
   gpc1_1 gpc1171 (
      {stage3_7[37]},
      {stage4_7[18]}
   );
   gpc1_1 gpc1172 (
      {stage3_9[42]},
      {stage4_9[16]}
   );
   gpc1_1 gpc1173 (
      {stage3_11[53]},
      {stage4_11[15]}
   );
   gpc1_1 gpc1174 (
      {stage3_13[32]},
      {stage4_13[21]}
   );
   gpc1_1 gpc1175 (
      {stage3_13[33]},
      {stage4_13[22]}
   );
   gpc1_1 gpc1176 (
      {stage3_14[24]},
      {stage4_14[15]}
   );
   gpc1_1 gpc1177 (
      {stage3_14[25]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1178 (
      {stage3_16[0]},
      {stage4_16[7]}
   );
   gpc1_1 gpc1179 (
      {stage3_16[1]},
      {stage4_16[8]}
   );
   gpc1_1 gpc1180 (
      {stage3_16[2]},
      {stage4_16[9]}
   );
   gpc1_1 gpc1181 (
      {stage3_16[3]},
      {stage4_16[10]}
   );
   gpc1_1 gpc1182 (
      {stage3_16[4]},
      {stage4_16[11]}
   );
   gpc1_1 gpc1183 (
      {stage3_17[0]},
      {stage4_17[3]}
   );
   gpc1163_5 gpc1184 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[0]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc623_5 gpc1185 (
      {stage4_2[1], stage4_2[2], stage4_2[3]},
      {stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc606_5 gpc1186 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc1187 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2]}
   );
   gpc615_5 gpc1188 (
      {stage4_5[5], stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9]},
      {stage4_6[7]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc615_5 gpc1189 (
      {stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[8]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc1190 (
      {stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13], stage4_6[14]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[4],stage5_6[5]}
   );
   gpc2135_5 gpc1191 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[4]}
   );
   gpc2135_5 gpc1192 (
      {stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2],stage5_9[5]}
   );
   gpc7_3 gpc1193 (
      {stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16]},
      {stage5_11[2],stage5_10[3],stage5_9[6]}
   );
   gpc2135_5 gpc1194 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[2], stage4_11[3], stage4_11[4]},
      {stage4_12[4]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[3],stage5_10[4]}
   );
   gpc606_5 gpc1195 (
      {stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16]},
      {stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[4],stage5_10[5]}
   );
   gpc615_5 gpc1196 (
      {stage4_11[5], stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9]},
      {stage4_12[11]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[2],stage5_13[4],stage5_12[4],stage5_11[5]}
   );
   gpc615_5 gpc1197 (
      {stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13], stage4_11[14]},
      {stage4_12[12]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[3],stage5_13[5],stage5_12[5],stage5_11[6]}
   );
   gpc606_5 gpc1198 (
      {stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17], 1'b0},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[2],stage5_14[4],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1199 (
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[3],stage5_14[5],stage5_13[7]}
   );
   gpc606_5 gpc1200 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[2],stage5_15[4],stage5_14[6]}
   );
   gpc615_5 gpc1201 (
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16]},
      {stage4_15[6]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[2],stage5_16[3],stage5_15[5],stage5_14[7]}
   );
   gpc1_1 gpc1202 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1203 (
      {stage4_0[4]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1204 (
      {stage4_0[5]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1205 (
      {stage4_0[6]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1206 (
      {stage4_0[7]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1207 (
      {stage4_0[8]},
      {stage5_0[6]}
   );
   gpc1_1 gpc1208 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1209 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1210 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1211 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc1212 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc1213 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc1214 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1215 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1216 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1217 (
      {stage4_3[3]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1218 (
      {stage4_3[4]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1219 (
      {stage4_3[5]},
      {stage5_3[4]}
   );
   gpc1_1 gpc1220 (
      {stage4_3[6]},
      {stage5_3[5]}
   );
   gpc1_1 gpc1221 (
      {stage4_4[12]},
      {stage5_4[3]}
   );
   gpc1_1 gpc1222 (
      {stage4_6[15]},
      {stage5_6[6]}
   );
   gpc1_1 gpc1223 (
      {stage4_7[18]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1224 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc1225 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc1226 (
      {stage4_8[8]},
      {stage5_8[7]}
   );
   gpc1_1 gpc1227 (
      {stage4_8[9]},
      {stage5_8[8]}
   );
   gpc1_1 gpc1228 (
      {stage4_8[10]},
      {stage5_8[9]}
   );
   gpc1_1 gpc1229 (
      {stage4_8[11]},
      {stage5_8[10]}
   );
   gpc1_1 gpc1230 (
      {stage4_8[12]},
      {stage5_8[11]}
   );
   gpc1_1 gpc1231 (
      {stage4_10[17]},
      {stage5_10[6]}
   );
   gpc1_1 gpc1232 (
      {stage4_10[18]},
      {stage5_10[7]}
   );
   gpc1_1 gpc1233 (
      {stage4_11[15]},
      {stage5_11[7]}
   );
   gpc1_1 gpc1234 (
      {stage4_13[20]},
      {stage5_13[8]}
   );
   gpc1_1 gpc1235 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc1236 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc1237 (
      {stage4_15[7]},
      {stage5_15[6]}
   );
   gpc1_1 gpc1238 (
      {stage4_17[0]},
      {stage5_17[3]}
   );
   gpc1_1 gpc1239 (
      {stage4_17[1]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1240 (
      {stage4_17[2]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1241 (
      {stage4_17[3]},
      {stage5_17[6]}
   );
   gpc117_4 gpc1242 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4], stage5_0[5], stage5_0[6]},
      {stage5_1[0]},
      {stage5_2[0]},
      {stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc215_4 gpc1243 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0]}
   );
   gpc615_5 gpc1244 (
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc623_5 gpc1245 (
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc1246 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[2]}
   );
   gpc615_5 gpc1247 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[3]}
   );
   gpc1163_5 gpc1248 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc615_5 gpc1249 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6]},
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6]},
      {stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[3],stage6_13[3]}
   );
   gpc1163_5 gpc1250 (
      {stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[0]},
      {1'b0},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[2]}
   );
   gpc1_1 gpc1251 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1252 (
      {stage5_1[2]},
      {stage6_1[2]}
   );
   gpc1_1 gpc1253 (
      {stage5_1[3]},
      {stage6_1[3]}
   );
   gpc1_1 gpc1254 (
      {stage5_1[4]},
      {stage6_1[4]}
   );
   gpc1_1 gpc1255 (
      {stage5_1[5]},
      {stage6_1[5]}
   );
   gpc1_1 gpc1256 (
      {stage5_1[6]},
      {stage6_1[6]}
   );
   gpc1_1 gpc1257 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1258 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc1259 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc1260 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc1261 (
      {stage5_3[0]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1262 (
      {stage5_3[1]},
      {stage6_3[2]}
   );
   gpc1_1 gpc1263 (
      {stage5_3[2]},
      {stage6_3[3]}
   );
   gpc1_1 gpc1264 (
      {stage5_3[3]},
      {stage6_3[4]}
   );
   gpc1_1 gpc1265 (
      {stage5_3[4]},
      {stage6_3[5]}
   );
   gpc1_1 gpc1266 (
      {stage5_3[5]},
      {stage6_3[6]}
   );
   gpc1_1 gpc1267 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc1268 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1269 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc1270 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc1271 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc1272 (
      {stage5_8[8]},
      {stage6_8[3]}
   );
   gpc1_1 gpc1273 (
      {stage5_8[9]},
      {stage6_8[4]}
   );
   gpc1_1 gpc1274 (
      {stage5_8[10]},
      {stage6_8[5]}
   );
   gpc1_1 gpc1275 (
      {stage5_8[11]},
      {stage6_8[6]}
   );
   gpc1_1 gpc1276 (
      {stage5_9[6]},
      {stage6_9[2]}
   );
   gpc1_1 gpc1277 (
      {stage5_11[7]},
      {stage6_11[3]}
   );
   gpc1_1 gpc1278 (
      {stage5_13[9]},
      {stage6_13[4]}
   );
   gpc1_1 gpc1279 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc1280 (
      {stage5_14[7]},
      {stage6_14[4]}
   );
   gpc1_1 gpc1281 (
      {stage5_17[6]},
      {stage6_17[3]}
   );
   gpc1_1 gpc1282 (
      {stage5_18[1]},
      {stage6_18[1]}
   );
   gpc606_5 gpc1283 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], stage6_1[5]},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc1415_5 gpc1284 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[6]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[1],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc623_5 gpc1285 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc1343_5 gpc1286 (
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc207_4 gpc1287 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], 1'b0},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc1406_5 gpc1288 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], 1'b0},
      {stage6_16[0], stage6_16[1], stage6_16[2], 1'b0},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc135_4 gpc1289 (
      {stage6_17[1], stage6_17[2], stage6_17[3], 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], 1'b0},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1_1 gpc1290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc1291 (
      {stage6_1[6]},
      {stage7_1[1]}
   );
   gpc1_1 gpc1292 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc1293 (
      {stage6_8[6]},
      {stage7_8[1]}
   );
   gpc1_1 gpc1294 (
      {stage6_11[3]},
      {stage7_11[1]}
   );
   gpc1_1 gpc1295 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
   gpc1_1 gpc1296 (
      {stage6_20[0]},
      {stage7_20[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor_CLA486_12 compressor_CLA486_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h75deb16be95f29af5978f4b36bd4320e1048cb76ba3062ee26cbde02dec159e62cdf93ab8f641675354d9a676612119e61a792031d1551ff66162fd78d0fce038a3041fa23a8d6ece655fa23391f7b4c037700812b5092330bc4dfb8c581932b0aa0e08464fc908ee5fcb1d2382b67787bfdf6cef8d19c7d270bd843d4647a29a083c33f29388cffab2d333af4357afdbe075aaded2d925a72c5c90d650f39dfebc1c89c3e0b13f807d66ddf07f8cb15d78b0607cc3723186fa4b7e79ffa0339f829acc688160ec180d40e799359518c9350dca7ebf2c198011a178c8f118b1e32a89193f3bbdb9ca7772097da396a47d6042fecafcf0c72ca870d16b6a819649d7d4af2f78e12ae5b8b84d6cea9d79970984f0096c03907f584374896a35f200efe5a5fc24a56d0cc393a515c48a0202e6ded054c2da8d36ffc3aa2838eb30623e8ce1a0b900ca0b2793890e58a0043c8a95852e20ddab3c2b0d5629585896878e99df6132bcee72f01123790d23c7b0050b6a5a6b66f9e57b32908cc6326b1d5ec9512b870f5bb3b38b2100ac495f1f91bbe82250500634feb18928b39268297fadc4e644f5bfff88f5e007f9312612d177462acbe763a4060b0efad995e678a91a5ddcab9cbfc3394ce85069f666aaf909889134d1fe62936eb30c264b4cd88b0f97a2c226eaea70e311f3bfb78e97f7283c1b1d50ce4d99e10da58f43d588aea334f92ff3c50cabd43eec42b8ce02ea5398c615addaf2aba536dab29f01bb2cb240b6f0f6113c6ac0d57bc14452a108c4fe12100cc4c280799a6ef347b6a401e31c019e8130352fbfea1978f6eea2a10fe02f0f432a2ce66c61960329a993fd6fc086364a0c7973471434891de6aeb25bef3732ccacf36b9708af4048b63038d45c2e1bb1f33734fa35e5a706ad5b864f92a94472814e026f2851d7feff8d0a5e59caa0bb8bd6f962bd5eeaa23cf7bfce3f9a098c3fd0674d417354489dbadab9912ad1eb0531e1a26f00467b50a03e917618fc5908d95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h26c94de0c0044c1beb591415bf3579600cd3bfe4ce5f1278315f2bc3e5039e1b88243fb28c468a8415ffa59996b1e0c3a82d421e3f0ee0e4c3a28a05a5a8e9600fab6372875f4c7758fd33299c72e87d1ec87c879282a5412f8557651ef1e5d5cc7adbb941e5f0976d730553bbfda0d98969131f9d89de1622c1ab87e92c12b4bd30121e681a90955109cd5765433afa0a379103775300e050dff1177f730992946a2229e641a31a754fe45b3ccece6afc46d790a76d63cfb2045dd8080bb4a00f65516f4d0a35b708e6b74ab2e49c5da3be160fd54579ce1714ff6be78b02bffd658635d82f0048ac4c4039c1a0701e5a00c38acca999d845aa6e98eb209300c287c8b525a2779aac7db1eaea3244062d589ffa4979aa934be890dd872508e40db061c486eb5b7b1e87ce1363b859d292b4714d804ffea7535f0121a37e9916d03ed7424355de5d11feca433bc06b7f1551ed2127100c948ef580d739c204557a9f27ef1379ee8549708a45b43611567628206da9abdd6e65196719dff1a4379f07b1c6010308da6c0ab3e69269c3221c1d777ae2a4b1b0e28a3871be9d8466893a745f1d5f973964c033fe7999df3909d293b03e26240700b5c132a7e4eabc05f8ccd32d78ee66c8603ff2f09f77866d251b4e7255dc7b329ec01e7c4c0aafe9515b689832a9d745d7d86eb6ad4f6f3567a5ac79446e7cedd04e7d9b716ff3838c40dd1a8acf15be1ff7bb94e652d07eae580f2ee2e2a8fd8d7af657f7e729f1ff0883cefde284a26c1854fd3933199e9b0e21c8926b4477c7a427473600474968368175f6c7d7132a9109bea95c791d2b230c3cd267f5f5a22eaa82b95f810d9d4473d0fc0c68e5b5517684c6428552c44c943fe644c6a1fb8bed2a81b9bc248ec08dc3c23ccfe49b3c07937c130db85abb44f9972074176187d6d6b8161c5f09a3c15c0328ea723b8d064f6b31e5d6f4279741c8b121d0490bc24dfaaeb98ac61c7e19cdb69f1ab66f75bbd8584b9ac2d0678fafc39c25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1185bd2f5147e8f9d2c2fdaa0b7a64990abc94a348abfdc7855810a8427348388c9d8df1206a2eed95bacad48c2f04eb8d2c6f8cc74085e812ec23d985779942097c44999fa542a78bc2ab56b5f69321f9632e57aeabec2656386b554895762d04fda47ba137a248c2f8ac06043b25bce3302300abaa5f082f47e02896771821a0faa1f3c852e613871b7368b7229cb3f6f609e1fedc937121d03e62f514ddc272671ac2f63dcd11c04301f4e5d68f44482ba06a7b73dc8033d881d4e4cde9c8d3b5b34a1f7f9eb8cf4931829edb502d2db697437c749f6b572cd2c8e5ee91377739ced91a46707fe1eede157af8d676e176d65ce0965cd877b9fe5ae4f12802b62e6c8a181f8cf61a49fbfbddd807fca609365eb9da508e468576239d747212fb7c8e97cd03cb7a729a49aaa5fea391e68161651e6152045a91595303afb4392849d0681438c473dfa201e9b5c3d4bbb82ce249760ddcd5551932a4c1ea108d630ff97c93e79dbdcdb325f950a9679682598cf71fef6464f245f522502a465e8b2428c4ea085ed80a99e14ed38a99f5b23d5f224ba8e7eb30ed0727ef90d4e61cef8d28c959905ec4c456b2d653ea8d103bdb1137793954277c855a048ab49c7476299a88f30f5e686f0b8521ab4b33bc3831247a2ffe26769f93fc974af091fc90e4091f06cce48f1fedee93fbcfb174c0e92088bb3eae288ab91f14593a71d36bc67603840fe4b6d16b95e4d85b1d4f0763b4249cceb1785c609124496bd4a3b2638b52ac0e743d7750debd66e641d5115a2f2404a9e41489399ccb06f698d49cf94302bda8629c571da311d0379242d3e1ee26b1ce121d2a7f4c30aa0711be309ee0faaa30980f0daa8e46af7cea9b15ff0993e9fe896f4b012cd568637c2ef21e229cf97453679609a4b34c4532fdf10ef11bb812a0ba965801da8d7b367dac1b70ec8b1018fba264ab3929f2b4918b0db748ebd374b62919bcd970bf013fbcc601273f5f2554f29560f5c00d4b25a11f8014f919cb9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha4cd7c9685dfcc731e843b550cbbc5a205ca0c81f0cb86b77096a3f4d3c916785df323b15b8af1ea29645740b6e9072edd46b61978b48a30d7cd280c32ad9667a85d7be9f1011a39bf156fadf49be6abbcda47a22a542f24ce957a92ad74d2fd34669834a5022bb773f009d33ac21e2d330d0c2e5fd2b4f4dabfa6d6630774999417028dceb3cea03d16f76deca3cba228709f5f9ba91c65d88643f356a5a1f9b133e7add5231b04de59587d123f6f707a75be060aee958cff4b87d4f928c4c96dd90433cd96af428c606291d609a0d7d3ff7aad1185cca9300a8b5488e3d9c271602d81cbd58e93af2cf9bc40c26162a2b3a8579d18ffe0dcf335331e8c1a277c79fb02c41f0c43317589aca672c82e3a6ed616f84594aa0fbc48292a49fe7cb649ba8e2bf7ad8d140a18db6f5a71bec6beb9f04dd752008ffa439ef5964b27d5489fcf1babd5c2ad0007d016ebe55ac9b9e5207397a9d1f2fb5d537506616717bc08115304d9a55ac991e9c67bb0b3165d056f5974727a5e2e6884274c5e0608ebf8180a48cefc3cfd4f22b0de78db67b9f65b3fc28297c53596f06ebde6581f3ba0f244e67fa390c42df0537dd315106edf4e4a90f3d11b19966670a0c57a279c4471727e34315ad3d0ec825e9409ed15b58fe5a46bd962779a1f0d9758387341abab8f88b8cf62dea54f27a33d0a3fa034e672f18fb5bbe8bc099b3254810881e458efe8815c77566f57fad808bd12da442d5a2f29a2ca85b9e983c031433777ff5fff6cfd7f7a5317944b4a22a2edfe789ceda83f20f25ac6009eb5f9c02f37dfb1aa2a35ab26a5d264e128d447eb87466705b33797aa74f9b6ee1f2640de40c592203495e5ac3c316c14dd5668c18d1c4a8e4d453a99a61a851e0964662c67bb5031204d61f85561b286930b587f264d7bbb148e3390f37edadb18e49ac3ba8c49511f0223e721a47ed6af5d0901c26c84566a84b66e9548e7748eb23477d130fe6b196c5bf9e80ebea57ad27e10ec3348bb28d51f42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h24c01f0855dc57dbcfda91670ec88c216c5937d6e4e5567b8a10c673798368000b1e886f007f664b41366f3ced66cccf3e11706f5da3b72796ac310108c5689cdf63955671b0d6cfd9978c866cf3efe42c60293bd5386d39aaf6f52f7f29ac17a51b54cf3579917c866b0485c77ef27bc1116140d927278a2b569bf8fcd10a6e54ee376308757471b191de9017652a1614b41e9e7c1e2d66260204e3928e65faa6f30afe29ccc075dc5499fbaeb36c7c7a2bf721330ddb62e9574f5fcd9763bfc41ef5f7f94da24c29f5a8fb9450bb387c8d125f75ad17086961005b16e09978370b066749d8ab9267605dee45b6ebf28e04e81d82b9a43734f3500e79e867467920515c6fa46736ddb4c3dac7290f905132031e91fc17564e291dea79df40f6a9589aa40987042ce2f5cd9180e9b8a08771098a921faf5a4946e2caeb1c225286b4bdbbc3e0008659893554023dd07872449f7dc2f2dcdd6d906177cad551434a2d85ec5a6e5ff38e828360f78b1405ec458a7ff4d70bb8df0eaa6253329d4a41f98842d20f421a0a40a58e9acdf420753877ce8b6f26adf42db110344f85e80316337bd3bde297e055e8d2f47186521b56307095cf9b84b997f73af102a06a2f69f5a1f4183450b3d0923281d890c9bb31c597484d74741e5e838e7102910c8621f61b73ae24abd4cd5205896364742591a460e521714ebc7dcb3a602d5a6a06b1b223cf2398fadb459ddc573951e0a6ba8201a251098ecd440fffb08dd7760639c1ac5299b168c3fe7e5cce25c093f0c6ddb870de2da5d89995a680f190180601884d95b2465538d8cf631f20430bf3f794d0a4f6b11faf60645340dcda42485ba980aa3202d2e2644de618ca6bf4e97d8e487a32473be87bd56a79f8893c35f85106ddf5398fadd4462a0bca4e804d42ee0626ed2926172629b53287bde8b4456bd7d3f1fbb729fdd999865051b8ce022fa0ff2300c546f9b77b6c10cf1d057393e927ae83751cb0a7538631b49643174ad63eda7062e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha4b96ea633baa0c82ab5db7207f01b56c027d88593079de07a988dbf7556cd39e0153d34692bba67140d9f853865bc1e47473415fd54446e2bb6431b096c4b698b0a755670ec7aa32981cf6043089c893587e2d31bf40ad2bbbf58503250df85629d322dce58a5d3076129f068e61d99b823f39a403e4937180a7b81f659a78b2f80450e6285680a182b395a8bbb7f3b0aca597c094d628ca20b9a7ea0de3a3812c23b695d651445b75d4508d3bfeef52d088d9f258eeac96e6234c0679e223680a7d8f12a8fadf36cd659c9c77dc4df6b7070163d6bf295ff5bc69b34de00b00c0c924c56a765550b2b7832f6529d3334e40427009a178ebc731e2e06c3de5296c6dee8c23a327d2ee15cb17644eed2d34450e0d0c604de1091026a7d35224176d46ea8122f89beacd800526b6467a61c1db7851e141a1f03e6409df60cadb2d0945dc2edbec78b6530c1589c383369392af8078b6650c458df27310d3c009c22333380503dad5385a95ee4de6a754710ec6d792c087f1ef6ef0902339784ae2908f235d4ec96ee16b3497756eb49f45078753520ace1088fa1bc793c224125fc3a6bb02ec041107b60adf6c45ebf3cb9221a1148dd83c6bc14146c0d3790686caeebab2103603f2b1c7d45aa4993d80f85cc97e6ba1207750734fc83dec50e01a06cafa816784659b1bdfecc2da4020a4b3be33c8ab58f42b1e3a0cd8138f188ee03e46ae15a8d02f6d73792553773632f9d269a7ddd22f7dde63df2832c9da8f0e19753526ffc5af15ac8692d19044346e2b786163d67631fae55217d2fb74c28c260382c43470b293bbd9ac23c8f4e8aa836f5124064882350183fbe67e5949b53814d6a50f87d885c44d37a3034658d62a884d67fb9d5f41767cb58edff01becda8d83481b5626aa60a33f1444f9ef13f1e8fd0ba46c8777f52889b2a65e86717cd0b07a96c6164133af15052bf1066a68ea95f1e7d98c6bc2ef8c5c16303ae17402292433f81b58d516c45e560498f88f7b6e8e18115;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2125caaf9061da7d24f103b728fd68c54865ac95e21a5f268adcb2ba9c1f5ebd3acf477d624eaf06c6c92a2aebdb8862b17117844a4fb213faccbcaeade5488ad3c776d438ee4530f99e0203fa8a1c0b9431f1ffc475520433c6adf4d9e609b3acc8833aeaa9587c83ab3f2d89e68322df66a71f6c444a1336ac2403516f10eee32f9c0bb53cf4bb842e897d55815a2c41beced2613fcbbf6bfd222431d405d3234ced3e53cd88b561e784152a436276f37160b62146f445a00c4e9d36bdae19ece3b508cdfcb3225b049282a43166db5c2f4340767ef190f117b08ca96bde716860208911ec993924a9af3e27f46fc4d1fcec3d192f12da081fa4fd036f1c3b13289cd5f122d4ff51d1674199c9f76ef9f1bbf6fd3deec437db8eb8163a14690f804d68b4ee7043ed0b99fae1c8475513c41e0cf3b136cdbe5d151a88f975c6e0ef927967c55b884993fa5d120d43e5e0cd98e5b9b071d3383ffb4805b7e24dd241576e54a259184e53b69ddae2f25367ec413d1f4623316dc60241babdb76cc14f215d4b625d34012af1ad2078d76ec649ed70ca161d960bc495f4171ef67c8ef63d409aa82c65934bfe21030bd2bb3ed74542067237d68a267dee727a09dc6fb691f97c1cb57387ead311ba5531b9f66fb1b550e5464b507176478da8252bb289e4c7309960b8c9af7602cbe7ce31a1dfd81cac4d160597c5168b2088cb0c17995ed93c34e063be2809df0fc51b03deb94a55235dd8dde579c2dd196e4a799f6a3b255787bda56cc0c6d840d842c91c7b6d059bbee408836715a93cc2002b9c27506f2fdce15e5a71eac9bf11c4f557b17015b07dc2e09a58f50b63a772faa8605d9674b8dc2980a9c478aee40dcd61376c5de27713619f11c7d0834ce46a6c2706b198a25745296cd552f613ef7a52c67aa5b13295630af766abc96a3eb2d344838b3036a679d4e86adeb20e5be8bab5c1a002b455ebadfd680124dc7a0af3219c8b5dec983f6151fbdf870cc0a77ca39868e8846e9b07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hdfc11e82334cb0d74ade47485e3495f3177b6ddca0189c2b7ea6a589f572c2d3c5bc08ddc437718635406712ed6e97fd947a5d2c75c0ba2921234cf3c53f1450a3eab928c4159379a4b4b2bf4ec09cc08c161dc612be0130a4e73eeddb95e5296e68e4772b0ecf12372d0bdae0d4b8edb99b3776a7f84e17abee9d0ba01d0df3348e80d9ef2e53e1a85132104c9a6f42011d20b02e36061cef828f9a960e45f51514511f94130b36d7f1838ab8fb8af1ca64fcb98d027f153be2bf64781b5db18b8e3358f18ac38e82146c1758e822c5ec091606f40d833e146f29cd61349dfd96f0678097968e7153c1cc5c0a5aea02d95a86ddca74e6d60ff12623b2b71d47d67497d876d66f5daf127b9ae230343ca05606861bdfe0fe83ff96ac270ff385d8b64e07c98342f5fa93849b459a107661684a7e8873e2d849e28ea1ace6353319b109248d4172d68b0b9bc03a98cbf425bfb64ad692576d11c9d20a44f55dbcd8ba5add15aea1b5e8ea25116a4634b471e1f5d0dc01c84721c44d926fc4d1739e63fad01edb49d3dede7f744d5fd29ef58f5a8de8fe71ab2b1c99ea3ba9b5c2d8183bb1f044e6323d12f5fdc1baf378901fdcfffc70841d2c69ad892d6dfa1bcffbea3a2511c9f9a6e640eed1ae08944bfe0d48a095e9aa83ef7d4154057096f33e332a2b637390461d111354b96b1998b98b32f4d626c554f6c785322d628a7dc11fe99220839f8c32837d2aeac9b1103178c586275264c4cdb4e2efa1adb2678b11679cd4cfbb0c2670aed1c118a05243d3a13b4d6445d5916d086e69b49f49d0e08f2385422a4c3cb3f679844f526e58e29a883583f86bf6c876c117ef2efd618169e8c0e658b19e837c6ae664bebd059cd00b271cc60552aafa2421dc7406ebb3003884e2f473059c52f7ff4221beb41cdac3a23564cbb29ed0983155c49f7cadb5e0658d5a449f6b02e8788c5e2df81786881617068633492c04389b702aa6bdb876f27a5cabd1560f87bb12fd984e9596b5b6a7cb1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h578b4c5d0232b13e0b4a1922936e85c46f70908d51eb78c8fe5d713bb50ddccc83ca9fdbb6124b29f3815123add3bffda4765db3e5c2c24e202c47ccb2279b11ea6d5c0c64632c6aaad45732cb225df91c904ba4f76626de78ac53918b6e26d9fd93a7ec10c409ca0610bdcfa85c06bb18142ee93b9af5beb69e9c8f7824d26e7287b4daa30b4d74779e7f4255ef393e1b22838a02bf9b8077ecae46b3ff2c8aa84c1be9d67653ce8c018c41b0542bacf4c912053120f0547e6963b6df27071580f40587cee3019f5b690992baac54066d36da45e9f1355a63610f9e9edaa5353eec2eb04529321f5b034ff1c60ab9a46a702e2f468a9f9fcea860566f7b735760f5b06611d190b0ef9e116f5e170a0b9fd7570253e3cd58bf95450fa65e3887511bf39ebad3bad57b0e8b8a38c6e439ff7fe931887eaae7f37308a308c67bc0f19ef655b38415cd508988c217b6f118bedd49ff86082be7aa02e8ada1a51bc4917dfeb67d1d21bdece724392fa0c2fe6ee1179ffbfe6f2c8c4b65b642490ac5da5d5f5ce5dbe46d05313d7b976f6d0394b48df3ff3f70b625ad1affe5632ee63b30c9983339a4f0307f57fd8c4d510271f0ddfa393f0c8ce9b39e582fed893705ff3c27c8a564d03f630bbf201187632ee0b9f644bc6da228da3c12f019997663b81210112907b19e29b2131a1a7975551a5463490ca36e5511b37bb2806bf74ca4d4a781ef2cf41b2a7f4b49874d59c503dee6adf617f03c8f1685f5ac60f175d074b26196c9374dbfaa39c082cb1c8f0a2b576b9eeb186f90504ec93dfda86caba0ddc2a69a88869b1a25c73003ac513ae24f552739dd82ae982aa3551a9fc44f3c1d2d81bdb3f9990a0a8c4a72a9cf93ae731eef818212bb7aad7150b343474cc04e13fe35f189ff795ccef72ff696c42c2f7865cefbd7ed53d3819f7f1dda4b76de546fa9e6bd469cf3d98de05cab64dbc3110f39743936ecb5b6717518f091ac7486de1f6003b0f962fda37bbd23d4909580a20ad5a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h46768181ce7000a2f8536c173abe513c72644dec5a287a9c72e7d451aa16809cf632368da1062bb75596da750981da10726bc6305b660deba6f4375b3aef795fe7d2551c7555ed8c42aedba66d12e79d517ddd73871b37c6cd8c679df81b4f5b7a089348c2f26b47162f17a51db058920e788812e723d4724cc3147565c2e602e1b49ff0ed98042380d989d9862099933bf6727217fe83d00a989d4d7c3a56b99450939002e75471c136e0c10e3ff13ee0e28a3b1b62911bf96bc4d85c9048be9fb27afc79542c8b2cd425a905b45b9f1bed826b13889118450e01bf6ad9b5fc5e383c3adf81be5c10f0848af29c4f9a77c3ba50f208b46947f2675340371e1115aeacf6bb7aa3b470280a5c0698299fc1f111ce0ebc0b6f2ce00f639118a96e3bfdeb7085df081cf36b42de009ae88280e4f8d14a4906f81f56bf6fd29089b27d804202e4c8958278093f8569e610a911238d98d539660edd1ce4e0365e4bb556d550c4c0ca5e2a4da19d98fd50fe789934ade6a9dfa5d3947e5b46befa5cc0ace8591b643b6625f3e59894e0f6c0bf3cd9244fe559b7aa7b1ca1038098d5953f1629c1da122bc94d62bee1ef4afe179a3cb550d4b18b38ad4588524a8125cf009a2de45136e1907e100436b567fb97422f75ad0495b64e248b5cbdcb8db60f143e4489d57721c68dac4560f184e1d805ebe6cf0f31772cb93efdb54f8b73adc63ab5ced9b26e8f5899b622c4072f39dd4fa01bef747e989ebd9a010a45f34dd88089d25fd4c22a47c7ee75eba8990c7125a5b7fb79ca1b2a6f8b75dd108d85b3d9a17df8428fa1a442447ed60e903ac9f5a171ee2220b9c189e767609a783110452e207bef11015b2cba927201883b408aa0b49175a4f52de23c812b1a809fc788b07e1b66cd5941f1b61cf0f6087581d48b23f89e9ccbd9fd9959a63abdb913b202956ef72a880a779c402372171415fa7fadc4666280aad46f2a7b0e93f57aae1cc627706f818071e867a6fd7df726d68da956a171fded;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hca9488e6e75255d350c83b51001010663fd4937bcbc8ac586964bac0430e16d9ff2fee314850a5efde81aff5855f3ca8e4fd000d5c88120105d174d6089fec20d71435dd6ab86af02dc2f14dcf44bba523a4760c26cc44a16b7e329910880de1bdc8e184f0aedd09a1b288434cd43c9a5d344a8d56bd7355cd5f46352feeeded24b73c38633d49abff6a7464240a3068dab729f9087eb03d98da248b2872b29bb8915e7b655fbbc118109d1d5030854d3af4875845d7546d3285f8d8873d0b0db9ed7d1399bd65272fe7c58872947b9303400de3faffa52c447a4e9852093021e1bbdd49d1bfc8c26e4a1b364ada99e440262cd5aed7c6acc8c5e23c169895499d8b63b101f5a692f0d4bfe3e8353779cf6964df904893376ce374792bd47b00ee539fcb19ad764e1b47c197b974db1507f7b2955bc3f10c94210d11422bf440e23d203b3144a2b0c5bbcdfccfcd21dda714b6bca18e4e07ad4b01edff37d48f1c961ef07eb515ce3f30448fe5b1643887554e580add6bf16b875fb56e4156aa2e6fac14d148f02588917c323e5ad8d5226b4772080a9089a1d39f72cd51bcc91b036bbad7ae9e888cc669ab422fa5c83888bd571b01969f9fbd5383e92d1a75caf2565d64eac285ddb9a67edbab22b057ffa009f48e20a239439a412e8c5e12669948cfcda1b7ddcf7b4684c6132420b045df28d3688ca86ffd7a31a923a1597bd0c976b204983d806df1e968f7dea63fb6908c4972e180c304a5689a32f323c6df17e71033811a0992c9dfa105b7258dada3e03ee4363d502688d440cb27b6187f924720fbce9ee2043efaf0127ef367d42873f36e3781997a33d166d5d568beceb81ea1ce72e9741f6e0de0463ec04d077b8877d6f2521c7c22e198db1ce337ce02d8a9af6b5a10b85276e7c8aed42bccb3cd2699c492b743231a74026c2dee3905482a69816562cb76eeec48c52e3a79f249b27fa5d65994a5cdf4d39def45fed4969f6c01dab63fafb0617973397127c25cdb5667722c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h79419715538bf82a442e26605c5afb7ed9bdab8c1d481cdb440cebfcefe77c39f8a772b0d41bdb841b2248e94cc5b986853ecabe22eba11b5274199a97a772f5712019b8aad7937c0873026a5e30c5f4999dcde954f9418fa10fe6ea5cc5b759f8b908e2f2c048d8a2664d585a744b1bd53e883579a17b9689e1a35f1a8389c35ad32b2922825ca0fe82d320802f71f0a7c10de6f67746b33e876cc04fb7a476caabe1cc35e855f834766facd87a971cc4e8ec0f586f32b365f381c48ef009608926ba8685457708fa7c525095b440eb6be2784e565e2a83e32b7e5abf7a82b9c85e65771e4df2b6d8e4b366d551a14bf5e5f91eff4d7075f83c9ecd0d5f57f0755906043da06d72e226eae9b6ba6af2b9426b4ff4b699f78cdf25ceb7cccfe089bbae955038f958e8eebd38ba78683e5a2067fadd77777e927c7e4373fac4d6ffd3e15f8fe142e8a41da31cb17f6ea13bc1c1acecf00771b46df6818844bab2283a7dd93071b83bca14c364b1eb6f790befa43ad0b6239e24c69ba64ba93aac664df23c96428d30e1802ac0a75d693f0bbbcd0febd0aeb9ef1c34f75c873974b49fdc7eb93d3ab198d6a298de33167719e3622f46920991e894622c81606798664909a20d38420e3abbd884768e55d32dcd7cc7c4cc09fdf0e8c5430b0f2acd87ce87b89e7fb8ca1f243ca3a65d8830d0527ad6874d885fb1c801a72a3a6dfd9a7291df03353f48ecc1a12e2d8712ae5d06f4b0f60608d080f1e9ca3f837503e6610ef5bad2ec190e684f9f0c46af2a8f525decbf55cd9c13c9e014b76df8c791ec412964cd0cbd8fa69a1ddfe5d908c4fed777966867d359250dc5f94466acf0659510ce7a411538371738a078bbc7ee5387456c453c87ca8129c4c81dfa5b55ee1a4a1098f86575146daf7d41d67e5c6521134707c6a12733c0139951edeffa0948de2868f71abcec8331e8080cb5f63b594fe5f5af01292653439f837e37fd9f714d981ba9fc6100e8a1d411fa0a72588e58916f9be0c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hee9634e38a7c5ecaafef084f7e81f3fac312266762ed5df7761f41bb64e590f6a9053c46d0c47e9e885eb67a0b99f74bc3858ad3ba268f207a4328798f3f57fd7514c61e4a59bf4f24852064c7334e242b24b20805eda7d524c8ed4c63f42797f0d1cd586deff8e51ebd30761eacbcdc5742b90080968f958689240853fd48f30e77d2c315cbb1e40b453dbab985d9fa4505cfb11a7f64d16befa399c0c42b7c55e46174148fcef3809f23a333f3a69377cc876923860362dca430798268eb1ef2f86f82a0413258d57458aa60595dd859f8a00b79f721f183ba6e4f7644560e97bb9f26bc3c446a78747de4f85ea865644f6767c7908d51c870bc4c7337f6e515bfff74613df5c52e43db7c0d22766ac5750fbb7d825df6954fb2a40eea0ebe73102305e571bad5604de5557f4209c38c5d5c031daa28015eed33e6a2d8a491a6f48c03aef9c0bf8bef3e2271abb4823c450e89ac8f2aa5d8dc023491e14f7fafc123b1ba3defad7937d5d17cccce7bebd42870addb52a5d2141acea537a21c844fd77ccc506af6f64ef86f16f22468bedf9311f746881a3f229220c8c90b5be25cd2e052af4f1845932caa24a877bc27cef63a4cf184554678090e1661f1ff2eaffa00cd7da6eedb0c76b9b65aeef8993e057b0b21fa8723d2280bf601832c060c499abeeeae63ccaf00f6de56e985cf44d8df59ef7045fcbef791f91a7b57b72d87dc373a6ac9bad78428ccb6f96567fa04cb536935381f6767028b1ac5cfb40cae8e9562e0a38b57ac0a59ca3343dcfc9e0629898d7fb0247bc4087ad67fad5cb6826f2915538515adc892ddf36a69e954429e8faeaee609315681e324417b39e8f228cc63adbc55935c06fe1c0e9c2d4f505971c306eb71410d5aa884b32cb189cf5dbff1d483db0720bedbab32e6493ab7c3ed0877848b1d1faca0e9b79513f2269990497e1ad962522306a4fd6208119dd94dc1d2f273382d97c0410a66275ba91a62652e84a295a0a340c9e8ad3bba9ba62fbe7a22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6677d7b7cdeceede71ce6225f585a734eed0f23f6f3ee1034395667eef50da70a25963688b46103038842a9ef10e72454865c5ec812587adfb38776a2b6a19bd6d101f942c86ab45196503edfad61e8f344cde3fc8f4cbde8a03f9f9be8415399a5357d7412d945b1000de2c2bac6e41d00b3c2e32e7ee602bd9a44e131f3ffd886cb44102ce1de2a98a5452b6920c56f8ea98f0e12855cc2567437f46da141324bf3aa960e2ceb42764ff7dd427f3be5c6771571f86f45d570b7afcfb024edc8fa31806e4e9290885de1662e6ef326cc1378ad023db076b8369aaf8101929c5720426e97136540c35f58204f158580ed660512c11e3ded6b59b6856c9fd07adcb9115474827d3485b784254160ede2c1dcbee4cb2b598746ad6c3d7259b0ca599110594a1ad9897d0950504fce99551b7463e55046eb2fc2192ea84689e5d110f1368b44a02159c57b74e6022a9ed7082c83408bd1ce27ff3896837a4b9e42ff141f511902cb72ace3f714dec38d956e2483da222eb4885b8e65586ae47b5abb0c291c3c9c4ae3808bb81f4dab4e1f2c9c80021dc5360e17ed708f5d32926bf48458e9917607f4c62d6ae5f565055a0fa979764d72c36a50b3b3f2046e1d8f96a869cb2396fe66a9cb9dacf94a47aa5e513eb4331e4e8d3dcab9d49eacf2271fa49de80af1e8d576bdd13aea60b7ed91a5692a81e46309e77be27dc60fa0dd578196ab7886326a716f1e18dd516528ce57f87e63b8105fd385629dc4ef9ee88934f5d50ff95a5d0cfffbd21a7eac9137bd444066d3d1ed20db7c14bc893a7b482e4c40590a5a0d9159021383508fd58ee042f856c4a3990495c3ea3569edb675d7b382e70fdcb535194a3cc3616fb95ae16f2d1ed79501860b6384c9dfbf0bd932cc9448d0ff44fe48a4c8a90b53067953bf9bed8286d64886d37db0db2a3605c78e9a5572496290565430f7d0b11401b2338537b14794dcf94b31892628334b698a2c74ff1513a2db66db41ce73e8279e6d41d6c366f2ea7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcbcfad4cab565fbc140cc83575dd342b3612b41db9913873266836525cc11632327b62cffc98b5c956f7cae18f3b0af3297852a6567ee00e1ba07a66d1a6229ed328171bc9abc5115bb231e50aa518de53c9d1c3cf72e61602c6d6c18facd0843fc26a37c570ad30068dbec03f0dc0b7c8b4ac24ea93506e5fb7b0717620df090eb21fb67e929e8bc486a6ef34f03188a1fff7cfe12ed36a99ec244a569c9ba003a45db3aec5c49de68f159dff54aecf5a1ac9f74275896ae7bdc5c51e6b1174a8bdb6171d856734238ac4d8c61298591b03f1718474b88dcda4985b0f8b8e1703a7cb844c1cf8245d660af1f6de5aaa96395b4c409d998e463f209ac09304cbb4574df3ae5b75b900d923ecd5b71c706b5d92531447491700af688b4b99efdce63fa5bb17fa78202128ab30bf13a3f27ad8166e001d3c5133662c99352efbe8e6d617be8493ef37e0315d16388992839d2929bc10d1865822969e1c087566c54de1da0d1f54fb025ae0e2553b7dd8cc75d030d599854969747367702ce18544e13ab788b50c15d8f54c29b96b5325df4a4db07f41a9404c759e829fbf73e46ee4a50a8452d047b0d03297b32552b5c094024b74cc14aa203cffcd571418fa184a3ab0907cb44065b22c72dc3a60e37329fcd6584b7b18502851d732323dccc2e92382d245ee073f0fb8421736a6193a6129783048d03501246b2c9cd82c5f804263ab9694e69ff3f2957e034eb7c89a79a1898836c6e908b3a352b45787ef8d584ebdfe3166dc9b484b12997383cee1cc10f1bfaa83aaa0ff55108446954dd43756740a4cc25b8b1f16f77867a030815cce23008cdd5168d23c5e0ee1ebb2615abecf6f648321f410a643a1065dbcacac36341b025f31c23c3e1cc772abea8f7d53b5d02d30292419a9f4872a46afc3c44b935678b53979b38499edc160caacf82562801242bce0a29fb61ecd9d907cfdd3d808402a43994578552fcb9f40e30d29401108514093455fd73213870c573bccfd3b420f5304bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd060f1673c7fca93055ba529f08e84d7d7c0f94b04f71a3fd6245f9214827b91e7d276061f6b60b0c0d93b135c8cb43ad2eaa0462c56c8a37f081f6dc7a58116e5cf4c3fbb7a4d86fa97a7952965ea2e66ef284ad963ca3922fc288a1cce586ed3f853371bb84674ce4a6b763a8bb2864ee6bea025cb4d8d37e4f0bfada51254663a5c9263a7076be85ddfa8e19f4384e63e5e5eb490b648c713d596e5062242a27af185ff091dbf6984da685d2d68705ded18fd2b9ff0b06a923dd6e6c7f1c791fb3a8154e9cf023945ed80e36e39b9c10207145e19fa41f37de9edf6792eb008590df4e8bd3cf9cc9cc633e0f2b3b94e2582bf4c590dd33ef50a1acdc1d0447e08750b07d569ea3df9e6da8c8f6dc6978c76077d263280f2de38fd0a216297427f5551984b728f63a67ea70d5d9310c7483b6e8268c21ff968dc1f52277a7104ac71a106d470f84f9d099dfc81596b1a71e8a0d198d0960cbc7da52fdc43195a9a70f80f20f321146760b5f53cc5efad6d85a4d668185af7d0c76e2fea1167951f89086b57b841d8968dfd83e883d908c10e9bd330e4f757e89dcc3e826cf4fe92f5cd533114b48ab2a9704b702f484d0f8eb1859bbdb722f73615a7c3055203d664ca79b94f9c89dc5d53ae79657335c3cb6f584106846a54dfb89ef257452bbcf67aeab3d4fc06bc786be2bbdb611c13bdb3a8b4c5f7b6b6bb11dec1e260c5bab89965a30cf14378741b3c6fa3decc5d1f5e9a491c31693fd498b1c0196fbe920f0af6986407311b830bb07ee6a43d20ccd29eeab37bdb30b5e2e5c67580f24c2d1073b861863d507d88f8071309f4066f3d8fe5e902813501a452ee0f5d7c78e43dd5ee740d9a5abe555a47f9dcbc9008adccc7c02aebf9a03c3839072c885933fa70e40d72988f225a26917b9ffe8ee3b59dd9a765d4b5ead33678c9b2c043fa87db26493fce8ae9c1b6145ca2c060782e40d021e7931a3ab6830cec599a87ebb0b2584eb9d36252a179cdc35ff1d5c832d4b8a549a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h306b3c02d33bc47a4d14cd924993bdabef4656af390494ce7fc98f8cda3d4e066328f41a1a0a72cd073bd1b6988dbf33463d10726c535ad383e1c25c55ab01783709948c29c90999306ea1321f6565a51b5749782c99a6160e8a3887c6bd5dcc180c074aa80b437de68463e73fa814a187cac69b22ee5847ca16b685fd90627b1be680b56e81f62ee4530bc60ecb2778b27382543079059523bc9b25f44fc64d2aa9eaf1ccbb043f02bedcff3c8955043e62a5e61247dd1466eb87579804004859a060c3770e7cb9c64c3626b376154da05251dd6a09e385abddf24710c8adb00968cd263953422689fc039f68adfcee2a687b77d4904e20cadcc59141ddeb6fa678b579b7750b00f062ee374f574e32c3083719d07285771e28a48a15036c1497074dabade37533a3871f4539e95fe7270436fd432e1663ce65d08ced44941d1030fa6088535e7a7012dfae86f145ef8633028dbc3d3e5e6aeafe918287ed9453bdc742827a17d9db28ea8dd7fc971964a1da901912398b75c4c730fc7eff1acce61a0faa6cb28f2debd80c1102eac931cdd15d473e2ce27ea9783a0cd8b759ebd8952c78e3c23aab08c3ced2d98947a152ffa2ac7493dde48b8cc5b931f212d7f932a1240d6b835e0aaf10684c4a8448463a94ec28efb991e5ab259b0af40cc69e190d8761b2e43e98ea8b1e1c6ef96a0acf949a6b073ae1eeb4ade0df7490c618eabc482ce9c6ece68b85286e4a2e5bf7306b7e1eb2247871f46b71ed8e0925c1567a64885c0d2f5fa54937b4f6b1e99314667a5b312002739d2c97aa2d2d5d20be5846d8ea8277e93770beeb691093f0bda41ce13d78aa01162705cd36d64a431ceb9f57fd667b374e9daec5a2ec02341ebc6f56d58eaa3021ca852b2f00d342e9a0ce45bbdf5ea4437654f88def0b4aec04d89c628c7b59ee0b4bc930add11cab516061ff6d478632ae302e496c91aaa4e79b0545dfd51f635e5e8c75655281321386580b54869faeebd1bde1cf51a7d43bff3c2472d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2e6abeaea88fe5f6d50915be62ec73e24f22cd31777203e53b083f55d41a0f023c4b275c7f19f3c34dcb58773b1f182dad34fc5f07cdb8c357658393ca98a079139561e3bd11c6d3036810e2e8f4ea0367e1f8331c43f67c9de75fc61996cda227df3ce3a556e2c9245c7ca2d590eadbcc1b08856f91dd654f09932403fd3561423249f69b699d8de8360bea494c467737c4e483b0ae5c83fc2840ad97cb94f4b056626807ee0f7c0dbe3f84f25493a8a07f05a727228ff0a60340ffc44554e00ff45ed0ff159d8f606ef3cec14e05380ff42ea43fb78d80ddc2b20ae391612b7dc63bc76a251e3b3018dff54e94ddb45ed2cbdd9ca2be1a3485315aa99b2d9a12ad4f144130aacfaf3a760ca5cfa25278206370a4b711ce8b81668b2cbd4e7ebc7f18530b937bea297966003b48ba64156f94c5fb7ebda52a2f0a31723ea79a0843255a233a05b0d165dea3674b6918c12f5871e49e1d4157b29211c8de87ada63344ff63e15474e0da906bd6b7b553d4019eaed7c80db070b8202883062c086b633aa3295e23debdd89b732be2c040ac5bdd439c328724292a74c12c56abcbb40adcd0b3520576aecf189f43bebfd1ef22e6c50a727f35f572cb38dd9a08f10ebc10072cbdc8916b1d5f94e83c23c27ec0ace4cbeff7d4f6e8d782163f2f75c7249885e5a2b2d961804ef5e76e37e16e6aa39f1934d54cb47c527a043b850521212ac2aa824b41eae8e429be94e57e7bf1158546267b4ac2e75431554f304c5cd3310930575e68b16da1e6a90fe457b2df68413ea6d53dcb12a1ccf72841711cae7c6236f1d0087f74cf94e5c490480ff6e57041679b6884228d07c8996884e861248dd7519943d111f142ab23993a573bd3647e9ff91bd04e0866d6669cdb5bd0374f58a80c31bcf08f1843682e9dcd433fe3886c9fa0805603e3ab07efb80002ecb18ae2f265f3058ae6f486a53f436d6848a5be4fa4e3891325e88b1e2744c53a0f65acd0209e47e07278c59844a5519b6eb697be7487;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h775d5ba99262cb42da3d0aefa638c66d56e58b2098d3e3d42426d52b6da1f85d219a3ea37a2443e254584dab92913de9d65581a1c2d9379bb6d45fa02969ccca0177dfab81a48ea3ac87bfd4080adfb80f4ddf643a26b3a0b5963adc44fe7aab898a37174831e556c7097cf7eee79de36b88e7799ccd36f0fcc2883ed32fd88003891810c2e8cebed0ffacf26e34159952afc65a15df192af437d8004c240d19ccb4ebd7c3c46577de8472076897877b9afa7d77b7fbe1b43558e0f9c39beedd5db485cdffd3c2d7c35696fa430e27f6e08c814af66161201760b8f76cba28d1cbcdeaf92e3bd6b2e0fd02b0fd3cc93a8a00a018d4f0cd7470ec117f232adb5211432d740f3a89162983c6db4a016e78f12a10b3265b2b5c541ddb4d1809bb4e3ba230555a4150d310e7c00458d89d99cc6b6e76d9303d9919761b1597496f514de264c7aefa59274fdfa6ca5b31f0ea2a1f2613166be31a6252f75e8d41f2578c6b31fdf1bfcb8834dcc095b47c500a7ad54f2104cdd73bf4e534fd3dfb24318cd48887310c74d49bb16ecda4290f1ee6586ff83cc8817e51343c878cbcc79a6ef391f70f3dbb7b7846727dd3d5be0718fc17fff73250fba3f7652e6bd7cfd97036c8a54019abe931951bf928f580c4a9538b0f3ef90616b6b8709440181eb6cb19358842ce9ea6207ea61af8243c601cf27a31b12e0010f4ee125bc078a3d80667ea08e761b2dbb3dd0f58ecfbeaf7538f7a26a639dc0b10bcd61b8c1cecad0099681f9f63d4769179c7e9396a6eadc7eae9a27b883b1222d5abfbd739c822936680b3573624111b9164c4a85ed8d74151264e6ec803e18a33c62a42cab6bc57f74bdad34c8fb282247e78d0bd892de6d813627d0bc2031878938f9818ab463d56b7472ebf2a6e9c7c6535e6cf6a40afbf0a1f62672854711eab8cfe0b34c1ce9e708c29a56d6f838fbfc2346be95e3ba92a40f25fed28baae3d57cbe35ba7bd97a2fd60fff9510c95ab12969207cff93a7ad2a14223aaf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2cbeb5c9db76124343a66691b802084f0077cd34b95d9d988daf8528be8d17350e3f6e34de65f6dd581a1d7b6568ee88ed77ea8a0cb03b91ba7211807d80d249334d005c33ef1cc6314bfff135cfc820abf9652c72feb81f0652cffdcbec3cd2e2175a6913fb3423df94158146075450483a0ea737f53591b674dd0654ab1dbb8cf5fce9c74b25ae26db216bc2269f39cd0ad33351592b8e643ab594a0daaaf5ed3ba2068c20fc5543592e3ffbe62aae68564bc517837ba8c6ce6c64a0edc7bbc09d24f98b919317bbc9719ab80e2a809202275efa3436baee83957c99674ce65f73f8df23b121224fe646289b7f702a39796446368be85ff92fd437523e390a5e9249c4114e58bd4195a8b35805259968d71e5403c4e32f5e853fa432b36b7a4e9053103298a954bcbb7f0e3cb7e9c361fcc02d917c37787d04d1f31a8f8db047326c1a4f6fa834b28404ef6589080507f56a74fe843e1850859b559d4622121cfe815ee5f759cbdff37961a7ef68779320ca07621aa79f781f3cc8f0ef20f414cbb3f64e95c53ef83b9d27c1d27393e42bd2e28d0111ea291b36c5508583257df4312a6f425f7fa1f02856b8a9a24e4195320eb1a1499986facfc391f31a02cae93c638ad0f4193e5e942359baba86526b16da9e766f3aed3e21c3da9bacbf97bc761b8f5958708168d47121221ab082bd4e8cc6cf48ffabb7da3e6c199f357cba524fb6a5a40d9a3a52259996939b1fbf09a67697fd8136233f742dc6be2af2639295ebb12d58e42d16e0b4a36d71a49b883f1252edad82ca9abfef641ce0b6b06fda52fb076e08755495022f3b80bc7b41eec05d4b7ad78601eaf0b1b69fc2488b34b17268819cb395732f51be95cd1fa607188315631c237bfd22b489665b9e3dbdcc7dbaf32065bb56f8e21a020943938a54e7dec9ad7f28adda29cabfae58114089b28f172ad4aa569933dc86a4662f172476e9f378f7886ac78fe7a1c80368da5d07e17bb6ec0d042d4e999538bd51b4a47f101742;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha90dc2e030e851ff2e7f85f7f166d3f350e3fb801c680c8268ff23b97da9ef08c2a08c5d1994277882b1fc47863c5835562fbbd7c5396446ed7bec2ab0b888a9bb5f4781f9f91f9cc79efd1118469796bf55c93b5e3d72d28fd9f561adf1d14acd2efe7be3ade979ede6db6a44e04c305275f229cd82fbfcf2ebe791621eb1c16a1d071e08ce2dd9379fd4bf57d9e67e3d899a0748f79d92076ee3f51eb4130ae505a22d1e80357424f5bc26661b96f1fa0ad9491c44adeee70037c702622b498e45b4395fbd448b8a22256dbec0d066962887f1f1e365dc823fac4e1a1e915382802bc28200073e5d1bb5329ac009781f4ac170357060b728c4f53e873308e1eb1363c19a961aa8a1bd456c03defd7e2e942dbd4d2fc3edcf87af1dfa6ce7d5ee448a5f4cad27bc452d05d721934cbc128c01b3be6ad0d501c5fc8ebfd62c8dc46f41a28f8d0acef38e98c4bd7c449def917a10959d6d1bc258c8c21e9c226e93792f1917380ce3c5d412f38ff2e75d33550e40f79a3c7cc1d7888d0b3946d42245ae2cd48e355fd048e186f88d89aa26e981f2eadec72ef6dcde787924fcdf2836816523d54a8e17e31a800e24be43a92586bf97ffd91ad68a480918bbd5c4721da4cda365a5a3f8848f89262b76004b6631cf820faf5e4ded26329c0ec3b7fde525db1ef13cae3b6784ae5f4b5b01adf05ffa7f113dbd68ec4d6b7fef5732f9d4df072f9a0c7eacc8c494536f260158819bb2a988251621b9dc979e5a94a76918efed8f324fd1cfc62c72e2c232a9401fc3d7f089ff9253028fc5268b18a8a90af0638c3d60804af5dc9280fd90c32b258e4e654ddb159b839fa53fcf4a0cda21e90a0c59c86f78093eb60aa59f5c9e17550147bacd16c4437de745e1b9bdbbe0c1ecdfb6e01013e6029e3bf0d07c163a0028090b1eb1bfaa998a89d6c519f9816b3c55f54b9b26e0aeb4edacc8ce71ab2a8940f748bbd1185316fcb9f3c7cceac1231fcabcecb50edc95def531c89bfe3dc68d1206cf5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h46ac193d5407070d8080e8336c69aca4d7343200e0370cdc83b02677546d95db22ce2963213b6f5d2b8a25fbe33b59339f831264f12f348412ae630b44f685aef8e5e45c49b34144cded166757fc429fd8af92e4f90b8d9d2aa0cb74f8f335b8d81f3797d10dc1bfba687fbb3bba442c30af8c4103d2e4d1b201d2fa2cdcbc55f5ff73b6bbdf1e376f01552262609d0d82fcdc3079029b2658aca264d852f3354a969ae35a12a7514e893077c46a47487883de004be26211a987ddd9b534a99f42cb7b17e0b805fc041a3d7fa5ee536ed27db74f9f96b171f5858718f94e3f9472b6ac44aef5d722e6f045da85d39df59de5fcd70d198ac5c9f628a2053659f4876d0c51447dbf3e797eb244de9502aa52925bd8b885227e08dc1054655c45a5a3387b7cb289433386e62d191f9fd5643aa584a7c7952ea7285b2d36fcc7042db982f739b072a55896fe3a73da04e9fdbaf4e788dfbe4eae404fa848697d97b71a56a9452edf54ca338b8b7a5391182c6ee95f8cebc537c3ffad1dc228184097119f628ac1f6f029309aecb8e01db19fab3daaf9c12f276983e133fb38bc3b7fe6c65c75cf415d253c0cb6e244e1b122a70d98c08c0869403b36c90cc30104e98328f746dc30f6c437bd091db674e73d809370bf5c8072020dd190377d74fcc39d29175b09031194240d5bfc0db29052ba066ebc6461d6adf35bb50be588ce64435d4c90cc352641ac61b4b849d62cd05ec30146a4bc0e3abb7bd6dd0af2042a87ccf0067866ce36fe77475d101868fa563c965d13b46428efb73d2bcdf44d204292a0bf45c5cb45911dc48d582d63b337f12c668b9384a838122dceccdc86bd708894531c9884cee62e1ec15e49cbc650869f0ee25315439ceed10b8d16b1e8d9b858ab8c0c4e853087e748ac8ffca6dc95aa0de2a9d30d560c594fc501e6c210acc490bd9fd08b22b68ecf0e6406d7718bd3da7ef954b049b0c92a6f20ed84051cf03677c6cb02da1e370e0267a1bdad0415c5426025a0a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h62a4e5e4ffb939ca99fc33fb7d85a12a4e65553062df936f2ebff60b2c140904b4a2dac106772fef9dea0b7117408b6574ae81bfdf1246d7b4509792736dbba32505a78fffd5937a0c43988e60ae0459105c138f9eb6bf115177fb977546c0fd8de87928a6677b0393a32c8f8873c597272b20c725995977b758ea470f91938d798e325d6ff23a3ba063a27981c5bc633e331f53baa94283eca17653c104802867a8bc17f8d67243c0bf073f44bca065284c5da30ae5c4b7b13803374f72810be53e212f347ebcbdfb4e12417a193d22da9546d3dfd8130a44f3e1158d10555b56dd2c367627b38cb72fc8d7b7561189bbb56bc902c5575ed170d640b7b0fee0574a20e8d22c53df33d1c19d48fc389656bf9e9581d9992b932580faa412a6e56d9ffa7d7bd845d9936eb8782d6b48cba8f8f3eddf17606280292ee37b32a98aa8d7e3d3ed6ed420d0ed9f1d1a51824ac4fb92feda9fbcdd17aae36214ace45812120dd02177877cc925fe9098b0e0a36eeefe482711b6a8be8452ce0f6e4839f066c242c1d09c037ca68724fcdc556d4b9183ba6d66c35505b0299d615aacdd83059c64995d7f9e12aaa40a640023903c27043def16ab03d6e47b182dfcdd4a0ca0f14038dfb1a4907d4d901fd5b1f93f0e9ce89111fd2bd772bd3ea8a4986a74ae007fe3bef33ee5add3d47dd87ff3037ff92478401ee7a82147e987773952db132b81acd5be1aa6e832d14c6e343f0f356ac4eedad522fffd7ca9905244877cc91d4ec787b5a09e41e9abfdf361ffa0ef3093da95778b11289df23d46a69207798306bee47cab5179062c26faeda7c7b90cb6e29d3984cc053948b0f99a9a950a36ac017ac716b1e9937df15c35c678b0e797e81e256ecf3fb344d948fd04285fcbcfad0228c4a3de0242084abc048499d3bf6c58a5a43cbd8781e38a868b5ce7fd7348a4814205cc987ee8c28e3e79539addfbb23f91e53b8d040c0322627fb13d67ff5c5a6d1b0ba1b3ba13174204cb25e8aadfcb6a21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h91787a8d7a2068dafa13c90d2bb6f61062465acb8310d9cb85b75a030ecab9f9ea55f121f62e6c4b244423e79195cde03c0ce6b45b31cb3c6dbbda241d285c914bdeb2b071c4cc8ef24163de495e2c320d4d71787b008150b7f06e13756a2d38bd55f6557b8ee17ea6550a22433981c78e1a462a338d56821c021502cecec11b6199e499fe03d4636e16af5f298bd2ab2fc22276912f6dc43dae075819c1c16295b36e19a7b26f23e14e82b18bcdd0870ca4a67968635f92993e9e87e24153cb3899feb6f149cf4bdd4a52d3f2c8ada51a2062371614bcffe2a8f36f24c6106e0d981626f0bb69be2ee925538592b67d917a707fd6b8b35bce62c375ee76bb3634028db830cd2108d217bd1995181c7763c62ffa0dd64eda182abe2c327867d1435635f48039566e1a97a365ecb54b217fa9cc1db521dc46aad9fd80849cc19e29004085bd366d1c882d914c7b80971b824cd1091fd96f8e383b94c35b192e74dcfba7e8405a7aff0cb954ab9e33679a886bb74af3b9d529226b10dbcda5f6f17605b4de982573a571bc4f33056b7afab1b81a86acbf94f03a2c0dfc73765a3a2ea45ac2c3c7fc3d5678c23e86e5d978e32e8b328b376b2b40861d371da28990e997b32640f868c411116e660989ba1ff8c7315b6fcbcf89a72b4ee72890b0ddb57e24190753ab46eea95d91fefc1575586364c0d13f832bc35a6d19ba9639d56b727a9b33c7da3c9f84526b280015445fa51cb6ca4530a024d167cebf4747bc942ef341fe98184dc3aa7733e1995496d3efb3522616dc66143493ac1d1c7c9e61018abaaa38abb66f55ddb89b04ea6b049aefe1eb40107997b577d2c23dff422b60d5066fb49db8d5ee8bb6d856861b9998ec25117f4fb25db713e4916a04e9c6e243aa5a9cd465c7780d55627eafa01c89ec50b7c290c7d9c1dde870c453c4539ad1788b09b59380bbb1e3c9998cefeb852ab1a603645aad33c575c558c732d760283c096bd64cd92a925799085725940505e4b3350b63ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha1ad2764ef690f8e4cc548522bb8cd43ec2150a8c6a89707d6dc37302b89c8fa08c411b6b58a5a2cd47cfe5c2594c15d15874ad6c2a82582d00613fb8a8d49d77d589589b936dd68985921dcb2ddfee42d036fecbfa9ceba11d17aa141e060ff58fbd682ab2cbe23f02c8e73b95dd248a1e670b101a006f28c78dadfe8f9e8826d5aad8de351e85ba89280a2261655e9fa4a08d73fb6bf06495c3b4a15a8131cb099270992b98a3f801d4a2031b0f2c085a12ccbad47e3a4eab93775b0a5625aa1a8134c8a5097f550affa93ff7c15f0846b2b9449e89ed06d96f928d771f07c1207770dd545c8e482f87f824eeb76114c38d5aa40be367b61c955704e74f6af444247564b04b5790db2c4681907edfd5934bcb00e84681c85ba9c9a1636a92aaea2e969802bf091950f599e1faf8581ddcc270b75cfddb900b7b8a59492315d8d238fff9daa0f6b79fb1c5619c588ec5b8803ca74a1e6f19c57e8dbf019682f12763ebb48afa5d2c3f476f94fbe06377240595032e822476078389b5b00f66bc35e3e9a1942d07593d0cd50ced40863f62443f4ab59edc577624d4fe9e1eba0578026ce136d68603da83647417b6c596372da3041a4265c9686a5f0cfc504510c8eb45402d5e6dd2c0ab3a6c4236291c2e5007faf6fb2b8a36e8c9e1bc4aebc2245e33df356fd55cacf0e31f69ac70af2accbdaa36691929dcd18187f18b30c26d37f27cd48bda4a39260dbb7010d27afe945ade0d8d9176553ec85d89d88788f7e33800d4802ca826987768b3ce27aa0cc2d2de5427304f2607725debd6c4afa1c9151de262d229c1d8426512ffc5f15924eb034afff53f69e5f4219280d3bbc3188852080d4e8bcf7af14c4fa4ec7ef63649bcd6243eb871b0869e2f713c996a28aacf28847832935490c19d8c86fa3e5b5d42409afeff43d9e02bc3e41d80cbb03e86de398a8e2472afc1933b63d1ee4344108071fc7e40a35f117b1fecdb6b208ec1540eb78efb26a754b36a1bb1b876a0447f1e7254c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2727f1435c21da1c8543c3d47bf606731eea51c79b943b2a7bc572469be824c70d6e8ad22933e5c0e2a49f81a5ed425ba4ce85bee825bc2a0a8589ae799138e3b65f3fd45ebfe8f5e74b95d15c85e9f9804dbd95a56463b131dfaf2994855f3be5bf5fcd7ad1c8cefb058059142a0fd4841b97709aec5cae854793bc16e6e38c018c8cbc9541bae9e22200d4d7b7c1ce4c5fa9a7b53ec7e0c3ff1550d2edcd0e08fd49e326ed3fe58693bd6277c62abcfcc4b413b4972473f76463b493df18c66e47cf48b95baa87d2b8703154e8572831bc993d4e6bef6e051f582fd206948aa9e45b0e149bb44316314ca21847a7a1cdadacd34964350f6805a5eb2dd5c48dbc3553f9bd8119f9d8be8bbedb1e09200c66046cb42a3d83476bb0763150c2e3b829facb694794ab188f4ff890a4edebc5a5e17ac378169f9c4e85cfcb225d109dcd310df863201d332c5b5d683c062eaeb43345eb2e28a2bab99438a48642daf3fbb0cf0c375cc7cc12d9d0596ba32573241e96c28be55fc9ac065e9626e6f3a4eba06fe24ac97c0f9a38f94b192894e3e730f45f6f58a0f7b48b46ea368feb260c13c7b6ac074e0e332c433276affc3a2555d5c1a9165dc2e544b58d911695e58b4987cfa97f17445174e68f012e42c3876670ef42c880bf1282010018241c11be58afbe09f4266160d1cf423b24699807b3d7621d07758f7224d4021c7c96f8c1aa9901a70e180edabdddf5c1a36e84ba49042fd418686ad4e6d61a9de16e00f5033daf6eb91e1a1310015334c67b059bdf2a7211d843d1b44878e6bb84512d449cb2cdb7378ae99232402ae3e5f9328cb12eb93ff9350d83b331b608c9f95ae2ce5d4dadc4102c5be9baf652b23f05c0d476e69908405f6c8101faa49eeeb19a07626a3f83713d97f7ddf38aef6b8aa48b91c2431ac44386df957775fe6385020d451cb9a9589d1a069382eac888a74244b7b7979d435cdc1432770ee3862775fa3617737493e1f3e68f8615483d581942358b2c4e5344;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h19ba3a6cb262e497de84d1496c92a43535ee2a125695fb6ed1b5d3cd921cce9349808dac801f03752787ebabc3950524e0362f623592d024ec8a6516b73b355be45c6938fa1b7d9a96572988af78b0939edf5aa2251f519bd0dab7bd22a2670ebd6415722672397b3f6d2d7f2b014c54dac8e5b056c496d2b955cdbce8ea4ac9422d67725c6b5cb3afa0f80ab006fcc38ce3378f96bedc4aa49a52ed7eaeba380b2911f9b65421d58abbe6d36cbd02049d2b7697fa5a60dfc4320c3bb2c6861f40d6e8f775637ffdf2f3e906ac1f1c960f08e71aca76bdc922a2ae6ce09d2ceb77973ee314e18aa93c7231d842734444d280e00865174b350991155a00dbea277d973e0702902caa0cbb6fbaacd820d46a71f36d8c9215260b2b5f5d92b74ee56e02680d081b8478e097151ad60e790d9a139bf9a4a0feb737aaaa00fff3fd15debb6c21daba6d04e583b8b5fe2cf74a7134c1baf094d72267b80636b853ef66c5f5fa1c77f13315eaedfe96f19e758784c77a6fff87b20c6acdd6f85b92df386af03199b54d1755d0fc348da4c138657754d9093e5f6e76561c0134acd2a0b9a20cc8abd3a5fdbe608bb935df7acf3b447a80302f5db4e263150097c2171a6393edcd9e8fc3fc222bb2b32906694c17d6d69d01f1a98fdb260d10ecebaedbd2c3997fdea414943b613f54ae70529b43920fc895bae0fce406a929641e8e16486d39d841309699ac2fad8cabe995ab8fba136dc95b5f70d34f4ec9742b8ce903fd8e1c6af61d711e05771e289f5ab4cca0649b29c34a98da2f1aaae62c3fcad2ff86bb5131cf57cadb7ef2b4a8a51e17017a4fcd5be359cfeb9b6ec7fb818f197a48ec11e5fd0266cf5f33cfa6eab2c14e1ec36d2aec5dba75c6efdd0b121b84bc1f551f23fd28fbde515f044044013c7541efa5272f7c70cc78529b7b824849b0a8d05db4d43f3199e33ee2695f765d6a2c9dfb7a4230b337d2367e03a229107f9394653c5056701ae35e2ba99ed856ec444d60eafca206cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5d4492cfc03b5eb7fefcfc8ad22da9243cbadac8235b80dd2d74bfdd6abb719a17e06da583421cfdbef1a19aa4ab9880cb07a26bbd8fcee69d89d650ab1b344acae72deb58bfeb1a462ecb0631948af6329264afd4631c09c876c979c92a1237c4a8188492eb21d6199a4486398cb6d857fdde2c6dd211089d50fb6fc56a49cc6b88fd0a67da964321f90b131f7a80cd7fcc97cf5f940ea7fb0fc796823f84127e7c168dce81e2baa70b8381bf165f54ed3732cbab415d681e05f03a9205498471d8118fd98d0efce5b284db13b98ea6c3a949503a714b21b224a7bc74c26d5e4e628f9824ccc8b0d97ba1a8b906e2232e450099e911d5e112bbda2f6f45199b5bef4533ab9ce9653e8b96f096a4b6bdd9ef58f0359f83b8819efa5ca1d4d597024beaa181f3c56f759d377501b604b1653a93b8af0f89173482a9f3c99e0dafec3b1d1a2728551a8cd0a121b6a9201682e5f0d49111ba9d26216882554348da63d79ca1b140cfed94792186951864d3941888df62f24dd57b24888cf637b7c9951380ac4657bac535f51339b5c82e1517c0b266c65315b11462b8c739a979ec0098d9e983fff7c205945e24422888c32f24a38e94a54b13b90f83e71584161c59db7be46ea1563ad57bd190e6933cc1460c60003542d903a159b63518dbc2fa579788cb4c587044425bd31c7a6dda1c5f1b7b88f4242fd721066e0e512bac2a9b054f281415c3794f20259277c0977b358586d529153f5cf518860c236a230254570b97513a3992f1b1dd310cde16ac064bd8c2d4d8fcb013c0350341bd8b5c5cafe4a07dd35d9068258ed930ff698fd68683cb3f4a6edb83506aed8f1d49e4758ecbb9fdf168363f88da12cddf1c6d59530f4a98f97452cc4fb53ac5927aa591395231013a3d783286a02466fe4a0289e879268cfa2b9e8c887d1536775bc02ca317e442d87213ff8e3b53a17322c2bce07e906dfe6e4228ac1d967b598772a018c4cedbf9450d56f96888eb629bf369be9e4ec1841bd656;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h310ee3915d562cb1343505052209c828008d39b83f67dcba067bf5cd4f3f73ce2ceb9474ef53e2440dcdf298a4d557fe053b5413f9775c7e0bac4e8244588cea726b3630bc4d3201fe172ebdc3b33f392ea551ef8de21eea20a8a4e4d4580239ecd4aa9a5b08420d52494fc3eff4c392b06449775006880d2da5128e8d287060ae1c4bcebaf9c2543d91526e88aae91c3dd5a9f3ecdc2f0ca805a9a76c7e33158f1c6ee804337ce07896b27fe98b1b03605d07e7c4c9aba32a0405070eeb2354ad6bc2034af95249780d32b8d3c785c73e094f7e0371b90e9c6a4437bcff7452c7ebbfcc88c5667aca393a4fa6e0a6e1c7c1ef277857d884d295e53faa0b1cc84bda0e678df3a41636f6f7e1cdddfbb66e6786fa4648fd12cf7790e431f6c5f55c8b6218a6e0ad37f5c11ad9547434ba94d181031b3298658d7d04b15cb378daad6879a7774bcc674a97e6111da7d5b97022926dc1f22b76adf6fc9170499d835fefc663c5220a6c8344b5df729449e8d90db9dd2924fc4fd1f9d415c9f63ced9f88caad263b0b65bbec904d925d7675643149f866df9ebb2867085631b83a52bb57e46b658c9664eb8e7e659ec6c48461dfc2f70cf2d61b72e4cf898d5b2583ed1649dc498a000b7ea3fe95df8a5004c8de4f6e7d535b2bc66ab0be032d7c56fca752375f0532af6c525bbdbd1e14acffe1039b69679a5f52977e775f2fc4f57005badd0f87f6500be01bbe17f8fc9dd2402b57a80ec3e63cd9ef8d201db0fcabf728079618abc840837941ffb52c19146270981cf42c456e9e8467523dc566c89544c76389b5560f5ec3a2d7f204eb98f201594c6e19de92283b49302a156e86928380331c47035128bfec3e568db053d9cad812639ef827a428b8aa8bf6c42c49f4b87fb81e37957903ba91b876b31b5b18cec985f8014b0a263c358cca6897c27fe352151c6669a97f1d7593003634aad3b8392ae018dc7a353e65a080a71e1b38ced576d9ad24ce204913722e31b481bddb1e4d0fe88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4340e1c0b8d343da662243e2f5b1c19d7bf066bfb50881f95ce215fc7fe856fcd1221c09f753dcbfaac677fcfdc18b4ca024fd2e3113702ee911384baaaf68a670797051bed9a1c2d65de92c7ede3f8891302513bbc496f8be9f54d56e75de4f896dd6f18e64352068c4c28ed75e165bab23d5e2f73511466f04e4c7b5a33c29f14d70bff69e598f77966a62341b9bad876b7224cc9fb16cc8457867622c2e8d5155a857e62dd56a167e3e026f7eba7bb56fbddfbefc7b8766db15518057893373acf809d914a8cfce485788c52530202861b556a629b4518c1499185f0379b993bb83d93a590ee89d8a9cde6d719aaaad5300c6e90c36bb08e5fbf17a48f452f0dbc794551cb46e952f2cd78169631afec4da74d93db05234ef2a5daa0b3334f9dced7245f4de1010193e4b3ebb29f2ef4c4d6de323bc57a8e6de245be735b2b6a9f78c2a41cf75ede40711922f417ab8aa106404708f778a9fa099d0ebcde1a16526ec3fe801a18a7459996902835fadc086d9bea462ed11aec19ccac4fc7db4d5734103c7bb111d353368f84c063901a770bfcdc2a6dd4153dc93a643b92187efba94daf806624ff30179de7876ece3eca9ee6c30b3e6ad17d9fcc5cfbbd4630bba65ca4d03f9773906b41d366ae45a65c7174c6bd89a62ccad9dd7b509e201215f634274ebadb169c5addc7de4fa48b3d6477fe76edc11dec3c670fd84d38720665bf1f5bfa7ceb1e3ed1ae71585ef4e880897f3d77ee9bd344a671845aa09b723070e489d8c7183b91a3c06dcc23ea862d4c2aa4b4d816a43ee32ed7b01042179cfa4332ca8e837aa680b151eb5ac8363eb7581e12c1e5c15ffdb5934eccb102fa591caaea5396c68b1e6ece06da65d28eebbcfc30764beb10a14b3140b928fb4475ece99ff8727c02e1522f4f5fdb5f7a821b7b7bd424927c935994b2933680f9e41954a672b3728d3a49ce32554a2309b97cc6a8ebe3ae734b758de6fa90dcc064c2b8d439982f1060e92cd24b2d0e1ed532e8de3eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he357ea691813b20d6257d3a6291d0eddc502d7cdef643657767dc91bf349c70024e370bb80f3ac35ba05794be6921165f2dca028780a0ca51ba1903a97b05de91dcd7f8fb6226d2d0c591770485bde5997160bb2a4e3915aa62bce148d624a6884b4068d5e054eb7a48700dbc2ff324fe7a5709882392bb4c6bf353e1d8a971f1684c6955a5d6000992c69ecf28e50410b8cbaac5d3213a1aaddb8ffc4ffcb20a29faee1e4d317fd2302c1c26b417f4d24bf9a75261006b3605155b5eb3bdc2f9d3666d7880bc7a4ca15ccc119ed5fd810fa560125dff1d321a2ed65be274490339a50724a8585f25e98d9a80a9033a849556a377f3f2469364b63a6727f5ad704d110274a650719bdf0b1da76a17548e3b7c174e88c87e3f63266f0cfd7e8ec03dba6e915e3eaaef5f3138c2d787597205477e89a45e209954f51d934d266f5834bea5aadcfeeeeb01e0d85a8a710fd1deecf7db8c42153daa8a73d9a2873fcd7d5c801ad3dd6e0bc424528315bf4e56e11d2bd9159b33aa9c90deb50864650f641964c71638af525fb8e4f261e33d7abfbb9b3d3156064fb9fa092a4d623ed665cc2199cd1f3344e12fb1089e342edb9bba5f1a77d12dfc1baa41ef9dd29601763ba78c5a8659f960deaf01dc8980e656092d958517a8f4678845483893c5d11cb6a0c9c4d9688ea4eb0148ea9ab9648994749f8f377177ee499071d1eda0c1a75c9d00f2b511c061f124c96ebf7a99d06e6f53004e718f886843c698274eb98e57bdf49a0beb215823e624edad833e33f422099e5d0c80a940fa057557677d056c2e37941176580b7fb988cb358e12e7a00cd6ddf266c2cf87426da696eaed009ed2e00bf461ee0a4e304b81f88734ac028decda61c42da3caae114006773cdad08f6556b8a3586bb364a6d54d55725d0bda7163f25a23de765444ab62abfcc847b8c260f4014dd65db4fa71b2b2786ecf6395a3d22047710cca1ae0e835441b56420ce543cc9be1a87ff465b8c32ae34abac566e5d0b55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1a5644d6cdcdebccff4576e96773086e6f6e790f567594c131c45046dd18ebdf168050c0fd1af93f49e1bb8c74263542ee2971de1567d62a92bf6ef21d842406e2e9e19fc5ac3b8a08f500a1fddd0a7e6ffbb2424f7536e470171d7b3bfd00a2fdcce4fc01e3e74f829420a9ef66e4fc200287a7429350bde81c9d89fa72dc32c308de317bd6a53af6984eb3255e91fe3e2f1db59a74df8107185d6e855abdec5c5ee46e8766eb010727e52d0d1b51d69d9b4313298a1df9cc67119a7966eba1daf62a20cfd76d7f72305b581f4442d9c6f3321745f4c61d8859365c6a72a1fb44551555cc486b2432c779fc531bc7aa2eb593fbfa24d1bb29b8564313077fb9dc5fb6a1981f6bd0563aa4d38317c955d0bcd394221cfe3bb06b2bdf661037a942e25e2303b5953bc6f6d433a3a103de809d4315303336b41b61c5a8b8a35d564cc48e2e14ad8111b372130b1c4df3616a4716bda1879d4c4941ea0780d8f1ebdd048427b89073d8ebc81f81e7a12e237ea32bb6f45c1b591a02bbc40b3b583f62a8c683f76c21b38c1249f3bf8a22694b919fe0517fe4e697763f08da07e814e0a641b6d104bf74a50736dad3363a3e8c72f4004059d89b1d6ed2d1a3c5630ee6b4b9d6bdf7380200b00fea9741ad7f940f50cd2937e1501c157146804eb42b9ce2879aa9ab7022f8a81dae63be8039f215d1d0adee3e3752e3092fc336db714abf7f31c429165750dc5a0e3a5a1b90adb7daea06fe3f790d11a666fc8009e5d9a9e5c085614d4231ae842087e9fd4e6dd60cc1b2fb595527719aa4cef52e1d62348820bcb1d9dd9b1b3d528d15658ecc897991222b6f35b11bc004eaef9817328f6c1854e64245dbe74c6c67e230937814caf85e9c85d27ddd7278ce3b9b8e301bdeb210dab32cf0229ba4f47db817044b34bd0fa51b2143336b694afe9718a85581b02a5cd9374c7c5ec0dd66895f14308171b171af6f701b1c14412aa36c5f9cffe736176cd1a3381df77fc6083b3a86720c01415bc0d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcea95a455740aa0c332f86de6d8f76c5de1069bbe00981f1b4f75d8f35d8402989e1405619f8e92b7e09144f2219cbc943ae74ed41d3f3bbfd0217ea33599d17fdd0ca1d53131b781d49559b1550e6ee7e812dc44aee67ca90d5d867b362f8c425b4709c9908e8fefc6cafb1cf96ee8600f28410ddc9ce116d5031d5c9fc4c233d139ed18859c0ea596fe0101288017cd2dc9b6d01e1c5b0240f5f6edd3295a668e0a5092a11b5b86a5c017feded0883e975cdd194359d66f14aa0a4cbac042df8415fc9b6cbcd6237982562a0fa270d58b52f0c6d50a0f35ffad2986d9ce07ca2dd019e0efb9bc454746c6894020164dd428bf5f6d7bb926889545da8a28c1443e45e8c0356316c2a90b2709f388ae6d519582f14534ba2b11ff75e14afdceb90b03d8842aba637b8e253d7de1107a3c34bca711509a9568de249ddf2d29cd8f51f656f37892b20585614f7755d8fd4d5238c3d6d6d56f562d6fc320a6c7d5364f88c662889774a7f4f6f33a90f1307884c569c1eeae54a62d163eddf28d4635bed7c6c905036328373614c74861fe335f2308d9558ce6bd82b8e31fe456ab7bbc0753cb8f119a36ce54d7a75957338e591400fcdca41fdaebeb0453f94d85c92a6d8c0d92ca49e314d560f704fae06ccc8d9264ffddd04065304480d38c3cbd91756010655bf93cfa142c1bb8be5faa7abac8bc0e6b7c0d23eaeb57bde9a37b8fd20a37ef94ed5257597441a7d561e253f1926bdcddf531e311955928021f9932c99d4586699fe2ecee03fd0a041c8c50b240962bbb7de946947cfa3fda2e584279999d1228ba96f0ce529a7a419d1619d206d40014a3caf779449a34078662f66f421865a327a5f39ea1ef1a0af95e00a93629b5ecbd3b8c7f6649363f318d2c0b475fb41374158b284261b22f0088f7e1a115c132a1dd1c725d895b94bd73ece4bcbdbf02efc57568219fbfe6a36a7e44f1722e4c4fa47bf28d8956a79c76c2247822902cde5f33f3ff4218ae4817548d59c3e52688672;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7b2f895cb3e8b7f3401ba77c412dc8bf9bc53be8394195d8eb64ea5d72c2b4d8322544d7c695ccd3a0468a95c2316eae5771f17e783b60817ad49cb67b3655946fd10d32bb1897205ef0f0be07fa58c0bcde23c6276ea9d6a4613b305a50d168a4e377d4ce7245ccaed00a79d1d21def353742607aaac74531959023b7d55c5e49edf4df4be08a684f3e288aebc5d376ce20e11f182e1d12f328eb6f407374324aa40809e131ee14918fc30bfacbcbaac2a6281b06b77a0daefe07c7c4691765363e7af1dba661891abb10d3d5c4df7d4376e142fba4fe4ed732139f0167e0e081e9c33d169b184a2795515339b2e635078d492d2ab95252ab3506c98ec0d24b552267dda06d7fd40c7fa683e106284cc28f5c8ff90cf902ffe925699ff148433739d0a361178888c51fcca919090c7bf57f064f3e677124e343c848ba938858d0c5b975e18d6c41c5235e21ac17ea7febb9e8d90d75271dc4309b98c71e5137d52a7983396df15e7db8f617401c5007a96b8bb8ff66b5594bea7d995a8380f80e074279665cbd1f1bb2cfbdef28295c91bf8ba3cc3dc3cd0a52683429ec7b9bd5d3ad2f4443eb58b37a09ce1ea676b66da55798046d8b163dd79db777bb0ec53291975ea87717eeaf318802c0abcb2d390344dd7de020e5ffaabf670380b341fd5da2e587af7b73fc0e294e794c27efb6ba948b703f9fd31378b04f5873058d80150491c11fd8f881d87d26f8d34633df43f0cddddb3740873b19c8229f8cdd250fbebddd2ab4294063749ec8f1637af841900b2d391db93ef57155b6b75d19d9ab4338c29ef6ae26553d40888fd601697c8ad1ceaab5f044da8b64e0cedfd58f641591301478f2c8ceb9c48d543d81314022f1afac573e54cdf136e6fd2474b4ff294ea0bcd2db602482e7dcf9929d6a4d870e9fbcea9a3198d6d498a8cfcc510864d6652215f11227a33b79ffff1845813c59c6e4297ae75ca821cf33b7b167691a0fccf0a1b9ae7f0340a6f96964f2c25fbc2c1e557d86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he577fb885738b64855d584705e27bac52ed1f9b5c221c61f135d5eb2f8408ed9de6670deee17633b22653b24c5673b6f25db0faa765cf73668bc5d55bf3c8faa0c07ad5663f75ad20fdc4801d19f4325553905767bda4694f5cbf6019b085da8d1e7c51489f2ad25fac7968bb6eedd22e7c380e53b8f2230967ddd3e8f6d7d30b5526e793e0b6efd78e147309752dfc29aaf088b8dc6bcd3aaeacecbf6e5944df8b547283d8fbe9578c9e310e5aa362e7d88d8b4f7f09716d9c62ecb16d98008c4c9f8bc562a30b3c5ad4465884734485c4e83027eb235213635af0ae53679733efa8763f0407b5b95abbae2204a143a3a240ecb4699321341eaad8d4144adc856dc25986c552928769bfa3c324ae6e87d9af0ca080545a64dd8a608190907842c70dea41d654701550aaabf4b00b162c3b931e70007434eaa1892ae43185f0d489d1e5f5ee095bfbd5aab0f486107becce4b90bd00777a2742dd599b07ccf00becfc4c70d5e1b4d159ce2d231b4cfbfb8e58cf3b610aa8271ba6cb1a391c117fea00701a54a20196623570e2ed2d5e9c9bd25e67d681bd4adbf1f4615531f41b2c4de7bac8bd6d8fa950c458d6cf38c705292b2c2ebf82ccf11d74dd4bd70cbff369fdc16d6539ab1119baf9fd6abc0bad5efe187517d5d764c913ce382a35d2ba0dfe8b8637277b31ee49567712c3003bc1eb04e857f921f1f5fa44529e7bb94df320393ea9d9a925d94305eb91e11b39b02e59d37eda3e1ac34b31612add4f971ae7315a8dedb15b68bfe50b41a26b2ad66366214399181465bf036443f1285bb9b1f2b5e317de9a46c13fe2e1153be19a3abc30b5056d7b1d1a6502879cb33c4652d23b3e090649514fbd913810c33d955bda3b6b028011be5c566ab139ddd77aaa19d61dd324a9853f5dcbf7e63ec56eae8fcaea6799aa4a1024ac9633a3546501a9dd18d3bb0dcf03520a2929b9b747272872886371cd6b83238158c92f9510e682ea3109fa35eff85c0ad13402621a06fd9f207bb09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8fb0cb32defb60cf168551ad73ca84abd7c37b49d17cc5954b85c96eb98034deddb617a810a1b4a1334665dc9ebd9e285e4b445458fac95f8cacc657d071a0d8c8a881e0be2373d170185677377ee0e9e6084bd138d9509ea23677a3c50ea08e824cf19fd9476eaf48751bfc7b28eef9a4deaa1b6acf32902d0fb404ca375d3e0106ce819a3864880b5869ad8ea3d250a992ac35dfa8fdc3ee2ce37da6e149d16e37e3a871268dd41edfc668f4b7513543dcb2d058ca18d8d499eb8d284ffff48db0aa5a21f9e357c56473badca74846c46dc7f052635050a59e689d8ff43e4cb9106729f83ce52700f89d0a462d31f42d0c5d378da0ce38bf166082fbaec80d701a951ea1a937bed9ebe63636c431de7ab0ea9c65e4beb07f9a98e8d6b1eb3520c99398678c3169e8417db56f0956872d19847a7c18e7cb690cb822d0e05900fc50da87a485987ea2fe10f9e04f74cedf516d1776793a13d569892bf1b0b4e5b4b02cdf7e614cb74622aa3ede3b0fae758ae183c8abcf8d0d7450871ca73ffbaf49f328450b84b41ba78d1080bcf47f1265449cfb471ea1c37fcca32ab2897f318e621fe3bcabcb47c60e1c9d2aad413733f60f87054098fdf4eaf3dc42c134283f617bf547be7f8b5326d911b7d6a07cab03f4b12d91b19502d90a1df15310a7ac4c7adf2c18b967eff0b77ccb50ec563d727202f42b51aac61f02921917a7f3bc3df6ef35630d8f18fa55fa0c4a9ef091b08a82d0629d258a2c6f209dc36149afcca204c5a4c89128027c2e7f6472e26553f5216d659de9d5808c860af1f249f14aa9c02634203fc0d82e4eed5f654ad8a869d4e6b1afe11463eb775775bf1a40573fb53d554e57f6ec594e0e3d8fa3d542fb2c42c931451989ba842478214f7bbb64e46df616ec2eaeb91500fc21202a0c37f467bba3f369678498f9b89b1e90afd867d7ca78a479b95985b5fb06c37bcc8e86c4f11400d7fbcff4b304cc8dab9ef5bf6eef009b6e17ccb07db93dde509d40c99144114a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h68b307152a2bdb62395e2cbd8ae9b5bd03e1df8dd1e1b1415f18051a388b628819cce23ecd0ebef34a90ed021793cf4d88dc01dabf9fc07c6c698db4120175f3878356a8bffc3d1dfa4f1d2cb0c63f7996b0487ae1890dba839ca028d4fcb0da1a103fb433e27ca2e05c947a1a5a96f960ca629bb364ccc3b55536387807aa49c3af36d88ff4cc53e8870f98ff2cd77b378272f4e0ad61709f3da88c65bce324b5b77d19932865be1fa56d467d0cd7a63aa71928770f1d47891bad6a48137dad0441870399152eb462a845bc988c173328cd15cbf0b2948c73f84e707f99438258293f82f73cf9f7a20df8d87da365ee6d013dcd26d46049ef856cfa8e6916bf9199228bf294e19f2a50e7fe9af2b7daf9c22194ce2ff4ccf81ec0522d43af50cb5ecd01d5b2cd675bdf3fcb0bfaec60ba0f2fd39acc3c0a0eb509b0733afcbaff41bdb9726cf3da72e5663c1e3b96f524dea5678e56f42b5a9950548ee9912de8c385603536373ff0d2c25d3ef67127799ae6194cf321ca02a5dbe26cc72348f03ac0887fa6eb6abd4cc5712c0e630a0b98e40db51b4e69aca589375344390374247a1f9ec43ca305e7d5757d4bf9b041f0d3e63f6b9e57605a64c02c0c14fe3bfe6d48c5beb9eae4930a6c20ed1ad284cb29b7f007b71ae77672da2ec77bb104448e49b675fa002035046766ff607bb171bb056c353bd74bb2a01f271661fecbb144e098372ccaf9fbef43bb5c168289a0a6fa6774dbc2db69e98744e98e1fb49e97e14445f32385db84fc965cfcc22122a0427b3a55c7c8399de30abc97c5260079e5f346165e312bb0591449aa70f70336817b84a42254049bfb7b0c19864062fa29793f1a9b2db9bb08f121730d4818040fb31789b6373149878be091143cda101fd12d095f74056d7fa8748e0c00eb56d35db63ad66120dc282cb4d96172c162744685b0720e061fb9e7f135aa73613ae3fb1ba01eedf1a0a5d2db75773fe3c553e11e8f6f23b959df9b39320f18af96e6d61ed8848;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7ad5e263eac99a8853c4bde5d2fbd62f28a8c51a06fd933b10905adff0c194edbcfd147f655640b66875484d12ee818ac419a1eeff1ffd31f95f071eeac963bf4a43f353d69d385a2290594c7d95b8f72d9d2dfd37bddf2dea3dfad8fb1c25969a558bb9890c3121078815f6dc1474a1df5fcc97b95c414fb55acd7ba76db337a3b38bf3abdda7bf0e8d2c85b6805573874b4e89bf34a92b69a81fafec2b5e9f1c82a04a6b7177167c78f1fb52b042047750345f93458a1947618e33e67a301ad0e0c448cae76863f5fd7963a3c77dc4be7570e173a44b19450b0110e555e0d8c6bfcb92c7e225569318a10ad9cb060f1c2741344834b045984fffc97c0bbca8a691c3df9d8327225fd851cb265febfa3f780a1fa1d2157ba78f240dc15f3875fa26906d17957dbd3d2bb3e49ec1e0197fc9d7c79518af77340869ad9e190eb47493d6c841a2fb8e90d0b3ee3be585b78938f723214d100b1c99e1cd6fb9cf9662bac1fc5bac7554fc1135a1abb4b301e8b9affb799ef9ce1e63024c8e1aefc3bc60981c97f41c27bd2f196eccef0aea6abba74228de3f2a71ddb128f12461ceb1adfd7505bb18f450b3c10b73d840b4eea30d6bd659ef8a16da283fce211d880718b1bc0c81051fda49e4196f4b8127af47c3121c25656e2546d55a228b14830e8a98ad4cd6bebbd16231edcc7574a6ec9953b9d95d05b74bd6ddd6ef3a79310545aa7a5082c4a886950a2bfc9cab7166d9d727f849de4fb7de1397e6ef8ecf85b6022db1bf6fc263c6a69b50148a17f945571860b6decf10eeb262dfb5dfb5563aa16ffc476a7729f9045f68697becdb12fcae519a9bd4d87623a6506d418c9e595eb083fb054bf4124153d1d34aa5425a1c101afbcddd6f54f200742d4fde7e4150f6bc1e4011e1a07624b780f1b301e7fa008ca1befdf541b93d451f784ff82284a7f445ccaebd52ee09333f8331bc623ed29d8769286fffcbec4d949e68801e5ef13b11112796af8c29b430cc75c41b833c2637c235d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf271311c038312e31474432ddb58fda0cbab7ae2136fa9307977c06c44a89a81a59449a30fa58b3734d7a6cf1aa70c7339b56b4c6667fe82200b0ddf817d08c51c36913606087d62394034937f3c8e0b15f9c9889bcb00c166dca1ae0ff6ea62cb899ec7b50c264dfc5bd612a8b51e16715a7838016a456ffa44cb08f4b0831b187d886cc42cdebae6d7c91202bfad984a8eff44b188a7324b060248c12c567e86feea004ab779330213c63c9e0296acc57fcf408dd132c114fb3ac2ce5e188f7b35da6b6d168476899d6418382d505003529539977bdd6c5f5f05e63b05c1903acf7b07fd0d57fd93873a50a48e7808a0330ee9e5b07d79d58e681d229994a4676ad56b37b18c3f1a97b1329b92bb4bb68322bf9b68ff15d7579d30b8e4e5742ffba92e3a6ad222cf42ee09538deaad9eb8d5ba61f947748cd63fea56f419b3ffcb8f571d25a7b33c74c38456c7ef16121a3d8a467f7162ca0e9a65d4ccfe27fbecca8b29b1fd04f02f4ac8cb12e40891c833ed1d259fea67e1dda8e152b0755c90f3d63cc28c0a9a8a690e93543d87f919a69ab84ad91563ede2b4b42c863834e8cdc34e00e49a56ee9bc6c099b7cfeef1208e3e6d69874eb5e4e50ba5eeca5205f09d4702eecee9dc05cf0552578fd0e596fcd8161bb8ef6e58fe3fd15038a37b1c4633a36862db49dc7262b2172b332cb573e56ef475b17f76136d5315be9d62f933b721c70262c371856286be3ab2581ca964f8b38581ea3667eea29772ccd90d16d96b5e9da651778153da5f0065e38077f57592f5e10fa71aacfc9bb5fd868cdafbb8ca8af3817239efff3a22a123bf64daa439a021ca47692abe30e11b494426afa0074d55bab64121fda7755d67538947ca93c739297369219378da28d95e41be6f6fbdf0a1a5a5e95bdba73342017c50b52ce6783a00cf6eaf1328d4ac6c497979f09e6a164623b47b3335a3c95bd9aa99af2b8d12663c9ebd157714da65cd5e6dd8257a1bde15ba0f8bd8d5d64237fbc0cb8f38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h49ff1515d3b44344d35f8ab9c60bc98f760e43b4dbb74a70e345a8646e981f33b0a0c99c2cccdd6fa98ea90802fee4ff9a1e6b17ea797c176e954436bad7754c07c512b82a45f8b554e51fc59f8fa87ba788405b1b5abc97108f38ecb29e715862eba79e3cabb0b27341154d874af9d23955e1f714dece521a6eba063ee2e6b217bd24ef67f0cf10ae387aeb060a57b03bced7e5ab035ac5db8f271bad39e78cbb5dcb336ea9704408f1dced35bd9e37ec696caa4d10364ec59f5cd68d0941a2d93a949296dd5d42dce9cc079b3d5f2a3b5634aa3e391632f54ff63bf130764c9435025383169565847a10f7a94814dd8777b135e6da517f42774f0dd0c51c549c8f6e580359e70dbf18ec5c432ecad6c6de763305cbb0fe66613247262438fa2de15f894b55521bbe563de5d7fead38dbcb4a4d7b67d09eed3f948037d5da12c5cf0b1559a0ce4422b0c05c8425b4139426afd65c34ebf756f6aef26a64b4b528ec9ee020f3ee791bf09c34da38b04688cef126c476cba94b9f110aed32dc1e11c313dd1736bbee6015693287f1e2a856e2cd91b6a4223d0ef4521233b2e3c27768dfe1f391b752db787d754fac3d4c032ba603551f89b97507c3d644510c5c592434abaa06290840ec17ddd12ca9c3de50c448f1677944a55292e401c7f580edeb0a3d19200219c4f85fa75cc28d7e2ae7eaf5385f7b8a8db2f822a967e45dfa6a859e6ea403e0c1d18f5234e154af219ffd106efb698ad677f2e6c50a4aa4c0702285330d67223fd65f8956f5f347d381ff816e7b3007d47040ced2da1cd743f4ddf324d295793bcf4cff8ecb9737a942d830bc6933875441d7312f2219f50a8386081638dcfef18c430c6c4113b74afbe6739827ea029e17d122cb509bd27b17afcb0524bb6f0ca17df368d41f9d26f9ec63aee2d2052510ee6bc02d838b2750946dbb2f0dd3ee69cb736d85a1b219fc0cc7f57779eccaf6351ef5640fa8913f24589031079e6b222a0e684e004a9c4b9c6cba2b43158c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h41d93e27e425c7e882208cf31a6e550b324082e2f687c05a0e147122c22f33c6ca51b63eed40de327aa77d02bee2998324e09b495cbd537417d789a002df896de745b83ca8c42176ca22f093772c6bdf417cd589262a0488f624ba7f1f8292cc8c3bc76964c664dca1cff8e3f557e6e539c1aa62d9d41b926f7debbb959d3b8180756b10897d46f900c561fa31b441c1a9d98f68415a996363ded1f094e83d535f2809fdbe19e495be60f0f863890328b15c3523d7d2296ad1853d38c850998c8b271a09f4a4a2a6c3ce6992d78cbd078fc28122622680fe0b20981f76cd40d3fe2c28155040e26cf03e2607df08aead3be10695f49976c59fb2102650222e507f0f6b5428f75a24b8c10ca53d98c1ce61c9746d181e350aa3a2f8328f88db7dabf393203d7637378159ca7d8d35921123fdd7d9b346d2b7b2da8088142113a167d31aaec28fa0c3e83b0a19156f38e0431fb94fdfc6676fea350fdde94e137f257b358f9c8c92cbc355dc6c2666bab6a5fcf46a387c62fbf63ba64ed0e1f1d211d545ae12a47adc7198fda94a2e30153bddaa11f39011f1f2d42d5575e1782314b3ae7407db112b87712e04e43e9e6d2e4664869746c1eebfe531666a2b505ae4d437f08bacd5958ae195806091ea331d60e4393249295c786f41ed1b583c5347ea85e6c6dfc22ea37cc63f0061da746407c3fa67d3bbd09fabd3f1147358d61b502760575e47c3f256e8678570fc52660072db4cb597a4b393fd4691821e87b784f63d81645a83a62cc19ad49bc612e3f6c296f6ec8d530529482bdd4c32ea4905ac0da831f9d0a1fdb658d1efeeadd61643abc3db0a8098eabcc2c2513ca0c4d7e72e70cdc58cdbee56e7aaa7c8af1a20bf62d5b0cb9d41ed71f33faae3eb550f50001dadb776fbf9d2b49f1b4af5ca9097249edc316f9cdfb97887efb3b9359524f1cf6cfb78ae7293fec33eeee60a1806d66d5bf9994129b22d7b71c095e2acdfdde9ffe53b3dd272f8072f6cebd13918684dfc011702;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2dcc0f798fcf896082e0d5db01c69499b9146aaeec326ccf783068ce2490de63417ee0e96d8f91b38c68e21aa393b425b78cd544b55eb827d8e31fbddf8567b27f4e5b25bd5d854b9553aa01b7ca9efc9a46e693359e9c9c7d1b8721b4dd6d34dd38f6d21da03aaaa421caf804b18f6a74a1b9b6c6c794113c7125de6226a16cd45a87406e75536abc170f81e11fe8952c275eed2f7f346e1af4d14d9a285bcb92828750b9db7638871000caaa7d587e2e619d5445d9cd7eb31e9ba4956372a1a19c216ad1c89c59107d51dd1052299f82ae582708d83dfcf207d2f745cbb7294e0aac6b2844e2f4306336b977bad888e3625ad518288ce3f96129497a977186299a34e6a2c6270f0b28533ed4ec6f3d3fe9168e442fdda3db1fd5325035560d552a87bc1b64a1f4e410e36640d64a3a5cf2e19a8fbce79fad5e4bfc6c97104b1714f29ed24eabb61a7e0c82ed9caff21c39733aac56a29905e688831ff8457ac6091edfc64e33b7e7bf6738fb5a4684d5027d7841e2a3f0288408ff45da1dbf39b2cf90389ec764c236ce987f171f7b10a0705457c59cbb1d088f700e980d9065e48bb7e4bf60575b3fbc4acde4a7597cf166d89ac693eaa03bcc126de49ee2234dd49ff57beddaaed954fa76eb26aefe5a48d513f6a68671de47f2988cd864de4e7702db538664a6478146a628d8e387cb484bb28ac9b473016b8ee73798f96e8184ff965e828e629ae4c4b4fae3127984bb51416471cef8e6411a785812c160f5c7de281d5a3ddb35d9dbae4e1c11bb87869fbe71b0375244b54548439b4855939cea46969977ec118c8165da4ad66c5d9de0b9aaf5b7a491f88b7a3cc4efff400a824a8774c0098e5074e2dfa215cfc8641244b63ec69a78f237e58c7fe8ad5bc41a6c74abdd0679bff0c5dcfec2de2ca7dedafc78d00d200ed32e21a48a30a7bd14594ecc353002b850650cb12517bd654245b67810c78012321fd1c5c15d0c0ee0cb63481bdfdebd9fd028cf1c09b955a30aa8ab9249;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'haab6d4e919fb68ec93982ca4e74f7eaafa8b684172813326d0c019f4a22f299d54e71b2ce44d65bb24471fdff4417949d081351a3822a02a78fcfb2e73790a1e91f93ce9bd0991df42b82800b786ba1676ad03d8b6acdd5d9b6cc8db4c764b5824e762830ab19deb4beebaf601b9d13b3ef615d59cb312199f0c80169360aafe66b324fc35bf76f15843fe44059263cfc480baa0aa6a8aef355dc8447cc0cb4a97c9c8ee98a7d9c160d0d2788bb933c7cc50920fb510c25d204da99cdb68753ad16db9af5284ce0d9d0aca352e4f5fcf8cf3c7c611807c1fb64632abbd4e4ef1122ab31d6eea32c7e3250a3f492635998d99d742ededd60533186a55671cc68940976f219a98885eb394f837f6dd1576d9a1b9ff43b637b94e9564cf2dac9712055dba5deeaee0de87b470fd009b3fc613ff76f262e7ff211abf6df1624e5f002942d46f2a45ea72959bffb4237a6b6812ad984b354ad4bbf385569b7f73ba8d0dcc30def17a9096ad61490fef61426caa01910f596cceade1f4b7d3e87a0a0ce253ba25308f97bb1534a9a376b46aa017efd898492d6651cb0cd8f5618d5d5cd6e3b7938c1f44299fcc84c76728bcb510b8b2c63ebfeb99626273121cc591e1da9cf330344150fa9abac14ea20449a1816dfa6b666d24cc94b341e2425e74784ff34b4e183128be40ef8868ab50db3cb25388791af613aaf6f0b5449bce48c9052d0c0d9edd22a83254691d8bdabd6b81929fc185079e9e85bee569671b76b09571f18bc419a3b8143ff87a684cec337fc3b6da136c3e91ac735427c7db747eeebf961cd1e961c3a0f2d278044767b7775ab27725611d5a9b8413027427d4831d2b0ae378b253214e04de87751d1ec808eeba62170c9e74a3e6d7d8c42bad3bdace2596acf44cdc169b50170ac686f8879626526e8e2e3915db5a3dd8e29abbd847d4366d38288dedce7952c034f8f330f7a12c2d99893ee5e77f82232236dd4945e65314595e40b549c99533305bde724995d827e495bf48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4f997b8d0c586035fadf1c71c8e31af25fdd86eaa55a3889246a27bc93a8c35093c4c30972f0dd73579a94421662087ddc9c12234968b50c7e70b4513a30ae4ccbe22e93f63e1279c7e94716c9bc8cff8063632dada0c02983f06cb5186a8ba34de43807728cbe3809f4c156fcf5f5e96e6ce6727a8b1f85d988e562bea360dde09668cbe7027cf6422962162c47dbc4395c201f7e111b6ec4de23bb21bc04618cfb585c20c20b936fe6ecb76f80ad72aedb08872234649b33abfadb74e537f035f74d1f2a1c0649094db401647a8325e841b072aed2d774f3a4ed0d92c20c69898b1767d6d448af61f66b65a34ceb017dd8c6bbd73ec69829f67555a64b4065ff228273a207c5c7ea66a8bce38d7260b2f406521e25b6f50b635c34c7d68a84fc44c0234a0faf7c56e71ae0c193ed7025862342cb685c060f24987e8204f148d60a460312be04bfb7b02fb97c947e2e215281b5c0cdfbcdf87f7ce399a8c337a8b1d7dd06f3fb015c02acd1f2f6b777389fbb66a0736dd553faf246ab5afcc6c98263a37bd28c63d94722090c4e05667ef67045a05876fc20e6a3b740c1206b71f40def66f016f205fe0b550d64ed76ffce05b05f00cf52289409b3fa5006646125dd79e705fea2111ffa917ace7d1554e0ece20144c6855a1e9cb78cc95a13dc262d3a83779855ec46d3c4a1af82742e36a0955860fe5eea3675d3da5029c9587fb806d8a69c1cb8c07a2d55f9b407c5b1fa89681fb02faa085d8587e6185ab64ab6fe767369c57fa0c12eb022b9d09e1d253abeff9e07ac44776bcc050fa87a809a5a51453a9b9675c6e6c4401a94f36bc9334d1ac8748db30c66e04f77667dc18fab46a2f8422bb1596dac261ab66474083493e69130fc18b369afa50dffde997c003e050437b92fdd6336c48029a31a3bd1fafb0952254887e0a641cd117e3a4b5da3f1f9fbc355a2f349b3ac188f2a5c8de1a612e1e06b8a4e7f92230e6c37aba726dc6ccb1cca0e9530d194ee54966d1844e1d2565f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h71fa9a370103e986f7e59ee3f21c635b52bdedee9edfdc9da0d5a15d6e9318a2f0c2d2ae183242d79218f2f335d30568e814561593d355be970afba470f1914a6773d082c5198b970792aaa64f3af3167a22dd40de7048cb3906171cea9027979f10ea7c4277af1302c162d51eaa40474e40c16ca1b533ad71f07b48e9090c503ab3182426517d3a1819a0d40c909892808052519ea51ea9e777499668de02ad103f22cf687d0ce00578820b23b24c0fa541aef7985038bf8c6ee94306a3433bc0afe8e619ae2c8208f1100eafcb19758934561f2daef7044c4d891d88f4ed8eb0dd62cf6c3cecd7585214207c9692bce5751259ced192640961e7d52a540c6db02f9cd7720b2784b93415d3020c4cebaba4390097169d7b59efbcf9f1765c6ee90929d62869ac74d71e75c732cf665374c0a8ce9a15f7e54a3990c32ca6c2515ad1b82a76d59265d69f014c524158428f2d779e93e4c92dbcf2ce4f632cb32346dd2fff32709fcc3b26b7ec0e36f04643d1d09ca8edc1feeaa9175b09c6e4f1baa1db25e7ed997daa0586a212263ff87ca82d25cb8137643e1dbce4ac33559bd1b115b61af6cb6af6352b6781cd9b69f9ca569d5280469b039936f00b6189c4132bc6b531366197986bcca94ac9ad9e52384a7b7eaf35e0d7415b8a9a963d70648a9c4f59141474d7382a2528df15e93dd504442b74038601d0dd0052f063e517a6d083cbf2bc223f88884dd7845517685c5a0196563bc7fa2f4e5ad0924a1db4cadf9f203202d1325533865f7959e1d294e96c2ab2266ea5cb2c1f8d747f3d058fbe7820de2477f81b795167049c534e5d6e6b805d719975c81960ba55ed5a24771efb7b8525be02492b76eabeee89f5069c343dc9541cbe313e0a5895b8ddb2c1fc377e5c71cbdcdce8678697e552c7d289c8d5cf5dcdbbfa4f3a8ad8bae98ec932f194ad16491a850cb0ef669471749943ac08221eec676593555159e1838357f23cf873f1fa90a7773dc024f817648f3ccfa7f03339bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9f221948af8325e3e9f8b344b41d57b4f3a1e959ef8f59c562797cbe3898f16407fdbd77bb86b79b7bdae4a72bcfac6c1c4fc07e8245ffca490ca1e2233f1ba60a3cedff4bdf5fcf9ecc37bb208ce4b5af9222ff7298187230b4ab7b890568e1706dd926e84cb8f39b07471f5efdb1ea416efda293da62f659544cd94e61f6f0d47ccac3e099d780475958bb2c0730db48d5f5187c99731d67ca7bf23448f26b3fda5d28ba905bdbfe56c77416cd1b150785d35898171c68d42eeca2cb036269ffba4ace5d41ebe30a4744c1f0c739f7c68b494178c5946efc368c81442b855135a023bf6fbebde03f68d81424f489adbf77f40c0cfd22ad1c62a3eebbe2439bbce936463f3cdad75ce94589fc6a1364325213c6a1403b65013a88cc66dc7b39a65b1778bc8d59be82a73a83bf06ba7d26534428d968fa8dee2659e16966011916eb6d7d5c2f0ed0dbca93e96a1d22b120c4f61b3cc3d684ab0def5163fb528a64dc2d344429fd64e549854cf9a062f912a9fbc63e4ab3a676a350e0db6de45e7d2fae0925ef77ca021e078e3a5c4069e6b5d9b0636357282882f575a7aa7fca5d11f171684a61d099d23ecddfa70730eff3a7a74a4c46c70cbdbf12ab907e2f6e210fdd4275c06a4f588d63330b2ae40dfbaa026dcd342d9cd5fa59f52684b546bcc1cb4949d84c6083bcd4d79f560193295bdd27825b80f94a20f17eda389108d33d0432acc59ee369dcc4145e672a941e3ae1d1fb01640c8b889c6989e1c67c920bc786541fc0fb651833d26d57f61ebb8c6f27761cdbbfea3a9e152495c21cf1b603698274328cf353797cf5e1b8748b0bd9b0dea5d0a692344551248426f39da6a5fa53c4c527d9591e3ec963c7f48e19f4a3d2b6cf2b8d87195c0dbb48d5f21e3290679a80dcc59fdf1cc89f7d030a9ebdc8a5ff6c9bb407fe65c92cb5845f2d78d59aaaf0614740ea4bb3d09677ee3e6363bd4d8147ba3e16015f6c26c9672b63cf0749dae478d78a1931dd06bb865d83a34f9b9872;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbb07bd7540c48fc3dfa3a295b0a44a4a393cb068788366da959918632fdf5eb444803c2197bc64389ffdec3b2c2a245ad75beeee3f30f5fc2897dfaf9cdc1984837619c5d2ba59c98192a7239d9268d63be3178835e64e410b7823e1dd3b090749ee39d4c98144b2614ba7e13307708273f2dcadba9fc7fbf9f882916a9094eae4182d5bcdd238b0f5c191b9bde4a2b47382ea4508969dde8f83516752d5a35e7e8f9263a75c1ff5b57ce72cbcc1c9f637e7849f32a2a03677f693bab8b76b0d1caa3749077399f65b631ea0b07ab9b8c94060197cc68aaf1dfa0b236b1bc4d20153a122d162b75c84dc72a0445a7b26b6f4cbefee83799f47ca2c7c3fa9a096d463f7201e36bbece27bd53543ee6b1c0e938a58cb9cf1e8df090777aab529bae1ffd633e837b44c068a79970a62a5b0917105f5e997c3a93681c0709ad71523894a9b19aa268c8ebdb79d4bd0b9e98c19080910b7bc5674c9f472c80f344ec22b9fe6658630bc8f2bfa2036b98f89bd1cb99935e1c6e805805cb9f8629c29b1963162c385eccbfe38faee515216b866ec87c631fb1cdeb9543e15ae4b692315ce51c0f01ba0498e457e65b56ae430dc424945be7152158da18af82f00ed61aec1f01764637eaad029b3b43f3ef104b42bebd54acef4731de91d411336c91ac3066af82c3e855a7df1af79f63cdfaea64535080dcb8404abe3281c414ace730f7bac32fab8d8239dcdc41f90eecaf60180dfeecf85f9b803fdcd8a6fd7a6be1ac6f50765d6918d6df82c5d6142ea1fe8d61faf8fc1e23fd84d4cd75a9c9aab27a7ba4e8cbeb77c6115d468a277b137f74b3fd529cfd3c36cdccc2c97c8dc5698226a82b86cf7a840f8f7f1aa08f4b22e7fdfc666bc87d79c1fa8d0b01e36eabda91a31aaaa4dd903f9f57b0d3fccf7731b4a65488ff7b77d1706dcaeb0cc3f53e32a7055914a19c27b595aa2184691c911b70feb112a5b4b840a201da494bcdd529ef071e856898f08249399bbe305a584246d3746d5ecfd35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h61ff914b8bd9f5b717fd65f2bf9d35fa3358d68e079f24244e588f3ae47331f0c3d479db0b888a397a734a8573da968b5f4fc6a6775df119d1654b54e43dbd77f223ec231b32349bb88493975292d6317056bcd01e00bb943e97ef6d7b75dac1fb7456c1249dff6d8a70edf743bb31d6a28c678454885e0eb54063e14ce534e617e0e85c1d2de5ede226d2578a6133765b642ab91c2caa3b3abff97279269b581d47fb5acababc3def46c521db49d096263abe8582207b56b8a16034aaedd94bfd6e28189484849e7e075cd63d915816e177cd50ed7b4f214e425cddb3cb53d39a799123cd913fb5445b803ce7e147448368a1b3bd13374c36795fbc870b4b5d0da5858c528ba7a6206db1dfe6565f55497bdfd97ac209b8ae2d7aa271bb28aa5ba3a8185c6116501b98afc53ec3bbfdffefada6e72e0ec0dddff326ef1760a44669349a1d94381d58c780cbd8f95b841e3929d710ae261b4fe5162d834ccc6226875f8be95c69d91909ca2b7d448aa2d902a18743f8036964b1f38e7239fbfd1d6541b577f9dc8b0c4cec011a673f3fe93068c213bda873389b24f3205a478ec8c17f831ec1db16da65f0cd6f1a6d34f0ac01bd9dee47c3de3df520291f2a12c546995e23ac5f3ad15c0afab16338c0788f28d1a1b8ea90d01f502d0cdca14bd318db7f382817e2fceffb99f2485dc02a162240869ca96e9d8fd130279d07d0f14df01c1c890004a770c469c9d6263d69c079ebffb1f8403bf7cba901ec7191570895077eaa5e7e357106653399e63a530e548d01c0fd6bdb5be5e1342e9081fe8e1654c61b24437260fb4bdd947335e476a9e27846c3c421ece916b0376f5a5096314e70a19e77fc03418fbfed185b33f0937398aa2f64f652d25eb4e76fa8cee00d7a8af2520cff107ada60b3b0220f97d796c5a15ccd6629b955bd377a236bcee1e09631cdc0f9bdfaf48700d793f17d71a3835cfab607ff474421fbcd0a83f580faddbd4ca6d652b075c1c2ae67e0c5aaeeff495cdac7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hff604b49d3fc5bf15e9aa19918c5dd2c7cbffccf923c4db7e9f127a86bf54a152a49a24a5bad5ed9e322fd8c4962e4552bf549c9afee1133858dfe6aa191bb93d7808dc2d8d55037896acc0687743b807dd56bac5876ba1015754abf8b3942d9d611bc8ee0c568ae25e2adf8ff4763aa5f4d705b5ddc8eb101b97554f2e6ecc0636e5964c5de6d9f167b321c9c446cb711e46892012cc791001e821a55903c4f436111e2611a5a3556e3bfb87be21e0e0523ddc428407e6c8361ca43a193dfd126adc9d2c301f30f0b1352e2c04cc93c903024acdd47cb1751e3031c497310d196bd943f5229977a84450f9a7646edaf05821ac26538f6032db68c24fa6d535c0c694509d179e56487ebc3189e7260b280974efe769b5a5aced9be7e78c7ca0f0792b414f2408e474d747502002d0dc14cf1fc8bd873a6a57855a2c3fef2e71d14eb432456a579ecfa1eb6b3a0a52ea2d7966ad91ed0490987b7146a909b8f9a8f84cb08b3b50c68a79a4442de22c2b0b53401a09c290751f6cfbb7e0d590ea09a21e2c9577684df663e486e6407e510f302d30913e52c38a64373a3994825d2c3339d4a8975b9b2e46cde0b572aad71495dba19d92c39e702db1ca89fe2f0872c4b760434c262184fd4d21312a87434b554f987f77cef9ed56d39af73d4130c0cda90b83be6bf44b5bce6ada09bf820f718e44d95af61cb310cb34e9e6809475c14ca1db4c47aa1162959bca3d8d47da6e4f1efcd3d3300aabfa9ded63d2e00241bcc04384003f15671482789bb58fe92e0eaf5264edc919edc6ea49913f33b796529bce385aac700d5df923330563e9eac2ed079e686ce5fad15f139cf9be991d51189630edeebbeda2c4455daaf974382bd8f44a3eef32fdda9c68e639b3db347e34a264d18466c960f77bc743789a8b3f82373a8108c2fa95064651b79b591dc7f566b9b92ee8201a591f837499dfe3a643618e673bb807c24df2ae2c4b5d160bb5f59a34e81478d3cf97338c630bafa683d871fb3f908;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha43ba657a63aeea2bf93574c499e0f08c56c9a7e49bd868e70d79009b915a91f2bc560f272f346b74b40b09aeb10f1fc7995733fb9964f466bd73c8dd10b8453958bef6a081425e795b666581a84dfb38fd17c35a8feade63f5702921b6b5eb41157820d5e7e6be7d9181ba49688246e1fcc564a96b473673b8e2fb7bca7cd0c5f87cb289544ee9927cf8b197c43bccf36e4a249ccb1af1ef42423ccc947c1ccfdee3cd3f77779ee95634ecea685e595d6fa19c6ee37b40883c3aaf2334b76fcb778f6ecbfca5d0e867eafe19d2bfee99da746cc91a84d516e628173b803f596309aa12501ec2d78cba8058de37710456bc8c800d701c3e31d0cffb96ff66237178d37f17abf59f5b49ff1b0805156a3516b4e043a769c320aa7d481f12b17d3fb16f77df80ff7889cc430de9f41c1345f69188c43246226e419a94990fa61ebf130d6b5fb5e6ed4da531a0656ff169f59e5bbe05c74b024c6e438dda0226bb4c9e7ffa2d72c075577e46c3a192cfd20797de0b978524ad21c1449a3f48f122b2a9d2b87e00a743447596aa884ec60fbd0f0b0dd3dc5517ec68c54474692e807d03dee0df45b3c971ecb49304c4c2364e5fc63c9f2404641171b25781e81edaff84f3ff2a3c73693ea16fd099b6a79551bf11381a108fc1243693612d6de5a51f47648150d771fd244c83972dcce476e4c0bd711db0985ef21845bbad4c639d82b84dfcdc76fa00016897573f886e7408f3b4ff539bf70354dfacfa5e2f434370a4be10e618a9487dfbc9f733ecb1d1cd5ef4978d8aab07ae8ccad039cb5fa8e68c944927d759d15fea7c463845504c5d22b2a0baa1753380c704a4461ea4b57e2f75f668d81768c43fdd01331f2b5e76ab67dccc56c21e4189e0ac52d51a0bf6cde6e3e6c810d021d2fad0dadbb08ae1ca74947a215e530f4b3c5a8985278d7142b94b69966c1e3381dda708ec0a761bb2f7f7b0f0fbdbfc195f8abfe51875a251714aad23860b799d794c7f4316c423804a5134d09c92aef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h20757ca4b4e7cfbe55afc0b3e61f190cca27db173daeb822f04519bb581832398ca42f681e4042a649befc29c37d8075078944cf52654e07597445626c20d942110c6991f1964ac3c236e72cdc32faf48332b0db5501445b4208b5bfcb9dccb60a1a28393348caa70cc75d0bde500222de3775472cc1fd963b113f423ce89da45edf8cef2fff0cb1ca5eac965ff03ef1c8182b7d6ecebd4ee069fa3b25c4c068cf1eff31dd04637929ca534286c25b3e7994fe4a327eb6362f84d2df3103ff16cc2b2ba985b6492f426a81df419cae1397c8389ac491e45032c090d14afe89f5d97efeb852b4f85edc937af53d7380eda170501d6b83e99187dfc81648ceec4687c8a171b25d7f40cc608fd1f7a127a6712a4b9411e48f1fe01ca99526039f217f8109b9dfc979965e312c8fb9f338216d54d13ea762cfe97ca70ea1ef03e9e3634e9b6bb61793309718b5573188a151f3e82cf3fbefa28ddcff4bcf73ee1e7a44ff85b6b4075dd1be7417c6850fbe17304ed4214c9e8698c100092945fe2e02154d2261fe8542c9f6f25ac78e643b86c43edebb2ae7e86212fc195beda9a1ff798becbf243053bfe04f9fb457247cf16ea282ccd54557611642c5f60e4528e1e1a5ed8cf39efd28d6e7cb34f6674b420ff5ec13009fd91885625b28819ec1abc5a76497dfb5071e12b6bb7aecb0d505260ae379118fbec61d642ce9f7be6c65e5f553af1d512923b36956eaae2c28e502b50db8e05447333c71334aae142771bcdea6645bf2891523afa482c2306182946ecb75b429f2e5772fe033956b7325ee708700109cbb2afc355eb0b180b8d7fdf54b49690fe844d3ef123652fe83d7ecc8807c5bfc228f0dbbc7f297ea34e926a493211364a850bdc37dfc759a02e106519ab99417a6e17ab1d58ae7a0e360aa3824e951467080a6eb4bff8dd242a4758dbb69cab3343bbe6c40f5e4d5b405e9d17d539aedeaa2ccb98d3a2210d31bb8c4a9aebb7c4e9a64796140b7e28474de7b2cbde0cf1df76b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h39254c59d9bb53c3916df22223fc35e4ff7fa827279f0429cee24486fafa1381ea77451b14f2e4683c6cb9704bb98a3f9364ee3d754003719d3ab50bcebeb85054fd3b3dd6f7a4249ffbdfac83460751efb81146e6237410625397d466d73ccb54070ad23aafa21067ba237197cd284b64120935fd5fb4b641b0bb156b73beb60907a1ef0291f310c2e0a36fd6f551fc8292acd2deb56af6a80f3994af2e7779eda21b2eac803d642626a8f566fcb8c79a3ab3a5ee7949c7f6758f512579a825f16cb4b9918462bd3c01c7b0a9c41931e52e9db3483586cba1075b0244293108cb90e883d4bdfc159eaee26d224cc33852e90512008317ed4672867ffd728841f8fc409248ee5de7bf9207e1b0b676b4626a0a964bf8a7efc228579d8570662c71d23d4d1fb785de5e3a2dcaec31d053379446be604f2df063954085c10287a8bf9b0f84cc68e68276aeaf812bef83bc3dc319f634bae62be30cd7fee8fdf4b360d458f123bfd5cacacaec22df35c8d75bb597a0868e4ca275189197fc5ccc31455b15f44b9fe8dcaefcf01b5171703229e36ab97397f3369e0551b780c71722959875e7715c694fb6a3334194b0d90208c94b2b09ac3ccdb413c295ea54528c856fe175b9da2d3f85b986a2c8da39a3e2b461572dce2ad01ae5891315bec463b3e6b9fc8b4e42b9e983906badad9fa590a2c50e52f86f91d168f0075b5110e27b0928eb64e1a08f46fb74e494f31972432ed7fb22ba5c3cf12929ec9fbdcccab08850b1c13d9f692de0474d72c5bd10c34b9d5087eb624997ec36368f392449b952d8276ca960438e8d7825172bef26d2c1f75ffa80d24269e0a799ccdcce782a9654c58d6bd88e3e32cd0e5daeb684ee812eaf1be43f0883a3ea902dec9229a6c0f3287acdb357b87d566b1d929f138b40a49c04266ea8d6dad407afecc576712aa91f2dfbefee0f193f4e173ef0e3b37bbc6cdccaaa73249eef2a46a9a54d010265a7e9d5ca877c9c71e24e3ee50fdf3ee1bafbd07002fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf6096a4f5846f073cfffa5cca471b198408a0e5b42d4723bccc4e079ce84863022ef3b7b206e077d463ee7797b27136f36512a3d3ac5a8342beeb7f8a37a80523052eca8b2632a116a6ec1fea5086c1d86b6356a267727fc16fbd5d658b7389bdc7eff2cd09797a46ad0bc623e1b3720a553536badf52e52889ca43680e54a72b9f49f02998c85223ffeb95ccaffe22baca875f7f08a523dda39810d56b97e0418586c5ffb3ce9ece27f42b0f69f106baec9ba239faab7316af5a72c821202ace12778c59d94d05f7c1324804f56a340370a75883b6f78885116863efd7cdf413dec768e6f87ca1ac2d5a3d3805d810d38653bb483e22844e582edc3efd1ff147c808ab3353f6bafa139a1ab3e1f13a777d4daceec46aad9e6f9923e924f46d3f8111bb340e1f4b764989454e2eb444976edcd3be6dcf977ffd7e1879c72c3c1c877a9c92255f1d3dc6d25774a60a980d4cffca246decc41563aa48ddb37dac7dcb6484fa64412a3c4399b438b6380f3ec8f824a41a3eb4ff58c35c01996480c3330dc09ab94424f5fe825bbe34f0656ef65a198bbe7a7335428853e2358dd269e898ec5e5aeb9834b6ff42a2a140ddb14fbd97fd85ddaae57025af55c9cf83ba5ec058f5dbfe85700020d8de0d5e9e56968d00a4e3aac6aa6727c3c8d4cb4dbfabd273464b740beea2cce9e696942d3361ff885e5b9fd1336022d89b49b99c9f32c57cb5f55f5d8f2adc3b9d9e813cd09e80d9730b4c80ef2382d2c6f1686f0edb69b04e6495df5b97b89053af4bd30539d287d49413d96793b24d0c350c61fd2ec79b48cf5cc73692278030f2e56cc7301d807c0535fc6f9141d0680d799e8e6732eec49b8f4a2ef21d68c558372cb1ed6a6a8181d1d96ba354bda5dcf33477670c56d3a7925138c845eeeb6b609803ff4a36f76e055f28ec171a6b23345eefa9143a58254ea3af88660fd6969d4b25518aeaac70d366b79e534a13c409c36bdada3052b94ce20fa47fb720d66ef2e122621738379cb96c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb7d46fb4c6402996a3c8b6486beb287f29773a504bf9ecde43b2880b5f90edaf18476d89dc0f44b32467b52caf64d03a51d4017a9a0ae118e0b5ed5208366ce23ea96de7f8842abbd73f09f10f709533d6ad4d6ac13248a7a2056df59a87081f68d5c81b730cae80f86d15426107d783c1aec61f7659956a21fa3c40ca18a9ca7dc56a50e0dc537f69ddbcaa2e49d78816b68abd5c9445088e4a6c21dbcf492299290c4b8e3f33833ef690ddcfc144145608e9961ab2f6ed8d7ecc70eb6bcb259668ccfe32e0a8bde683f1cf0d5f69bc87d4726549ce13e1a36cfc9f24ddff168bead17b529167249d261d8c66dbdee14c4a16e8fda2c515c629cb1c65f0fc26a7979a4cd89a29fdf1a22943ca3c00bad40c748e3b46d0f31b1a5d8f83b0467234948af8d4bede05b2bb6780cf46b7f4873f9f6bccd946073e96f722827e1950b6c17f76df72faa13af1a31fd175e4358de55b4176dcb5b9c73cef687d84387bfaaaa844db82188477b848c893b2ce677fb06ffe9c777d4324ef45d540ba3ae9fd38d6b791a803d6b1766113cbc868a8d9ee9b704fe92f3930619578302f78ccb56d345683dba2a1551fd682c858576776d54e0d09cdd63224e66f64de8b309a04be1ad29a13e8078a289e98e137018ab71b9b02a2bac72a785902ffabcf2e6ca2c2de9ea3c6a470eaae139dd66624b5d689d5c1c3ead756654a2152ca250491b8acbeb290046728eb639b9b38d3cb1c57c92b131a0aa48da2afa81348e4b8580fc6a9a0ce88c987eb83998c63b927381f0761eaad66b573f67c21f4b4a5cdf628ffce8fa4c4c9982b8ed21697eac235d8efe94a4fedb73993ec808311ee2b814608b393ea0a2e713c26d1da438400d9aaf19916cfa6329a24804b92284e72b851797717a6a170f2dc9bce50ce5e3c8fee9c6d79fe1cda792f9d56d98c0bfc98b837a50a8f0f63c1229e5210a0398581be99faebbfbc34fe30564fac14fd182858893df253dc9d79efc62697a27fba0f909cbe2fdc53c1b83c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4f34c0c8dd40a5659afaf8fca761b3a0ad0210bb4042f43ed970abf4432abb504feb14f4092ef015dc11fea7106793e57bcd719762f5d064744342e7db531f52970af8eeed448de9002fae48eb0348f8cfe66ea8e2b1b51c12b2848ef3042f344b727b5237776dfcede24d4f6612ee571ac1ea45472b8dfd98ee1ee2554e997c3f6848a8aa0e71512bff73ce4a4498be7db160962c27ca6dad9a07dab8c5da28a8d77c522f1c0032b0fd8608b55615c220aaa248876a8fa8ce40cb151f85260505dde12974c8c08f5e1e15745f92e3796256d120e3adced28aa26c633e3d4eae186300842c7bab6a52971612f684cee0d9e4b64cb793775ef49683e455e0ca7d7a01f486f9c18546a806a8e290527e4e1c703af1b39d5b927af4f344c06ee09cb5052b04c8f867fe58a55ad314e6224bf05e55260e084addb7ff616126064a23b15512e320d53ee12c073dd74ff199e4048a34cc8f8d8b96d58c4e9506e8e8f14b548bb63be96e1656bf31d17239800ea242654a2f277fbcb99b3a1b96bb7bbe4c95506c22fbb72e2afde499c67e7a1c31f61d95566290623aef4d48bc00da1c42d75b0d91c86c4595c9aaea40b09705eef4177cc833a366bde45da004b6ee2e77bb3787fc340ce70bc6dde5e062b06b66ebc2669ddfc645c4ef976f3ec74fc8649cc8d1e532192a52541ff96521604bb27c657aaf463145dd6ab4c7a1a6fbdeeeb32e1b1cd9030ddb7187f808e7b51c501058d71d9d923b66c44adc18e24a681f089bcc1dfed748a5117727120bab5f58f036b6e9a1339a25f67dc643192f973090ae6183827443fa1c5d2f9c6b45412c690bd78d686f883c09c0c86999769a5466c9b7d99e44f92c8fb368a7047bcfcbfae7fcaf2e4e7b7d5b78c21ec0b1f0d25c91cca7d771eb1eb26ef87415c9b91d13f8745d6e652bc62329fd9d43376ea36bc8391578ba0fa0624eb2b3343e1c67cfe3852067713a2eba9ec278ac7dac366982ea3043c6d431a51c6e982d2b7ad54fbfb67360092892;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc1a4344a53f540bb6c97633d987c5c50b2c754350f1b7d9623413cf6cd33cb0125797c208ffe6d73e7c767b571fa383a2cbec6d2e47d2290e9a2f4e9c79e4b9e16b44e38acf23d401d6dec9ba3b72e55bd293fbead5f22ae966df31659ccd2c20c6a49e70d8d56aa5a9babf6b8c5481b457dde08543eb0a6fd049acd62b1cfe97d2f66eaf2a600db3ef6da3b8e9c1b18193df6633e601a13c150a6f460a088612621891fc4e1e15b53f9a0767bfdc24943200da58b6bf0dd0e9260c82bdeef916bc893ed9ddf76368e3eb567459e6e504247dc78eaa043f92e0fce6c884c4409c96f9090e43cca1d20341c57a0056f9681ca06b73e75ec078c9631c06ea0d694e3f6fd380485b6579091e6f11d68227b04cde84fdde5418768b9c394f2f828f6d59fd6fd942a5812db1e7be1f6e764fc6d06c064a3b5b6adf40764a2b7b6ec31a0286b0400244cdbfad40e7d46ebbd1ce466408bc3a14a82aaae7e845fd68e8fb975fbf2453d7bd6a5b968cbba14b1f5a39423e137d1266f920898545dfefbe6ea19297e1b06a4e0b9599349fd1607ecb3e7b4260319fca13b15cf2dd7f23a2847e5a409d4e86a852858f8101dbc4b05b2b8fd3b947b0f05af53bd61a949b4c8790d083bbf057877a170a0660c2953c90ce535309f33482f7c366e15177e2153522ac1a754dc98f46e0bb4b2df96a601e7a40fce8a8c332c21c9adff3942b2db1d8037d2eb9be6c40df798382de68d4d648bea1de5fa7f510c84927dc05afaf044800393c5ea2d0c15d1921a5557ce3878e53537456344534c7afe96a6c4b6bfec195758e5095f3a574782c24888717c470474fa01ab4d0d6d24d36392fe87fa84424fc98f0dc8fca3456ecf4f2bcb3e35c1ccdd23bf3cae36915588fc385ceb43478c383db14e3d8626918a972534788c91549ac3fba24541ca493a1ad5861042bb5ace7745a19cc86bb70a558fec16cfde1fa466c032640cf2f38cb1081626941d58aed2fca71289a6b9817c82513ad4a6133842d2ed3857;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h10d6684e7cc1e39b4bbd7191f2878a72d71c864b013eb60e484b07bad32c4102dd5860c0e128964fb8276b20ddb4556e0c0ca103aa5877e0faacb8a7a7c7a1e06bb8d5f886e28eefa09c4fe510797d3160c921ba4db53844402c4a5adc0f9ac1bc533f3f3a622cbd0ec92d30e5f0b1823e4f6ba82e65417670c7d17101f2cf43985f0f7ba368282448dd191af8b01afc39c96ac9a137b726f322f93569290785204f6a3e0334fb7740e5382687ffc6c76535bf9a83c42b9bf276394cba93207f145b5cf5c622efcefa225623ccc830895b56f062a8f5004b5a23e3f86abcee7d294a47ce1f9f698e4bbc6d18f8da8924555bdf7572035ece9958567a9e818bfda93528ff580e605221e758cae1fc7b8dd07baea9800f01eaf9a0e1002d393b1bc591f150736ad0595f05905c1c4f69bcb4f2346277505685a56bc6d8fc56e5d6de578eaeffbc26f9f0647ae1207fc65ebad8a2a41407d630e0288542d97476614ef6adf5813fac7be085ccbd750536d66158fc8ae387b13064171f0e109aa6ad4a7945e76cf5347a678b2a9bc1446aa8520a12884e3d17bfa834b9218a3bd22c57fee417cc2760a68b118d4801525cce4a30a5f388f31238a6a3c4bd6b5a9adf6d960ef44f7a2b6e920fb2705e8b00ec13291ada9214df396455e2a54c92187c40305864bea2c56a0b7eb1cc0c269c3172b6b1bd937612557c121b682191484c4d98ab7638c56c2e34fdf672536fecf0df35cd5612cd228da3d36ae4aa007ab1df65f759fd84ee904fa0d630da0d296e76e47b6cc90e324791e0653b8b41b82a5459fba63a793b587a1286da7953d5b6cc2491bd3d3dd8fa787877e046ac714bf504d9bd548a3ff4ac181b4653ea364c9eb45b9736d2a2e63042fc8e665dd9082cba36e2740f4f139cc5a5d5cb884bb940841445f090a22d09c44aaa6717d88865591c4d428cb05b1de865c925ed5e74b763df164cf957943b2d69a538616f44f1f090cd4064f7f667622efc515c80810cc7de81c75a2a4de2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9841adb9fa4694b4871b1d01ba5b7f090fd0100a6b94581cd326a5a17d7a91018e627c7ae930191c908cbfae54904aca3541753e7a455f340252e16d4f3ceaadf0f36355adc25f075e79356850ba715f3356bf2509daaadeb9b8c2556f44159743c946bbff866ba5f36a4044f2fc73fd7c293a165a8e657a56e96f723d06b2bddb4e1066af7d5ee6fe2b47df803a76cc05cf0963fdf254572f4c4e3f5a9298961b837e53b8425441652069b08b44a3152cd6b605884ed2f5528920c4f55442f398924aecd7882330272b88b2b13a2c6bbe5f7a89834b64a922706fb0aad81cc3354eb6cb428f283884f10cbfe1ba1bff2c75062246d9d9d6d8670ddd0343a0a1b315f2c185731f4ea0eac3fd67180faf46045065ddba6ddceaef201e6b1725571a91cc203a223e7a78baefa6016dcbbdeb834d01e150b8080fb8295424936637a416b1ff99dd89217092c36abf74da69951f0b89c402e0ed34ef4f1792a2794b59786e3d6af888e8692d0874b0ef862afd387e3f923f6211b45b7ca3699ce3e4d439832aa24e56d55bb0eabe1873310cf6ff3376ce629448990dae3d3817345924a29b7c56e3fa50d02b10d8b5b2ab267cde59fbfc11d93caad33d8283126637c6ad97882ce0b1c656f58dad88f52eee651a46aa11f7ce7bdacbd7c167b44d9e3601954a5615e0068f99b8d19b9999b0b0a907c66c323de31ed44912ffcd111d2496c3a70cf6d4a3270d79dd8afb4127d3d7070e05c9787210cc7abf96660cbc5c078e050a935a28601d94c2697a9879cc07b65acfd2c0e2c36d47ad243441a1bdabc9361d82358b1f663f8332500c72de529c958cae6bbf09b3e76a451948019b7deabf8006419dd15f06fb1c6351d0f4aba5b29719bb5040d21d3cdb8ab0cc3bd7d8861f84b4fbb92a5b6c7772146a106468dae6b138c947961a8678dc4e1f41ae2330c5e5a20363039e83d0de42c0e79937c148fbeef77a8969e18d356834f6ce0ba08e273e419aed49d3772300238e6a61f99463c81318;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he755c84bfd60287fa123159c75b2f20966cc89b2f1c92598aae4c3ca3dcac280c9b16835b0bfc7614d2eb979f5ad0712a0897812313e0327a1144bd5be85da9c090f050494d18ad37bc375c73d212dc6e2fba135f69a30149ee97eb3d2931b478a5b9a1b1974e23cf74bc8b5a374b2eee8c56223ccd9f8142e9963471d180d7f2856953a5ce131ef7b4c3ed7f44cf23c599b253f27f7f456194c2ef0f76f01fc059a49d08dad18ea42ca39811fc981c2ef9ef0bdc8769310ba45bfc0576a9aaf9f589e1758d2c1bf1e747863db6a4fdbf89ac7c2e0241fbb036103e844ae00d549ce7647be56bf59c951f21522b89c99be325eba214280889e424a7b0e0304d0fd229c78e1201adebfb84b73fa9d61a15ff6f62e18a6688d8d5175f51431f1ca796317236b357dd4b6ff99c93c5e35650274d93ff6cbfc7428f09083b2f3bfeb51181d35e2f7b75f30b569e1b472ea07a4c698797dd69c10b39292946091eb9eaaae4c56d217866f9223b13ffddbe28dcfce08d0bf04556ba768a25b15e857f3c0e5f285d634b8216cd3596de821b052ae5db22377726334be5141bd450b81e2193e126976d02068032f3110d18a2f823d082664abe1d10831c4c318f98036b470e87aa066f67bbd72ea8e4bfddf022e657e56831ec7683e93d8c673fb040cf4fec52c633d8bf5e366baec041450c4f679c04ca16606ab777225b42a18fc52685888d2dda1b7f339c6581faf202a16d0ba3bbc975077a1bb6f4f06fa30bbf50a1ada9e55c3ebdc25ef2028552df406789e6b7496eab4facb2c5b719178a3cb46f53ef44b881cba74ab4ef1529005aa45947d31b16e2639474911892f69441a19d064c6ea56273c1f9247310088def4a8f4d330701624b2ca33b353cc61240501fe024112f94f6f65b537d0d589ced87b765ea6ac086277c99b39fe11fda86e4109a64addd276674ec931862183f7d6c7561c8fb36864b6eac53d848b9304630d541229cbc5d2ae357ad0410e0050ca3d72941632db3bc21e29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3a3ecea853b365238241cac81ac5d4a21c204e68b225e7f6292407a79ec2c77e536df2aca3be1d7a5b93f2c732ede4073fd5dc327dcb6d4bd7da595a30e32f01fe81b4d5a2d5c6e0c1884bc5410036c607e6777e8011ea4a354ae538f9e28bec4282fca7c258b436a7a5a1f96956aef6b0271e19808d4219c4d8ef83d0e31377dc45eab38b0f56f5e9d7c674d287fb8a67b1aad5a90e590d24fd8d87202a5b277ce21ea0e99afa23bdedb428a06a84ab25f663dd90b691f705373db30787e813bfa2c1ed37ec5b7a06a782b78b67c0b6e45468b64f6fa56dd219a5b309e41bdd44ba96159d460e00adcc7176eb5ef313aba022fdf757634efcb0562d3c7ae2409c72d55991a9c5710109559bc4e33afb4a0d6c7f59a250776e7501fba9204ea0ff6659904aef5312b3ef67830f2b62e4e5887afe36d2e673cf47cd57a1b641e4f116cf22a1f031a6c4c59e16e4675eec0c564cae61876392206a6c7741e84ba86700b6e7ebc796a968c237c582e6d6dadf98d9bc64113d1bfed9a297a94c0d6b5933d979d3bd36cf2414dcc518ecae71ac388a2b7512aad7b0c855fbbf8aba773a3c21a931a965f5f0b71f6303271ba92ca322fdad85f4a61a24a9747e3280b077dae7e3f0c6fc09f957a1acefb1f72142b84ae9dd06d4d5ae812e9fb89c294fc0668867cfcec8973c7a8336d892a7dcf627ca55b303ce61734bbee1053a1135e6a1f9b323c51d27ed67dc3d4b6faf4ec04c10a9e6b30930e01a5e2f051eba5370dbb72ff3477f74b565098d125233653592a18be480f23e26f7548aebcb4d3e8c0b779d0ed87d70cc3726690f52fa628f6d9794b1b027e2c4957fc2320d2517797b48ce784f8b931f4ad3ff53128b1ed4415174e23b1d7eb285d8149e45209b95e458a6a187638aa82f1287b10f30bd995412f05728d298009f8a2a37a5e68d9bb6fe42ac0315323d34296474f8147ad061ae016aa2f11b61864832ca8a302f49785cea1233f0f0a9e82ee67bb230a8048288809e307fbe15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2ed54ff31eed7f103c78b61839aa9e0a33f3c2c9bae43909f307fafda70eb4ebfe04a2da85df3b6fac07f3a545b45463442c3004a1fdd6e95cb4e9075c3f7e2bd62ce3a355d7b5bd654ecde36eef496f3547065245ab4064d2d6982dd964d439b76f739b52460f425ea4d0bbab88bf63def20a07145ab0af288595be4451570d5d3dd245f14941fbe00ea40d1f5493687fad4d684bd7d3fd9ff5473f7293f0dc4af3a267f8111c3c4e487b4912e23700a6984dc3db45d2a0489ce4f6c0cb4a47bbb7927acdefb693347bb9336bc8b4c6c43beb9e8420262119afac8b66084eab24da91476409d31fb19b9d1f3b245fb9878ad2c3ef5cd0f1ebb13868ddf3b385e144535739753abf7d5da35e0ce799aae7f76edd1ef3f729f5f4a04a3826811a95b9339f787c3087381091fa0b046966d849dd89fbd756fd901b32ec80dcf599c322cadfe6cf6bf73c935a90e1b937f09980d335389d3a3cff2acbf85797f0c2e1b86f8c8acccef651dfedd126e217f7f64a0424cca113350466a238b7819cebba4ab7788ce0f35e01c7e71f1b18cacdb4fb9b7af9f22708340366a8d36eb9a5c1daa8b500132072403b68c8e578903f26252c67887347014a960a85efc4740227dc0640372f0f47888969ef8f7562e19149ddaf7f8cf19f9bd7bd468c7a8fb734d91ef6f8c2cdb87bae8a2255c2e1285cbd7d8bd7c779282e885588c5c1f2e732809e08397158a5ad2cb21a54e726cfdc5fbbfc14d4156093c6f18c41b2bd687c5f595095ed9792149b9db24e1c74c7a4e57deda89caf8722925562c352ca1370b09cd6385413879dbe695789205f57f5ee6fb058d5d97374ad8b5b316b9c584b33eeae689d7c3e8dfbc44343d035732446b3d1541aa8913a6182366b9e1f4f7fd1e5e9d4dabf15957fdfd03bf147114e7044b64ee5d199bceb1db7156650216bbf4865b65d4cb353159e69787bc3946b6ad1095397667ec4270d12a614e6def741387bd90c834f3e92ac327db50da43ead49dee138e1ba96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h985796e14090ae52a29ef697cbae686b664c2a3b1a9351fb079139b2b699a96af0cd11531714f43b1d1c1b8d79a389f8751a1271c4e822ec054cbb5fa4c25779804cf19eeb903a7ba41492a02426ac9f0fd82976851c42e93c22b2857357909f549a19f6c5f80c8fedce53bcbfae6fd9b6837e6afd6f331b9e8cae6a3d579bea0db3ad0b5e12694d1edaf99dcc3c5b2b29205e12bc1ea34c3ac581d3c6546134fa543c6a0d2a35c6c93e521eb596609796105a1667046d3502eddf7f7227a3990e4dbb7798fbab10735a2f6d814433486f8cef53d56975a26f4b78b74a847117cd3b75ef8f30cf237b8cb54a71d12439c80b0a61161fda42f95387ffa4012b37a8f0e68a80ebaa19513d29d9ba1f6e02d316ceca66de0bd3d6e600177beb345da18af93a81e1652c327d0400802ea60249ceb4f3028d97dc941f48bdf80cd83405013f2b9c3f817b3dbf532df99cf683945d73259a007b4fe5baf35407afc1d96e74e7deed8a391f11a4b18efed8fb131de0667f48b29f58def02154e22a7e1ce707ff0f961d7f58b7fe89b91bef4a1b4ef6d76836cb4dfeccc30503401417448ffccfb7cff239a1371b9e49a7b5ea89a6fe675cbf71630987df333e8a806583b05c4a2235e7ba7a5f3e56cee3886b391f5b88a1a6c09aa1ad3ee1e20cae3d22ebb70ba7e69c9bac1cb2d60faf5eb8bfd8f53fd9301b5ddfdf7b741ca5c1d0ef880c97be46892fb2e451f6d2eec2c4de86513141875c470c9c339fa10cb2c3a624b5564b61b7cbf6a7d44fc441ed3914fa255b3e76f1e9c13d68ca74ac536f58aed65a78b0c360db5b89c5d97cd8bb800f3ce2e4dcf9cdbb525f2468748537c8bd34cd1bfb952abd886f0cd6a725fc7dd99b6c004305e1cecb143ac3e7610ad87a770c0c2374c78bceeaff50bcfcc7c3cdc1b2d9ca99cd5b023c189173973b11880a473f97e9744358b539bf55fa0eff488186e4630a467266f2196a96fad1077be6be17d7e9f960254b50bef48c8c066891d9f7602daa542b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h97d25b31ea940a0ff3166c2f661b1016738665838de01dd63afa8a6aab6b7213d6be3f9535b3feb521f944dba8c1839f68f71909e869958b99ba1887bbe2450cc2f4a17d8cac23b9d74a44cdd694d6fb4af6319730e4c5f1cb37fca02be6c247648552089ebed66c03770d1fc6e0efe9d47a0ecf0fe0c2eebfa70b5ab06247f45b01f901188f51105713dc5f4d9fe6b33edf109ce09d789c05b4ac4aa9cc76ee0d6234cd73b8734cd094dbeaf915758a109a13aa951099f3114e3ea43c4cf2438e9f47dea6f85a31c7071029b233a3df0f6158981a3ebd491cc4957a704bead921f5d42d4dd767018398f0b2ed397acfc96f22b6a3abff94539a87381ef58edf0f9763a551d22bdaf601e1c73eaaaefb3c184a51a8f87661c6a61a46a94a6f235ee8df65d6f51810c0b3541648972324cbf3fb817152c83959ff24d739ad3aa9a76c358a67849ea3d90c891d880705ebaf203584af43668694368af2773836487e57846a9a7b9429e6beadafd2dabb9186d4f3a3618c0175f84172fc752e4a3aed18511eb53f0a8fe6b1f27a199846fa5a464897bdded342517fac0edd34c0e0623bee130d25094442e047943d54021f563dcfd08cb7d5444969e3be45dd5305d5bd4a645a6e6a5585581643bd6f148bf16ea6b37ab10fd3a715c7c7cb2ecb25097edd2a5cb1b01e8bb551ea84f8c560c3412486d1eb4dae41737c804b32765c1081429de157bda9a2793a33f8d84c26ba716aab2607c0451b15e3d4e8191831983e5a3cd720156cdde7f4d7595cf7850594a87341666683d1ffba59aec6904746ddf876e27dfe65d5e6c3d928c8a804997183e37234c337e11aa40d2d16ae38eef85c1dbb35dbe3cc2676218b7a70ebdeeeb8175e192adad698a2531b50f72c292f8f984870926bb5a9997ffdb7d6f81da32cd661d2ee2339531c3f7ae8a59f7f93101f8dc0a542ea766ce0aee3651b592892511fa67fc258f5ded942bb612d323d25d540b91d5b9886fe8c6bf2888097b2d807a647a45d99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4db9e0e052a02ba06598c2aa98becf5b77c3ffaf6ac65782b21640501374bc450b58364694f1ed5bd20fabf364c8c0d144c1f3b3c391b7f74212d38d2845db05a63760a3078b1cd8cd66d0d461a648163f21bdec7e7d218604d40e1c6b36c8293b785026252e05b575bb147eef797745a55876bd60b9bcefa87c8c65f44aadce8a0eeab36e59a2d80bd9d74c68294f581233240a3bf4b5ad9ceac1b025e1f0543fb960c20b129d66cd0409bd899ea7acb9a1f0f6ea114e5f82603821fbc7443ca594d02fa3b9252c193e4c2f46a3bed663518c9d9453580ffb37963182a329d5ed933a5e614b8494e4d4d698700e9f93f335377faf381b3d6c89fae4ac9c7e535f869d6d8cf04d4575210769428de4249b4452deb6ffd9ca58cc72e415297e204830415cedb3f57bb43488981a807174411b50efe1dd871c9d66743ce49963dfe9562487b363f10a0a295c5c0c6633e37183142391137d05ba905dea609e2d17e468f33e4a12ab73aa165f8d15bd677de4c2dc0ca6fcb837a9e97a582fa1684a2dd9b9f6b0746bfcbaac1c2fe9f4c8175ef0fc01e37fee6a03ab65562ce7d537d1716c221595c5cfed13d964a257928be16f61db6a7b8e72d01b68624a867fe6647c200d51a96f83c2d788caf7214204b020dba0499d0a0e09207f71ad13021575c754ee66d828e3587ee30047a64e5dc892aa0b39991aab129a2c364bf7b440f4e5fe72fd6a15f1dd2b1fadb545be5afc48915c64f5355396b75cc582972c8d882c216e1d51430d123e00f98044d5842708421df2137f572bc5e074be1309d44d87fdc6441c532c6e7fe38f31ba5c83fe83594da120a9892e0bebf751bdad90a615431f8716e4ce881de20855859371cc105fedc6cbf56f4e9c8eb1335b8a7bf46ee2a5a8f856083ba17ce187cd7a125e3d207772821935ea5bdb8489e132432282229072980765ed23d0697d58c4b3994b6abc8a4a5647fb70abddaa34460196521aee6af618de8aab0519df2864e4d039555bbe28a16249;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfd4f4eba936e5ae506fa68c21902a58235d82508250c6307b49d793a58d0bc6d86d2b80aece12c85e31ebfc21754cc0cd62bce0e8759a26a5d887619e02e1aa49cdfc357203ed1dfa99c128aecbdba2dbaa9e6e1dead1d5bae5dfde9baa887e6d05dc2d56bdf609138919758308fa01082802693b7a6cca6744a5ad06113e15610a9a535e9d9b18197c7ce81600b2a915b50c775bde55e32e3b95ab2a7529de6b03cbb0e4cde2caa9e39da537c0644e233400d7d0da3f0505250ccbe0233da5a91c61ce23f868cf46435ac1e22e86d60ac3466c63fabc0b36c74f22e3510d457a50703c30a36d72dad108fef3d6660130b215b424d95045bc6d686e6d42980b5956ecdce62182ede3987cbdae59edb557213275f853769d4fc19bf9fc5de067df320c1cbb2182baae5aa16b62dc549a91c919f0f6136c9bb844e75a9107d52632cb7cc4dbe8e3bfbe907721b4f367942bee6edd52a363dcfbdf40144dabd3d3f5ecc0dd907764d92fd878d567bcc67b374c0e1c34611c3e3f4801927ec9419ab9284df71f277b2efc33b4b5b4646ba73c0f92cf43700903dbdc3988276ce14263370eb03343cc139dfaa321486c4975c96d62887f7473fe704f2f3ec6b206ce15b2da3586dabccd9c3dd188b96fa550d374eed7f0be6d0cc2285c09ec596ee6ee5b806abbc4b372c2282e8ca6556a54d6028106b6e005c7e679844eac59457dd90b8d28bf564c2b89b24d91ecbdcb72d3e02cac55d5237980362bf3aea9ce50dd7737bb7fd9eece50d30f955fbdba2d17e73ef30d2e667e174336d5daa7f1f22cc361a1898d86c3cb8827695d1b374cd4e3619265f2e2b472a0b6feebbc563d870bae4cdcf176f04f0b3d1c2d5ef70eb12d97e92775d6c42a1f7872653c2595f6a4da02fc4a7cf923e190c021532e43674639d2c06d616a5dbaddff17b7b0aff20aaac48413bb8b3284f160fb3ac040c4f39c0fecfb516f3f65be1604a35838655b3fd8be6072debec218781f3c497ba677550e8d300684b2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1d14d3c159f8fd5aa2197cf11540223dab9c5bc794b13be0a146a9bc3c861ab01c8625d12fe7f24a09948ae296912ee824584bad637f0c908128da4778ada5ddd62aab7eb3deb9850e9591494fdb3887c93d2c47d57f9279788320fdfcb507028d31eb5eed032620f4dc0b2016fa2a8b1057fda53e66622c0945974bc17c6b4f6d5eab61bc45708d8efec1ec5aa46f24f07828446b4d5c3b69565b6f1abf9558b6f6de44defe123b10eb2c7e7281406ede4dc1b0d71c07a53f3ac32da7d7997a4453ef20c1aa49900cf5c2a3083dd174fef4fed53b2ed0b1622233a43524f64586744b4e70e2d1cf991e6e2edb8642360d3e9c7d950a503136926a121e2951c7f24e3f1de64ddcde146dd35069ff5fe878122582f840ab6b298c2857051d7a6ec087cc3f5b770511329564c1aa03d7bb09ad025ba50d34cc1ca45a140ab8ef41626d05cc591b1bce6374bfa609e1a4b649ce51affe97532ad52eacf80eaca93002da6f47beb5b5d03c6bb09630edc25e295feae3a06116c2f6c29c88004f8df64d37b8be1af8b6d4f3c9662d99796afc88df727e6fcea31b7f312e7eefbce0971b631571887c483b4ab328959012abec86bc62da70c5b562868ffa17e282ad51025b1285e26a3ca6d933963d364b18e470dc0472c109d20e7a44bd2dc69781ffb1dad301b16458c327060de886bbfd399318ccacc2d95cf5d30efc0e2f261096fca3f136dbc4bc2f9bf0cf8051df89d1a005b739c6c40cc854f74a517a4ed4c4f06881fb32586daab78cb121debfa00e153ad31290a269b8b1223133b6197172c8c0fdab45da084cc117be6451084d9b8eec6710d7a62913b8864e42820ba86f26417d0d6963cf2a030bdef14e87d44ffbf14ca37c38b129e96b05032c9b1d0a12b8c19b64b6cd5633b9e91a4125e14cdec75b1d1e310cb6ecbd818a52a178c74cfd1d37c922838cf598b5015bdb6708cd165ec35454bfe62b6343243b6c2b8c82394d36a64237ba66990eb04eea883e727a8409023c3a065a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h338311ca9ac9f6cc82363f449a05e57d1fbc1a474327dfeec00a4804d64831dcd86d1534f182fd6056a19c9a84b7f49e285c3bb9b12ae7ca29c1e6981651bab8cb5a42477ae52869948f4ae2dc3fd13978568c94469e8991b954020aa3ad660923aa61afa4a138deaa3316a58f4d373e9233b7652cd25a638aa44eee14120360e122a99a1682591d271c006178fad16bf2bc30e7dadda7fba2b41e5835a02f9b449470598350c63a364c1e99db1edad5cc5f92eacbe746e28fe195ba1de951815a0f8b7d5f4e2490135caa5eda7c4450e4260a4024f0b9f9d04f99ecb5999cc891a3996be92d0c379af1dd10fe445c7b206bb01b1123a2b81b018ee9862e7ff832ce41cc2889f802f3129fe63c4ef29624a8411e72618a771b0a3c75bb4ef08d2d7333ab1407080ef9d480a189b269ad3a48d1818370a4070716299bd3db23b84bb5d0681c138fb34be451434124636b9e2f66ef74232068718209700f6fd7ae65722e75aadf3200e80c5986011156fbe1ed829ff9292dc25a2302e06b4b48ed1e60b9fa018121ef2be939fb47ab67c5780b58b7c9e0b32015c6765934f5f5914166a2eac20d166830fe7b2a684f854f3accb654d09d05f405b7806414821be198f50f3a04758b95a90dcd2ad48dd126b647f8db645aca789c8b6c09b5b7159a879f9228d4a1d882200f8f884e4bbfc0fab35ba410fa861724a7514cb78a39d9556a62cf4a8200b8c6eb3b06f698db9d165109a7b5a3bbbe0927e353cc9be1bfb65102171040fe99f242b96205ee19b8af61ade0e3ae86d177ce7dfa35e0a59cf10e78f08a7edb6b5b0298e44237db2ebff3453980d5d1c2e1f21cf7a411b727e041557fb59424e861ab86e52d280c5a6e043882342572925a70ea5339a7c6f67737929788b19bfd64c0ef1d055d7ccde0c611873b51e9ffcfb944461ab4a0ab3e0f2dbb9d5ed645e283add4ab2dafb90e2ae13590ea7877442726bdf6ecae54655a84070a1a02265edf0b4386391aeeac17f02307ad4f0850;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he2986468d06ac48dace4da5f5ec4e0ed761fea6a5f91ae66df26ea8813a7fb4ded3464763ec259abda09a6aa1bceb5199725eb124d0ee00212135fa9663d5890ca95646ca528b2c2046d19e62ad1d8ace3b84293d0bcce899134565c280cc58a9ac33ca170abe968275dfcd0d4ca57c1d0086962bf5b6212b87f213107145858e5d6c053a9f6e8f8984feaa8f980b56d6e793fc7141c965e2c2921302f788a5e2539c44a9dbb15bc1a408b48109ba1b35a731a3333f08b33a7b309a2174ff773b18a9d1a09ceb621e98633f1c4d8a73bc703f5e2d72e8b9c2664849e6d9de434927cb0aaba2f8dc2aec8770fb056dd99535a7ef100075d6fe09b19c145a1d072047af0e965b55b4ef9e049d0efc470a04ca8e51be4a5fa8ad5ccd95c9c3e38222da13dbe8409de8c88d5cd86e15bb54546acef35937459af7cab67c3df114ba4fa76dfa0d2cace8c1c998f03941de85059774f9ecba14d3ea26e5db4dd5951556ac99f450e55aed5bfb8afcb121bdd3b2ecced2789213c8858078d8298c67c639418d466df68bdbcc817ba47532426c7f1c7e1c463b450fee57441c9189bef4e0bccefc70016b0ff00496f655aa3902bc7a4ea12936ff79fa31fdf66ef0aa01ad3fbb67406044fa04f7fe8161d60d2371d7cc1da7fe8be61ac6d5fd79891e9ec86c4ae695bc277b9d5f19069328154856d36eedbf12430d45285ccc94803a970aab38ba1173e516f45f8cdb8931918ab030e9e66a2dcc96bdc983fb606cb07b47c99430cd6d3401f453cbe32efa5794752bf0e44c707bff671109cd7e13e3af6be180a3f002d561861f1d0eb3f60047eba12ec5e7207e622a760d759e36f999b45c4b32232f7d8d8c3135474efbdfe8adeef8ea46c80eea2e19e3d3c8536c3df69449caf3060ce729245c68ea9dd69bd33e6b5e5d41d7c8a6dd57e8a560a022fe14a41de4b665ceb09bf5b3ae6672db1355f257062b68df4afcecaadcc12c1d9e16a4ea1064aa74daa7db8716031b2be7dd8039c01b2555454;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfd3d6e7c6cb8e47885bac9c42655c7f2db87f1b003f626e66bcdf900665d45dfd9d313bd686ccd7405d0406b1236ee05fbb17eec755c1740f0679883c096cddc2a60b5698927c0c633530f088e04ed7bdc6bc67732a792146b7eb2b5698bc3a247cd9212fbf9f536a9195714e12c7fcf7953e95da87dbda0dbde744515f3ba6dc2c8a0fad93fb95c17a06339abc6f630a47481aa5a0fe91e5e2596d5afc3824c867d096490595f4f3b46a2b49d73394327bbcc585467103c1403a14190834359731edc5ae946c1e86fa28703ccdaa83687007ee653a10d99d524b8df0fc5faf56b4cd83f451b2916581e8ac19d5c669ff803cc51a26870e632a9113aba768936a128f6cf6d5972046ca82d8ce18b1251109c22c9f1366e2b41352b5bef20f12e79d842c7fcadf2fa2d7a7435b9c9e769853a0e2322bee70d3494308ced430d5c95c998ef383a64811a35b907454017a3548efbf2e60016d26ebea44936439ac17b548ca7baf1c7e211c5b4d15f954f93a34f1eb0cd32a449878686f2ec7e2bf800c1ad5b0f74b4c26c536ee1ee094ac38241809e60fc10b69f9f1f18126721504c7b2b72a732e541ce4a42434d21275e8fe5ad363ae2071a5184f9345aee23bdb1619af0966a922a5a8ea127fcdeee7ba807b57e919b47736c9e1300edba571919ccc05c9bee300181c77cef5c7de53516270a3dd04a2db883d5fa42fb435d88284fc0a27034ff54d4981f88c55405c395ece3c264493572f8ee0f234668d178f1b2bb846844eb328e8518141929a246e20fd2cbd05a0441feecea35ecc4f673a4bc0843dcb3b5fcaf3e6d486457bf18d14828f4685fe98407c09af9961e7b6cc7b6e68ce7407daaf9a3048f72ad82bfa0a6717db398f4bc06fa0956133db9ea56bedbf3aec6b82dc0e54bfacf93963e33e560317e81e6f2dcf168107affa5c9480994cb9777dc6e86574d0c9908039ce2a5d18989a853d782b1f7a57178ac32fd9c7358d953d6796a7ac91549c5cf03059963ff8f76193f11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he6e891cfff59ed72c530a666c95715688421faacf8a880e01baae4ea968daeccb16d76ee5ea36b16e3eb9bdc1c5656772688e6187b382c02a80e28f1abbc67b470d7f0d4c5159d5623f347f7f97b478ec8e4e00de8e246fb757563685427ecbb3937534c0377469bda4518b86425f67d996777d9294de0896aab012454ef8a84dd802d096bc7220b159f648909d88a6ca5b0902588aad6471b652f8eb59d22fca86da5f6b37a3d352793e352c25a70c18ab61361e1e7d022b2cea5ffeaf33b539ef0d73a268f41807367e113307c3c116e0e2f9b277447f6b5bda45a209c47064143034e350a0b8578e0273a069751502b50d7919f9205d47a69a057b2247180434ffc9930cfbcbe47b1b7be21402809615ad2f3567625144e085ac13b0e271824fc64606d1d2055f76bdd6c523f354030ce96bcbcd4e7df4429765a079dd4736c06388bcbaf12a64db6649817decaa6cbdc36a3ff3dfa8c79fcf0799f6f43caf741c847dac976853f245a02c6655996d77ddfa1051321f45ac159ffe819071aa03c22db10d517d0772536272bec23cddf25dc761a7a2a400cad926535796ddb5e9a1b0c66c06f277bbae06db9dff30927d40975d82c339ce7bd8f73735ef469e8b01f54d0face9a1e37bf1fe10b188110602ce27cf4b50fb154ef5965255cb8d0ed324a0e61fe3cac8fcb7302ce47711c8255eb60d618ce3ce4a6b96794fe6aee7c1f3dc322c6b3075c4dd676a402a41b2ae6e734c4f8a4e9d76f84bd5466f8893f0f10f324d0fecedabb1a85c33ca687e561f8efe22ccab50ad63d721b7dc2367b053dea7b998cba6c7c06e5b88d45dff9ec27b02fdcfc241ca998e181b70a94694a1ee18c870f31920528acebadf46dbf3f574ad922def630633a2621a71fc56f702b4899db93de10d587eaddc3f73074cbfa7f101446ff8491fc4a885cd99bf5e9175a940b88d6183461c193d1af946b3f9fa409520db91324418929932bad9a7e3ab49b5f9d5d53efb8bfc396c271f7498ef350f0576;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha8dc208ff98ff6612608b0fd8900167a7b2fd69594fb8966b6599bdc24716ca45c10ba852893518c09ad74db5325b4598d06b2df32786db26f95981c0005fbee589a93d3aa83c6ffba39b441298132b27821aa7d737b838cea10a7e014fcbc42a42a9f21fb0d4b0d74b91e0a7ef3e1808d20a6512957ae1fe860f4371e810ac2b7a5fa5324bdc45867ab8dff064f090671034328cc74598b011c9828083dfda031fce69b77258593afba3484cadd636500afe614a59fb6d923278472d5d07ff551c604cccaffce91e77b7601f58795419d2b612082b9d1b331498d7d621573a1bbbcfc4863284595ea3a6882b5c842b0e635f158ccbee88efb6c6f776e4dbd2cb9f64c62a4bfcac1df05e64a273ee913544f456bb4ea5529bb53599af1ceef1cea6c9815b47a5f8db678bedd77d31c08a235c08b72766e07a3be10446ad862da6f2f2c434851a0a2af45073a91b889a33ed69b0306066219a108af699a2f943a99db92a7cf816b9b2cf8f57f183691293700a74595abe59f1754b220c3573da5dbbbe1d97419edb00fa7fc0b6c21c1eb82081a7d7cb7a985b8a7254ee9992b892e8dc06aa4aedaad9ac512b7f20674eabe8d8906dee7197455d31a4de4ff8d34020eca5363ea7ae733b4978e6a24b8fd0b57b32c229592dd46028566b88f9890f3e0346afeabc263e922b2961e7e3e5233c8969defd5c291f1fbc8197e4aed46c8e1795a694134ce873719d404dc07dd6e8e79576e9296b080d843734febee145d321929ef436f329106ec43b38971fbeb6e8f7ff043f6f8b78f6c4c2108c4a589aafaa01721fe40175f8aefb2153360a4a69bac5fb869aaac2e9a35c443988ebb49a0a54427f51eba30f35f0cf18c60bfdacf3f6f51e3180765e563a99ac0088a92a7ab498514ffd337a87f018e4d8b1353a28b4669492f1b1ae623eb9be896fc45f6e09b6dc4c89b7e3224a5f9ece366186e3fa263c9c070cb8d2639305a892dabbf8b80b38b8cef6f0cd8fe23becc2c5bf5d0e2269a3598;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h67981d4e8340f99834e6b1c40f71f801f5049af8ad1ae20e60458660918d5536f040ef42c4004949d23bf9f494a89a869b1c9bbf672289b89a16e6a68c4b1d88202566c0ff63d99f75d2e4f6a860ff169dd2f1795bf7ad0bf88f15a8d9b756106f566d7902f6ba1b71d39fa9ef986821c67fd3475bde5f1d264a2f44caf2ff66f7c58dd3867306d043e4e5a104696400fdff91830b563a9aa420e44a00f25ee47dee3dcd622bcd848fda6c56b9a17ab8acd6895e79381829792a0508ed316f89e42c7306646b44d52f446dad4329ee8b7ef5efd145139c74619c3a9ddb8559911a4e5dde8417e45fe3b5052dabf8bb26be0531b34f1290fd164b92c3afc8be08ecd279ac759adbf5d8f3eb071fb81f30e51ddaa87c16a5cf64abab20fb0e34fccc8355c573f58dbed54dbc3af2dcd136c82be66eafb68ddb99899bb2f25a92675f4d7d1d0d01a0472848411473d135373b095f57c348a671ecb21b96efb5b512a832f10bde2810166b29e6d6a89d58a99e68eb3038587a2be74c6f6b0b50ca964785b3c9ba09d3c50b2337745aa3bc764d33a1d33631858a074018bcce78a1e2a8fabff20c4b2cae60ca363e7219e03c5fb81b835b04308fa139be42c36aa7845f7702635092eca427cd2c970e2ce7826a55f065b0dc3a8deee59325108ae65926c1c7a8f81d2c292a37d4436cf091a240d0ca77288c00535dc1100fd6d5823c318c69ec1d3b94e42bc2819b2d490b2b88c1690b246869439bd7e5b5be1cd4dbc2bcb9ffa58f1455ecb2c942a8b9ad3d6aac06b2ecf67ce0a51610046a308d3e213cbd01cfe612400b4c52123e22e7e5caf45bc459a308084bca685f3f04c4d617aff9662a05992a5ef8137b75281cfcdc393798803d1c3c2b640cc8454ac3c172490cfd19825dc7f75ba6b67c0d2168ddf50d141489f50968f40d9bccba688c333f1f902dee68e9651cb21a1d13b97d49ab7c489ec518ca0cbeb548cc6c44cfda610407b9bae69bb1910a35032117f2083f346a406bd4441e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h382244deb4d3dbea28e8a3b6ffc8f4953831450533ded8eaf40bc857fc0955be5425aaf8b09f9179e186f737bd305473252c2a0e87666033ba5fb7d52e4ee50e305308c9f26215d96f04a0a200632b40e2deab0bc828fa4d0f4f97d6092271be7f5932f75ed307083b4ea4d2a0e08cff2a7f26f7f23c2fbe363d44940801b92f2facd61e92c101b53fc8f2efcfc7b62aca59335f5c813b46ae8ded857ef73da5feeae1df6eb661da196f781f0e6cbf867a2800d9a13b945e4184e981fc625764d44f41a9c2adbbd39cb3dbb2d3b8159e3baf62139567e73b5e73de071326222c84357f5e3deea0d100ada103af1f22b74cb281f337c2eeb84a0b8eec6174ba1533df7bc1f96334286b3be1882c36019fb63e565a5ddcd5d3fe06d1fdec83e9bda14b6256ab3e519b4bcfc9f41748a216d576c9f2373a9e105101d4e3879c7eb5ea9f2310b567e4269266f2a7c98ef57faa6f2d02f189f959c973fed658f0039779291c203d7a5139386fd98826ef05b5cabeb8225641130a9a6ce0827eecf238ca3d12d944587358cd9ebb1e48456e8eaf20cccc347cae6600ba58646674e5e651295320de1a69c0304dac6be80b4c75d83f85489df4698d1b8cfbfbb8cbc11633d4de3b73acd01d20365dd9dd1dbe83fb5cc0ba38134931412e9ba265e29831a79c55c22522879a0cbdd3220c64ac2b4a5e4157a3f67806dc21bbc14eef6f6fbd97296f34e031bc288ca50ea29b1aef0c053fa00dce80e01c7184a68352e3367abb148aa7ac1042962021aa5c55d3bf9ce0bdba4189cbfcef8be419afd37c255ff6627d6a1a6e76f1539cf6ff09203a15480c9bc9be5baea4dd2c7253485b0bab10d852c5a93dcaf776bae9b1fa60d0ad4988146aa4ada2a0524f0d1de2b13aa536f352d889cb8fecf12170e32fec2804688f5a4e836417887610dd69fadbfa62951b3de6e7a75977a31372a5c4bb17aa51d8fcfdab285ccfc91021317da6f537762310adfb37fc9f11d9bfacc668ee10ea96241b6d7b69c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h66ad54819133ed238b3e8aa0c93023a0b9720338ccb7d59894f43ac7c0ec0b412757ea5cfa89a509b42ad09bfcd76eadae05cbf33fe02beda0b0863452b1fd1eee429d1e02e854614cc9166ae5215fb4673141ac49e82c642df5f350c37932cfd2df6b7a27dbd0deef34849a985dfab239c0f491b80745ee2c9d3fcec6173a1600e2f6feaa077a0c9d7b792de18846da8c51030d08da06adb7aad05e44349bc3b23977aeb57d7d4a19cfcd70e2d5e0102d33700f40cf8f5d1734690bd84e6d1222a984e06efb972815844c9d6340b8ae367bc046666874af8d790de2f12bd5097d97653d6304ce48819d27efe0739dfd3deacb4fb9b81807326276b830b493b00087ed6e4fce29c157e4d172d10ca44105e920e32819d948507e80e9572d41ccc0e6e712bb70963888ebe43d26e9e9473cfad4be3dead6178798a1b6a822053966b7c2bb217cf1c78b872d40068122be5e26708eeb3ad6083cfcc5198eca6d2e4711f03cc97cdce28bc756f9125402f5175b8d4b197ffbc85f78a791cbd343cbb9d8025c3f21729eff5b437cc08231211e6c25245848bb631ae6b855bd7e78801b08102691bef5c9389e2a02d257564fda2d9a91d4519de7b0dfefe5de50dcec6ec5efa13fb5219d29bf6d50b7aaad6ded62f16a3f220611ccce22f4d479b045802292770c8ae6badb4638822de01c9fdba9edd5840f679e58810c9106b5d6683497bc2932f722d6cc12ea3ba05dae299eefed751744451fd71cb8483a75eda9d9086d4e4faa88997d29b8a6e4f739f3f9c721b6bbed389cc2ee2c613ce7fcde130daede91fc497bcd30055081ae22483fac278c36f5eb9a54d1c1f0690cc8b58e19302386a34164f484645be7981810646e21699ce9abf3d8bb85f00391654200055d09078bb9320a9f3f1c7ef915a2ac0d2b1474a3fd9ae6f802ada3fcd3ed66cd4ae31db66e7907a1b9f373c34f5e0aaf1f54cabd635831d839f6d750220b7a4a50585dfed19e8dcd784be1077f9299c91ed7b7719c6f3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7afc743ea7250c1b79a60fa8a659dd4b41fa2a55ab010423895b1f2fde29a1b31aaf38b9be43a13d8c5fa28958c7f04d42a2e842d7d39ccfa20c6a38daea84d4c254b107ff80d47886f08d118d6da7a5a822b0849e648165643ed68cbd8338ffcc6a178fcdd6a5b9c4114908f78ef6354b47e304a503256575392d2bb562482f9cafa89016c6443bc527f157840cdeab7720d32b05b022f2e6db7ff9bdebc39e79c5ac6047c75e6422584f243561eec98354df7ce1aad6c693eb42a79093a6e81b48820c058e12b5b2ed7ce57659565430abbc13a5aeeb52caa04f0a09419b92bf5b42c3625f821ca996cf046839096e198e3da0d23999f3f274560fb3451b1ff0daa53d9fba33c16010e367b58775377117836581d1998026f33bec44c8d9d189a07c0f557c7be12efe815ed54a92cdc06f94bb17068961563787be79e7007e26ad1b23fdb75a599a6f3ef905506ff2c16b1ed857d900f91adb4b45c657e612e1097949bee6c74d92eb87b6cc418cf1204c748d6c57f969fee10e4a0e3c626480cff023a2f4faef8f33e34bb08a760dadddf7baf104e2f0bb812a8329fbd7f1020cb2c2850204ddbf2df9410e7d0388b9a62a7d11aa699fe02a65740f2c129743c158bd0d685e61e95bace93fa11d30f6b3f3cc73c9518e76830b9ba93c168a253607c5cbd7b768a9e5a76ae5322d1e4a842a90de818c9032cb674d3c53239feb000620461b0ee526a3fd8e925c7b1a77c769d35b1742213e5dbc1558d0e19f0c7c33ccf3dae9c1ac6dc8b03513654040a4f6fc06d1b2a79fbaf524843ef602b500e642ff62ff105423b4ce77958ea84d81d1c56c843d2114dc8a78fc50a0112a8c0c7f6c74ea99bd43021075260f57eb9068fb2187944242952016dc7c7794b3536a0bfad26df4a6dcbe83c53229a892bc9bb1ae838e8c8eada0f595176036e1a1e796cb6c979d58651adfc71e1dcb028a9a83bf7dcc0cbae72f96acb739332202fe333652d05b75e8de4184988f808ce8a5336311e4a9f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1a75b51b40572ae6d26b3d310d9616db8c7d240c15733f0b8a7be7f367e561c90131ed820293490320c800054ebc105dc6f66e84ba833d827a3f90f2cbab18b04b57cd2b460b611889153c6d157d65a90053be02fae4b7aaba5cda1fbbf4f298b8ef25bedbe5266abaa03cbb464d4ca4b9dce1dc4323335348dc4536e856ee010abba767d32b673168d4507832850c9ee5403a003f284d29b79bdad21ee09d15be86d7ccc9bcd5526c4d0176d0cab93ef6d7612f5070910cc7f606da7d844e00466a135e49dc20bf310e62fd0cf21c1a3e94084c85320bb8c93610d233f847da339850a8d463adfd0d205d2b55010d1e236422bd506f85673e73131c050065c7a9701f8cb6b88da364d65a93b7fa6048d1f4e5f849e0d02b0a3871ed31506df956020195034dde863bd857b91baf40f7a0ec8d95e5d73da915cf2882b692203f5c1e053cd3cb0c0d8128ab76cb8ca0f847764505d811d9939e911f74980ed668da871cb89a984e9b8b8bed6cf3a04feccf4c22b9c1bf010fbcf4ff322854cc112ca8fd6a7497c1d1088c4b5dae4dfcd17c74ecfe4ef54c805e3f362685b3e1547f11fc9d4369dcc060ba3e438e82774c5d2b18b5ddfbf9bb732e87de20a8112c9255c45b9dda9a363909cd8c7e3e8ada6864439a79652a690048edc73e92fd05479308408ace08e30a804c56c3f103a7f80a5800744a03980b2d281428c2f13dcbfb7340ad148e69dcb398fba79cc956da616635268b4395733a0d19bd7c247d59d627e696a82fd1997611267baa8e26cc596bacd7bbcb1cc18c8167398fef0faa742c5e026c27ae69ff241053ea498c78756e8cc085464f386549ce399d4f728cb62d2bd25ba5b029bf7cadad7b5b3b5af0ad6facb90056326680108411e2b901675daaebc67f4e01bcdeca92a318e2f18f9000d869a54d88e10d84e6269cf81df713d549af84131467960f071de77f135318f3f8ee54c8ecbb1ce7e3036091d85bb4e75dfec18723be8b4a22c2e0b49141f24390cf65e372;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd8b661b4766136e78d4f7494650deb7836cac44b75b84b671863906c111b33c1eeb1afa44a49e239f1995dc79b9b1b14a950c0d1267733960de3820ab8f8f3e6cbdf5ae62da1fed42233b3de507397ad8c729e33678f19fc3ca29c96591486e5b092da50ceed2b1974aa75225848ad0afc2c1b8c4c97e9be34c27aa89a97b4ded64214f8efc5ca7426483bc2ab59b3a193f653c6945ad3b4d3ed6a4bd06c9ff5718ae0dc47ffde5a3c84881d35b4463b98dfb0981f0cbdea41360e145ffdd6af18997e8d870185d3bad556987df1fdb6e0b7d59115e4aa9f32a02590d235492e9ac75789adf5ab57146b7478aa232f13e6d0201af79c720fdab217f2aee47e59f0e59ef0b9130a4b949ff4984c1f0be6db9c3a9c305d6d1d3266d485c5e74c8effba6b23b39ace2ae2489cac34ef7e55797cc4bd3581798688c733f03063b82c44659ace32844fa829462db2e311e28156aaf3833cde30dc1fe9307d257dbb0abdacc0029ed45c81c9dd55e674f3eea3e75aeec4b5a025fb7b1d5d654fe31c3be6fb900ca74fda82e9a68db37cf0ded3921124b36cd16f074b46360b336c1511338fad83efc18f1360d8dd3aed579c2c96e6b98efdcfa6d77b32c181642e5228fae9e65b3c9be882b964962e204bc011c7475a89e3cdf995c4641d72e0c97ca6213dac5fcf88193661497fb36b049f013cf3431ad90da1cc4c064b5a4c709f7dd98a88b4c1fc549f9489e5a485b4bdf290f053db5c68a496b340f6d740ab057b653d038a21a910a232b571f52e617ff54086cad468e7123ebbeabf0dafa58d707bc60c76183a870279d303d38bb2f74c8ffc09f23ed89f2ffc184f1464dd606b5d4f7453723872144c48f028449094d715c9ea31e00a4bf6b5beb45195d6718ab5b2ee856001637b7f85bdb3b703dc3404ec3de4e41ab12e7137ac46493ac74b066cb2d29b3fad555709b16d5a24ade516fc8e143946a59d02deaa7b70b33ef994ad4731247afc8b39af6eb8bec6fa8abe46432b41f13a1091;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha7d92c96b4021d7d774d699c0cf30379f47cda7aff0398bb0c14effc825f8b491b32a091beb7a7e8b1be0dcebe4422de4b3b14a739865585e63d3c72e1d928086f8651db7e2b47e63bcdb8c4bda82f4cfe81b5e82e66c131a50639d0e0fe0a7b51abaf78c39fc91940bddb80a8d2b04d136f6875c133aaad6ae6ccb6cadd35306623e187f19ce88d1f98c4228a388fcec4b75242713c346052625f52e52e4174ec7d1ed115d05cd71efbe1743c7ed7c12a3f071a13eb599ec3ffd2a19047943873ebd069cefb4766555215f62e5e29dfc24820a7a076b7cc27f3bcf96925766eebf54655bfcfe27d140b5590a2678b2ba7cf27cf06aa578b60869642425a81d36754b765f93894bd9f281311036b6b4023a08a133d4b4d5e5ba8da2dfe45520fd91b85186fbf42c737e73cc6af8e941a524606d1dbeaa3df41d5ebefbc73d86f515578513305a272e58c6ffeadf473d4fd4e0786d79c2a88f2027829508fd01aa0902afdd54d594f132e9015a493ad7459af4baae98add579ad26ad5117ce43cbf90dc7beb21c674695dd0f85659a5c74d8f353c0ad28976ab3942fab6a8c53662e71225f25345890b1d111ef0cf5465fff02e5e70c1c16915f34aa63a96bd0f95b44ad4f240feb87f9ce2ff61c53eca949faf2c0f91c82dd549b5fd3da7e75762f695161fca0add875565a4701eac86d2dfae64ceb40f46bac2463c4198991b7bde3e376c2b643c2d61bfad6d55c2ceb90fb8301d5e4abc281d14560aca933d7a1e8e284b68e8ec7571f7352ed2f38a09fe9ce663f895a31d3d35168b09cdae3d1a266c3bf1b43d80e849b630a27842a6eba65cd94c6d907f58d3cc3d88cbb0084186afbfff602d1bfda4262447410bce42f188b8cc3cf833a8b69c9edb2ead392a28de454036c7106d1775a1d0045e802d9c754e288e46f58b7a26803968eb23efe9cfe9d8e8e691afb6cdfb44079a1d354ab3e0fe5114fd8f4af36fe1c5dbf7278df45e09b12dd1970fa48d92331f30d58dd90ea4c7c097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7b936e3d98ca52cdb5bcbda0ee1dc99c57970d3d58a1192fea956fe3f0e342527419b585a0591547306157ba2370af07db8b81a6f1b99971baeadd3dbabdae15e50225441a0002df55cb6d10fedf19e454b3034eac38a3d686fba8da002922072b166801ceae2185f348f3cc496499737cfad4213143f7c21ab24ba4a033a985bb88b28f3bc9cb26d0a7f5f183f01fb3941c6f9edf0d9caf885df8dc6d039232c5c72d2fb0122bf65c41ee673121a2a26666b86e2e62b028afbeef78577b9067821b58717b81baeb2dff406320b7bd0213a9094097d0a7054703fe869502d1a16ad723358f75898c001ff77bab36a82ae58916780a9d04c1d5e85716b1048426019f414032ebe57d257dfd270cc6eecd4500206a71d7700edd1b69596626673cbb24e5a5d14fa2fe0f9ae3827dc697396a9098dc81cfed2f83d7e093be9cb3e7ac0a64914e807f0d453d09635013637fc210c8f6e543a9f001eafb209c134694dfc0711f49f357b903ec1f1e930dae3fd2e146eb0d6635da18c552355798134d26a8cba74745e242fb82718026a5ffa12bf21b4ab96e5eecfb46b0f4d7e79bbd165ed77080d84fa1542df1287d119bca5434f5bd8d36947f58ebbd2c4200e735fb20977c8761ea4bed524946246cdba7fed1414b8ed85b0d5be54402312ea3e0cf5d571cc2d804889537f6494a0925ea1cc84f37bb300e3ddc867959af24cc933892a6efa675a451e0a0886be225d4880ca25aa1237bd7c23daa5f3746cb229c56912384c7992a5cc939906ae7a2e16f6641d5cd5e4dc9bca0581efbfe943e0e22cf28874dd20a0fd95ebadf35e8bd8562a7a53632d44850f5ccbcf0a09f82fcd7c5746e83c9bdeb06f4d18b0e3aed89c7fe28220bd6a3e9851c196526b88741ceed354bdafd0f1716df5a90f144cb56912d1b49a4d45ade3618ca0ec91a22912f2ccd2e820e6fd5d1cceabbe8d072a7c2f75ec46674c081d1ac134c789340b6db4bff8da147b5924e6db76f3206b45f7a2021d9648d736059;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h76c96bd627c12d2c50db4f1c29a084f420f81ff227b5ebeb03d9c1faca8a30dc2020ad83368f6ad93aa1f89ff1fb430c275cce7ddfd169b050c1a02723f346902ffd847dd18534a94f225ff1877cafec8ba8223cdd12980b3a8f8f331e4d24e66999feb0196e5319632b3e6f7216b895982900706531d6bc9f353774d0bfdc714600503e55a8812acb0e615ca8ec976c7b4df5d29fa2fa2cc341e15cacb67cca2a032dd33e0e6bf808bf336c760902bf153af02cf23a6a95c52046cadc219bd3ae66915df4a0f15f2eb1c2abd2027c6df74dbedea7ec682c499157ddae078f16452c1db1095f98b8640b4363d67a3a90e49ee9e3b1f6dbe8924878cfaa8a29638ec7e25be42915081df8323166b15d9bb63a23161900f10ad7bb53e73ee2c9fce560272f342635b80172f500bfe58686ab0a96b135d35eae6c26faba9e4aab754215c85f212a5b7d6d3c9d8d44b8b177d03f5343a2e0fa2a5029861f2cf2fc9fc6057820bf0da63db6320dfb12e591b5b4c6851e3e414ca8474aaeded4d3d4473a7ecdbbe9c4b8f6e0968e2b14de2e72d47426554a3d449fe46602fd432d1e3b5a8dc666589a269b5e25afc9ea7b5bf95547152ddad6bf322fa29e9e978b476c9b7bdca79014c218baf0d2e824f648c24ad232426398915e1ebbd8b12285e1c6369c15bb78d0f10e486939e22865e8df73df182b8972c83725981bfcea4ff96de4e4d2637bf6e33761f9dfbd6bbf62f3b83ccebd80049198aefd78eaf0f5695c7b3907eb1f3b800464710f57da7458a223adc526f9c0e22ab95be2c6b00802b978abc257758803771bd34d8506f11a473f24f140686970f25402f7201f9b2677263486cd3a1fb27da63c3cff8dd5552699731677142eb08eb6996b244faed6a26bf6dbc8a35f61b08e000a1e3f78df932cf5c0058904f7a1c3a9b8d6c7811a19affe338be56bf75ccffb5b20710cf59c4f63be625ab58b63ec741143c8d3f75edc93cae546fd487ac19098bbf9ca7643f5513f8d4eef66f805;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h80de19127177a4d5b5d0628f7314e8716f71cb6affba457ccd9e0aabbe69fa0188146f8ceeb7d83fb6784e7c0c50ff4c66bdd982b14d71c1718b45a7074501e5c2c47f72d7be422c8648c8e71ea55e1aff2bcfe492ccbbf66993fd71f0a5dba4a3b05fbaf6f02626a94b23ba7f916c890301ae1f2086f7bea66bc3192654742c22d86b1533993292aaa09edd86a23bbdd6c40ebcceaed4d364c3448d8163dafe6010262674df6c9918a39af4635125333beee9791c65b1b53e094b16a2a2c6f555a6d277e257d0bf13a4c77f8eb57a559fa37553c7baed3deeaa66fc29d1eb261434db1dfabcbecf95a0d62671d0d59020c0e195ee341c80e610593b46fd602401a52df7b74d66fb14a6bf35e13aea54feb9b598fa609d29e45474821c727404d0594b0c3577ca36a21876e684df4560efd560bb311f68fd1b12641101820f553d195968a0d6b26231f9458920e2ad33cfd62fdcf35f8639f2cb96b016b762cafc57f5bc993c884cdd0f77a761acdd9832f670959e5b288376e464e9c4395f436e6124bbb4616aaad4d257b01ac869da4c0e1a35ed2981ddc571b385ac86dab9d64ebb3d0c6fcaf5f70724e2ccb1ee60a338a0d514d5e5f9ee095d815385249149b09a56a8f201d1efcb286a05f7b06a199fe4e94aeba96f8a4e1acf655f1b71f4fefc605b64b9663bb7fd3a58d27c45d690e7f38d621516a3189ac403ccbfb3f6cc314062c3ca8e3d4f73c0afd33d2e2f47518edd1632d8d02502f5e73b35a79784718dd57896d8f579dd6a9217df685bc84cd4b7a4147d3acee7a322b527c670a461939fa33d2038e3eb9ab393ca466a91301ab2ac5c30492a41cd008f4c6c1469d400408aa4611e9d51a110409a5ecddc312205108ff49918fa25903be70e569d21b43ee9c3e9f50c4ad9acec2423ed87be1df24a8a95338b244419c838750e5b15f62e1d65bb8a92f442b04d05b0622d46fea3042d1754295eb1a44162799b63950765bf5c22e096c2828a4bf0d2cd92cbf3d4e3dbfcfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h44b58e1452b85456e8872f9816f6addbf561ee4cf22feddb31ea0d99d33ad1867e4371f11187f2647d1923c062b1893fa73637d1cacc6f40c6343b9061a2ccca5198cad0c7d3dd2484a6356e664ab34bca2ab57206559fd0984b29030e278149757685e14667d7a639a64172a5825ea26710bd6db8beb12625eab40d34f2805d2c28f0b3b8644c80b8d3e62fdaab2f471649f9a0c68c53414f3cd564543bb0849e65dce55f4d1a52ae125757abcb8dc9d027b99a7e2e33f3e014767d46f9146edf9f548aa2a8e42c0a34b7a32260f3f3dd696dc90ae03671d293d2186f43d7771e66f19410f0a79600a35fdcafe066d6394b14048510acf02cffb9ae4576614f5ac469101bff579c6e00bce61f8b02d0073e37dfac969c600214d6c8f247977896f57fded660712199bb09a23046d6d8a6e578345b4d6e07b55cb015d2fa4fbe9734587b397647f5b94f9e3157dcc5923d65d6cb3e859a6da851feb23a9927d8b2e9a6fdfb14837269db3aefca1fff5d1b413a7639c19c3c31885e62c761bdf82c5efe396247716a616a2dcf177562c85a53e11da04811a2b1ea127ca487f0bfa164a63e50ae2faca4c15207c731acce28f09fdc8b7acdee27f24ed048f90b32b598802f068c34fc24e4d3fbc7c6643e12f16180620ef38b9d382fe6d1738c90696d018426cc0918e819178ba6edbb423b3daefe6dc2e3c3e8a3a0d1e436eeaf8ebba9d7bceec376d9e56310657e91b3ba59c739fc52172144c67493ad82ca12dba958b6083e05e7ae78b74895bffeb083ea1d9a79738da4197dd2285055f6c49863c24803a24c98b0e5ae7a61251b604117d70b32147742c458289a1c1932484ce046e518767f0df8edd40c664ab499144a05e09e750e5e5af970abfd42e8a019f3c5fe9ce7987760773a9b7e3bf1a4925666177d3326fc03a4cb44f1d570e15b65dc2c242a201cf378ba365d2107d5c8ef6b1ae2f2ef19319e0a4392a3e6752f72987e432b40311df0fc33a9f37857ebc9a342a4b34ecd64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h982da9a58fd038559f5c79441efed83ca015b152eab2ca3c236c2ea1f93f1564907fd03436625f6eb16ddc93023f65e7a21eb4a537faddc39751a4289588c313d734ce12c104fb78d10ea0f31ab08eb8f23b8b6becb84a5b698006a007bb5e4062562ea62a804484a5a52422f99ca628423a6ef2e9dac68f4b727dab401b726e7572187444fc09322f77a6c6af781b828b07126027a12db271dff06cfc086dabfda7f1747ccf58ddc48106420a7f8ae8d3d89e5f272cd8dc1297092b23e86488c9f2ee3b2207f9cd7048c120bd8d5c5e33fbf2d34d4bc5b0ecb6991fb0ad4abf710f92cd77bf136822e8e86e759afd9167c119a83da7933dae00ba6216e982e0485ddba72ee78fd5334f3d493cdac22798b55e31d3eba7aaf0e82a0c2fa946dc1869a26b9eb3f30bf0b258e5d7051a0cac18c2b8cb74c3d331ab629e56e643844e3595319633891521aa9abd347ffcdd9b297a017a68679b422475d5f6f4dc938ada218e2e3ea988aacc8f525f457ee35175a79b7560b14f81abf1d5028e490c7c2c2dff19df0c0c0762dc4186cdb6a73102cd78dd1a9de93ac0d0f8e42576ae9e084ca65b0716b34b059a092d8013ae5aba8b04abe99ca284bb96da82e765009fb42ad15d50a4ba51eb5b321f960c0e2f6e025e8e720beb7eb9b0da4c3d9afa1d957c2c0fab021f0777dc3bd8025015bd1548c1587ec22214a96e3b8368d9ecc8f3cf3c8dbd5d5c58a7fd2b7a72b4f2a18a2dbbd82ffb4e762c50ae6fd8dccb234d3bb85f8866bc437e25c715d698551c08bafba3a3d818fa6f7d1e7934a92517dc6ac435d63e946bec9cc0d6b20453d3b9682751d8b4f6779972e38b4db264ca82ce2132f610d434ecfbf1f56501ab4482be7e04bff40ef14a0973d995839c1c10a03abeaa5b51b19a134c3b4f2ad2908b9d89da66d8f9e926502be7c6a22e6e181f5d37b88b9a75a760e8969eebeaddf9830265e3bb725bb2a33a57085529d2eed952ea5687b3b31d28ea165fb451b034ee769bdd12fe11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbc5442e50b2c20ea7783608bee4db4df191ee155102d7e9cf6edab9ed819154bbeb07d22ae3da761ada62c6e14b597291419210291ff2690cc7acb33303302b78173fb40f37eb2c9569ad60b3bb35aafa031c5972617bf969516162a2a60fe5be6a78e0dc0f9ccc38b10803f2947390d0661ccda294fe4ba3f5675ef1c36f2109fb27feb9b9a3ca568d9b0d71a961d031f75cbe5f0ab9fd8c0c2c73fc2454bc8523a6370e769da277512bbdf5f7eb73279bb4932a144f87d890918eef10cedc225742d9e69528b42d0bf0f0c89b62718ee5784229bbfb43965d157c331d6dc9c400fab44de5cc9b1146feb8bc9ecfbf6e86c2b46ad2b629e9d4cd835453f666ce9fb9561f4acd2241c9293a5f25d3b2fdd410d6cd9877f5adf3c1c9d1bb71f799ff4a4232a49f176ca90c2cc941dac14152aa22b6b07519d1cc0da4b55b70d804927fd26648a6147889bbf506d6ca5fc08a39d5b40b6b7164cb0ed241ef71aee3939f01e2a4baeefca70fe1b83e1413578f569e1e8eba8a8938e4dd1967902c8036066e6f6d364534a12f9ea85885029f467dd4643eadcc68fe1cb6e4d30ee240e76f6ea50378ef548c59ac1b93340aa33acb099a44441887823e6e30c6f86f5026995a2616124c608c1b789d301a93cbe7b0d01f9446d1ed3d3c5e98750433edf2b78794167202674cc4d28873644a5209c3135cd9aec219f13da7141a3811eb29f9e3b98c1041b2832b1a56ceb673db5bb24e29f13019028b7c7bb02910c778d3e5d094fc3a4ddfec94b51cdc4a92c23ace7d229360ae3a8f7e9f33e349dd580151aab29cf669d151c6832dda43eb550ae37dbd826ec5b1d36b8fb8889168933530a9dbfcfec7cb5e14988c609716eaae01f4661d4bfa4c145b1d3ec33c2f32f1afe0967a2ff17b1d776057d0cb1e791bd22c2549e50a663dc254133288a3d54f2294a1039c713a5838fdd8ecf5993c0de0e28be7ca4437a6b77527c45b9877feb6459fb741a34a83274000d6bf82eb46a832061f493fb02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hff438207ef7918b4ea95bd981905e510ac627204129f5dd5cfc9a0144c354762520655d68bfe70f28d94b9e1bb7d2b87f63e1e25587390d5d62ac71734f24e24bc206fb7b1cf4b144ce66df49112b2bc2ed50a5b5da47465b78b11fcad6653ffe454d306dd91b77522bd3c4d517fd2a33cbf7860f948481418b74ac5e3674188f844f1e9f422d29f0a633d7683701d573a4c8cbcda994ebba03518c3abbb64cb09b15061590eb48a49df53ab4812b2cafd22ad9ac506f48adb7cfb20de7f689cd62482579a0fed3ed46c27f1182fc92ff3c57085b9f27bbf74aa4437948945fe791ca75f93b8061b86b2f5f619f317a9a20938cded6839bdf4ce1c0b4f6937ab19c7c3db3a576d6bd739744654ebd0011a7b01b7b6c9a7ae2dc54eb65e4dd352bf9c042583b7af7b9861ff49652f415bd192c831565b5dce24d98aca8497f13fdab92453c03fa77c822094f1bf52cd190830bb4ffb4449428587397c68619bfb2ed7b14f0ce9446bef2e87eccb043d426135f3571691b53be0dd623b66362a31333e551eff0ce9084f5b01d64a8796bde50b00aed6d864f17eef349d769d47997b1227347c4407505310b62261c7eb7787da37e67d9a05e5e5291613cc14224c042b3406f644d5788f22fbb425fa39a186fd975e8394a17d7b2f0ec73866815163f60427455686d91c3542f05a722b67998e7fb9cab9bed7fd87c56bbe3acfd1f9c588cb35ada7ea09ec60a42e4f67510fa0f10e1e27f58fade9ed3025b9ec7b4c2fb60c9cd687a4734665a48d583d1cf2dd3a229a0307c34f0ad03887b8b16a7eb2d99969d0bfe62f645c771fb517247c485e4dcc14b74c0341d578349981425d95e9bbf67418de06bf3f9b09d0c10b5d4bcc228b0c27772448a05d6977271b4240fdfcc8b18ad14e6096b0513a633a650c65a33fae484672585dcade7dd1a15942ca3d95ee93d32384341041f76ab54a51b0f4b9301fdca37cf2de7497394a60f7fda5fc19cfb8cbf3d82b2a8ebcb85e55ca73d5c95cfe7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8874b9dca584fe9fa5f41f5533b3b2be53794a4eaa03ba33d41964b571af769065afe7605cc08afc228b7260f899124bf3bcd86fe54626a9f1a4af851f7d78a38c43691023ffc0c0e09aaeccaad67448ce71df858b42b38f7649ef350fee915dff403c12b12ea2b8c00a6e49abdf2ad1d5dd47cac4a61e8322f62eeabd0ad02923b272504b8656ca695d26231438f7b4a25d24d3155f2f9d181a54458f7ba2e8f503a1ac55583bf6c4cfb7810e337ccd6ce9f81373b4d1ab2b7bbbe22754760834bd5adc5e23c3ac27a7b2eac9080f7a88d998f1722815ae15e1b5a842040f7632d5ce91ebd6d27f61b368136804a9b67f0150fa3f3608ab5e23e37e442b44440e71e977fd209209edf28807c0aef27b3a974e86cb51c0960c8a239434b16217ed516b9e67dec075c2efafe4f1adbc17e9dc4dc9f17b32932a6d1d1afa6f04911bbf35beb7df04c71309aa02619a44f39a5f324d73378efd24c107caffd398f365f975588f4ae2b676b256d6eb1b80a270f59c504dcca6cf062dde67a3626b74398e00fc9eab6f264db537b664b8d4cfcaa01225be4b26828bcb3b7091315990dd365bc6530f3b18235b7212338bd0469882928feda148c8d365662e9bb481c0e87a17fa005f71c947b73a511f324a44d29fa2238491664bb087f4b5a1f6b1d4c1782a46a5500056f2e30dbdf3aa455d5959199240585154d7b54aa46b4137779765e9f7eb7ae104b3e46f2573938464b64d6cbb903513d63a03e30b98d319e31427197522f1f59037316335ecdf14990228b74c26f64536078e6baaace24f30d54f2132c447a4a580414138a3bb544e00fd34bd5c2e130da5b422ee454993d89ac083bc5338d346f3b76800a6aca6a7e6e074426f65147eb2c9cfd608a7ac55328ef050b4b990dfd90318a9c7237b43c22ef0c1edf63bf1aedb8f1f357ef47cc70b66c4e06617eda80784870caeef2543a39c5f238791a38e6709cd88e835441535bafee6468e391f6a0374ce9797be1ab767bcb47de10e18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5aa43feb0c930d14a49db4609aff07296840fe1c6a692aa1fffa632920fc3a853d35c91711013ab347ef8c0a8ee598e44e5a2f946a4d1fcdc698b2e85bb98c08e7995e0f318a3c41db174fcafb9e4f996b68d5e4774fcf6ce3b50924fb39d2d35d82a5158a0fca1d14550f6ed3fb781e9778bed86f084df3d85302ce15d7234a53a189b1f0f59ddb556fd602f0522cc77768ba51258e353a23647188045575e8cb077f26e7622e3b7526721848afaebba8fe30502a3e5d7b796ae2274b4453e2cd07af024722d1bd88b2a883a3d2b7c57215828979478b6bf54b183ce416bfc0e33cd4b04729320b6d3614e9b2bc38765a56e6a9ccbe6f6956f3ed3d4ca0d08a9f262fb262827e1c6b09f16143e0a67b9febbcc2f6b3a632628c9c7bbb42852169f6faf1dc3ed47d8160bf81b3e977bcc5b8ba48b2375082a2ca77ab0a55caa3e52148340f2a0167d1b212119408db81a53bee84b1fe223fcc44a8cf70df2b25d7b43be06862df2bc7a38a36cd045824c043564aa5418b007834acd9b0235f384bdbf1f1128e690ff7cb337cc2e89f6a19af56ccb4cda6d5eeeef54cb95451ebdfde591c0ed9750c3688125f4161075d9eedc36c09792660ed07403cdde857a6ddd042a918b0bfc01885a62a1fa307eb8c23c58554700d23bb20c8d005540ffe3616cd9e987f4707dd589faf07501a7caee0b713cd62375c932e85e43dfdb21dab55af14ff6204ba542c88ac42bd9f1729052d14d29765cec07dff7d8d080cc7348ab0ab3badd4320c28d4cd29b9e7b1097178488ae4e0a1cc300b9477769554453207d29dc7ca1b8321f7fce10eec2d66045b2038e7b04c706aa9c5b4370eda0075a1e0afbca6ee2ca6d9f4a182395e5f6de28447352a0f1c57b8a251979d1d62df6e6f906fb8be90f4a0887ff2d6b27c3e5b2f1d407e878807f3ddf7cb8821d75c7cba4d56bab89580cad780b4322e5055f3846819c45373c51cb2a01dedbf4d3677b52ffd82028786f3539a63ad5330fb57a306b362b170;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h60b5548762a5315486e59a9cb4cfdc313333ea722c5c98dd40a58f9f6e5a8efd06c9d6c129803ed0fcee68f47f309fbe670c5f79224e64e95b69611c87b14d6ccb77b30c829350100b97cf74134959f5807f887d9579fe3aaceae69ecf3e3997e701c951634cfc8a70e1a4ea6c0e10dadec4150faea171ef0eff314684a9c103907e2ffc9e9fa99e097a627d0f5f29342c9ab873ac15f476da6b43e9fdbcc004790c3ea7f9e026135526e47a94722048e57071a20527aa84bf9f0f601eadf67d391a05f0f73de9c40b392814994a5c6ca0d73d2bfcf5ffd7c92467ea057cce9b3d06fc822433a61022c2e8e55e0271e436bdc5548115a73e3bc8f70cbc4758cf18ead91d17e9dad9bb32632e212ac744ff4c7a7f87d471a2745c73714cd8edfc84fc42c207f9cfb372e5d4621fe581ff2e5d1e00fc05fd282bbe8fd75523c2fe5ee3aa376154a978449616e910a0c8ffc0fb2bbb5157aef84d6851059ac5912be652a1d8a99000912bbc022b2cbd76b1a873fb1925f845cff4399cfad96f2e38d1d5ae519063123eece5c73357fccec9cc500f5a3b62c619aa70485007f2c311946fd2ee93af0a127772bcfa6a5d81334b029e17cc9945d9f2dda8b061e397abfe42bdab4a9bdccf7f454ef7d4284574928d16dd3471eb0e2344c92820fa9c24dbceca546644192c2a9666842f4d69fcc57eb0c9e98c5f5d4966311195a79080f0d5cc0b999a4b57f219b0a4f09e3f840b63a70fb8b932be84509b393d4f530a4863500e8b01bc16ee5c083dedaaddceaff9025e2c917a4802f33cf7d1146ff3693c9e6c1dcec4532731f4b2ae6028b22d9fd91ff8c8cc0d09b0d2e4b0683c595f5d623089ecca55cab499ed6dda8e24a86f0acb0b5ecd345677fcb1e537322e157ca509f5edf8144de2fc339ecc913299ced62fc2737c11030fae1388f2e35ce892bbaec6a957603ce7a5f555afd524397f40cb4de851d712ffcdbcab4c2bc8790fa51384ede56aa45e276368e3643cf615307628a2ef0478;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hee2592e86c5c0db964504cbb285a312c8f5c2926a4c440d2e42dae378af3e7325dbc23c2265bb47e5120ca2d6313cda1b71cf38e22b351d280283cb9335b00bf6a6a860596a1007819f3d7070c72e92ce2631d284b09158e60d09213b442a44ca145cfad83e60824d90823909d1007fce03f6896ad99d07d027f06e6a4a508cc05f10daba5a81d1cde61953db78e79ed1b872e4faec5d767ba86752ef13bfac10f34c7175530747e86a7ed71760ace3210ea5e408f190b5cf883c8812297088946e5ffac4c6a17b425d931452cdccc9877fd84fcb3896136e52ae0bbb63c4905b22d7e05de4537d6074c0ceb9d69f1868993a2d498a4796137f5cd7f11879b2744c5698ee730fccee81205a1a6db2115e8aaeb594d7c818cf6c380ada8afe58dbbb7fd5354f1dd33df251dd6360e2955bcfaec74b7c190853b2162daa726669977a5356d930859d46abad4606ccc76ad7abb0403df1a7aed815836f1195c4c599a39698674c97dd5c5846d180398d6191eb884179f65a46ab2a293f5b051fe61c3ceeb76d30361fa7e6736806d3bbcabc80fbb4ad86097ea93525b20beafba9a1a1674e503c28c8f6271570ea1e202abe6aa2700ac8027d654d0c97a6e3b6c1569c532d3049599169ff5124993354c6f391f1a12c01d21db843a79044850d99677d77e28ca51c7818b539f3d9187b69bfe5cb48aa5e5ed70063685b4508860ed50461b69a1e1be323091d5357f375622a343027f98f60750eb43cade655244483ac886fd673d218d9abe8cf2eaafdd2ca3d8c965bc82002d1b6e66e6c44c0dd55ea71c22166718ea8e68e714cb345da78e2854b4e4a9c4ef414dea180cf3db3b29eed46cdffd1a67ca3c02cc6fa52c7a1cfe7273a69a364af2598bb3634ce6468ab078a5e2a699ef9cc23b302c9390bf2d7d1235ad4da8c25606866562b8ed9a02faed550a7862d16316d84b39de2bcccd3a163bbaa0681b70a036fdd8730d959efed5d500c5b39a0dc866c39ccd5f9eefc9c32481906b2986;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h81b9596e37e74f91853cbe506d480715c0bc5166e99d14f16fd020ee7374549c2b8b8ddda41397d048b94b1e370331a7316b0d2e1dd7ac70557f17f6978b2173d2ced7bddd921c5c277466e78989636ec9c3b241180391c3e586e59ec300ba046d2363a775ffeac0dda950d5cd6aa16a9bef6154d11f87a8e05c8336ce95f6ce2ea18414070136179fc9616a9ad8eae1f0fc142e39c097fe7b885059deb69be98de787350aed04ded270f3a8facb3a09638e8e0ee60c1777d73c377b630638f112b7f357fb89b965b540844d366a432398bc606146d2481e4b27d24cd2f8013d94ae165e35a925291e48e2a690129fe21a0a515293f28339d2d0257a0c9111c8ab061b6312603f4bee367739195014b97a97854b3efa0d886ca9a330b42d00fe0c57ab165ec8b8c74c46bd3e414e85090e551ebf37474bade070f6b41ea970a4f380acedf4534203cae6aa5c296fa4019029af5fff33e328546d6b29214cd38573ae74617126848266ad951d9d342d3754dc6547e117342987e29953dbf209745265d77915503519ff7f80f94c1b885c8c566e2ff2a3961e53c9bf9230bd164c216bc889b6f0ba0a31d60075cd5808602a31d2b8504821046b32c57a0d164870243a7484289d366542c69b572be7ea62ade8f9b1fbdafc6ceed8cf59aa39bcb2c0e96a2827d9916b246e9c06294e09d625944a4fa4af89a752780532efeaa74f1367ae96228f1d074dbf9b745a415fed7458c7aaf2dac309594d382221ac9d45bb67421f68422607e4d26f9bce314aef6c164114900e0e471dbef44587fd2fcb844ec6367981569c66319a6c05fb8992501abc0d3eb4a135be64631f5709c6d183ed5fdda29b99ec4e1156ed105412f8ddd2931ac30313e7c6c3f1c7ff6973e3292866b00ee6bdecad6904605d5e0216775647a8cda9e32af8162cd0a5181cda5d64d830b4ae92500dc3df6d022c343ac8af84fb9a3a5f2e60b3bf0d38323b8b4eb227c2cd8394a3013233816b4820978cd4bfe0170fad313e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h606d9e7ee37813371c247ef9601961c34a1fff0b0e2eff61066d75c4cf5f866b72704ef5c365f38d70ffbd70280bcb97a204822daae0bee463367149265c644321d60ebfa882563f9877da07ff0c7ea1ad24cb92eac4d3f200122c710490d333a2f6da27d2b01d36b7547c940dac1c9e959b10d588027e9927695de1ad2ee859b5ddcfaa348d0db30364303105318c70869322a5c757dd6b4daca609673e0cb8ff77c228c4ddcc0605e8296db20b365f4191fe41937b9faa7a0afbd52d6eb4813f6a6034fc515979bd168a54d41057378ffe67a34b3121c50844977ba44afcf1b7847b72b6817c1825eac9037eee6ae0f0ec0de1adb506861be76f8e21500f6c217edfb8d63ae66f21270c565a3f7148516dbaeed675832bf2921a2004d620020dca4346f0bde238a1ea1c640ef18dae44c2bf9dd814e692ba5fbb016593dcf062d5fb5c1b1b525709ba4c9847109e07c715e1abe2e480d0461ce18d3e91874bb12af02d5a8eb302a65cf10297a12a6e4e27376c27c17affac7c5e28b8b0483286eb2e98ba220932e41ec1a91c5633c360c3727db4b7872f1d85a5fcc1547bfb7b1e2531e9a8b609afebc984e2982458843e77d760de2044569e9db8a70614b9700566a48d5e968d0d4a9625de986ffdbccc3f52af70df6d3ae8904f18b4a5d001a3ac678fe24ad1a3d543afc8e7010576fde73db1388861d059a73caa7e9c8d1ff1ad4df4a2c68e77fb2a3e93722a23890d28b039dff5874e53a9d47db3e7c520293d5506d1ea603d5bb4eea31917fa893594b658df2fa90d498c720f6f1afab2e1d407d6e631d2294bcb7764ab18261d6b6cc56e94b275f9aa3d2cc239fdefadc22d612f0e88e7a4ebb8be58049c3c28fb238468e6684f579278b283477a383f82d0a4bd5b3d8e87cea517b3a0938eb918a9b763108db5d2f0019f7e7a236fc0ec25c1d7422e737794ffa72101267ab9c829a2345d22c3d0bb5b6c82e96814f280923b87501eaa0eab377e42049b46d7cc482ca06f8a3984;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb84f719d1103ece812b9a2c76256bac8d8fa5f77a5ada922520c4b434c05f17524883862a8bd918f3a8e0c73e25c00c35f0e9977ce8fd444ef15fff8d1237a587e6b96c5e4ad150307aa38cfeb25ff30c3f34dff1c692a907afbbf58f0c647c26f50de22785d79980a22d90701eb351b2bf8bb4e57502be91a00d7a1616f1a188a9ae78fb49c51105e0eb64f986af46ebd7829417a66b87179f552ee7964e074ec94348e2ab2889acd8ec9cf757a1cea98e95b4511e7838745ecb59643e33f383c686bf494047bffb53f17d76fcbf013019c6383cb4d3aae4bf210e39446ecb5d55eb6d7058430ac5af7cb48a4a311cc0db4aceee379121a85c50ef79e0be84f107de4a96068b1a86f5a26a0963302dc8d8b5783a9a9113858571ee95d86795f79d4e1810ee9cbb430326fc079c10d28d25dedafb9b326784cf11e0c27963bcf89402b1294484bf941b998e430c3b3448cd8c6be93e0f2c1a7f317c2e71c2f40d714ca7037a19538afdd588e5d2b2883f0b9bc53bf12e3c892203caaabf794fde88e94cf5b485d31ea7be0b4550f38dd9250e50486b76b5dcb1191cf49992e28f346ab31bd85fadafdafd83ebf0d2ecc9137c7a514876247ea8aba25fb8576d57fcd2ad9457c68c80696279aedfb22dab017de5d5529794c71cbe230ad0dc1eb597f66876e09ab3c5b6cdb93b756e432aaf90faa96cb389ccee91e65407110e8a168bc65e29e154abc51b9a0b2fef051c55185f14d0942dcc8cbfb5c42e81822221e434e250c060fed4b06e0ab2ff46027396ed1920118c6cc9e8e928b8866be7f1b3639e21cf61a25ed86ad2654bec1ee4641684d74eb55d5e07394ea62d2081a4fcb9e5b4c312783de2d6e70dcbdb47e24d1283ef8a00f172c5464e1cb943c880e2b460536d71ba0321fd8d44ce8f743e62968d63d6d0fc36a1fc9a55fe57fb0c066026b14f3b46e30bcf0a6b284dfbd49f7ccb9c80dffc07e5128a327a893760c4b380e6a359484ac5b33c1563756751379455a10a2f8ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1df7863d389e481cddc047013a79cac4930336d2d611eeba1ce5da357dc5a5cc837bab5d3bfc9076351d7aba23de6c5021ee3d5b58ac080c96800ad6ce781819124c0fd1d264d0ee5c5e05b9128425e2f3f50965107c212d125bbd5e94026d0585a2499b01ee1c1d32b5dd3ce3fa3fab12ed0446a07931bd440b0fec2ce9e41b9f9a85f851278635de532bbaefac038962c7605851b904183cfdd834e88dd046ce23efd6f5a100e58ec6aafcdd0850939c8146243f8b34f06cc0eab459e452e0aab921fa3f6bf0a1e986dc51d256a3dce877f4dc1c28b7aae7b9ad4a47ecc0b68616a645cb1a52e21b209c50fd1cfcb935a479f5ce3d033b69b4819057a46db9b378633851acfa596701d83b9d7be11d1dfa07429b55bf3dcdca99a9a0bded331046d46b00a79afae5d8b188b1ec1c8780d05a5e0e3df8f79e878267edbc6f0c233367ae3207c079f0cb08ab8840bc27769e993efdb94936f43803f6759fe1f8ba594364da329f9c4a4ee2536ea72f6fbbf706f11d38d88bb7bb2d75b943af9e3a6cec45f2fbaecd017cdea7cc54fceceb4cfb4e9a201887232fdcad43c80121f34ba9f37bc9681e18b0a72adcb742601391051671ca5c2d08a0d10d75a41079888253254cbbcea14f61a184d823979f2cfc1efb7767c59cd3206477f447e3474e5c570c533ab523c0fa3e9e9c8690e352cc1bef2ac8600262ff83e9c9eaf9ff4aeb936dab88c4fd471752a03b8d985250310f1ab50ac6007c39ad63fcd3e51bf99e97d170f49f2bfa68ce167806ad4b1e08844b119433f9e3d7156a71e7f10ca67a0e32a45a7f459c7f9e1c35d5586e5ed6deb21781b1db43cc0f447e3ded5d41737ba335751b125df2241d8a69ccd5913a95c9515485291be150abd8426f030a2a751e82c5f46568fc0ed98d515da4786deb41d769863e8dd7bacdfa97b2e918d7425d21d41e95b592648e33d2bf514d8028621032694280fe02738def38359a26d93dd1beda57b6fdc50be21e7096fdd2951111402af388;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc6fe2c305d030b8f2250d1a9ffba78dc224626c5cebf0e40154da3128b69f7871d0cd86735ddf63587ed8be6d6206fbda0094860e80277e7b5c6783286acd9f890083037d0746ef4660a71f5036bee64c64ffb98ac7d8ef935c7d541e107751bcf89fc0273328b8b67da19fd56ecd4bb16b83fd86cf8b3c673c9a6ec76573b9448baae3e5716a1ee255aea9d85cd95fa8da4302844b614f25df37ef152e722f5564fb6594d156c73c1db991f0b8a147710e22f7e6bc0caa9c2f39e3daaee64ceb146e1196468f6e8f51c2f8353d38e387beca82ba0c73fa117972c26df62f03bb4cda554eaa1f1796c3927136b26b98458ce6c9d1dc0f8cc274e39fce16afa680ba4767a98d457beae81fc3a9ad94bf05267b40ea12716d1ca05e9eb9d5c6aca5fffbb54344002ef0237739b9f256de25a5726303dca253e333d5121d3fbe16789b4e4d461319d5cbc6e3cc8ea8763443a3701c53c6615f88577be5b07c766eea50d731e0aef96775475a48d50c96fb917d86061dca0f86fce25aed5d002af137e235feaaaf54cdd32d3f26063933a72fcfb7be4a25fb42ca00334db91a1709410cf1c2dcc7899edbcf7928b5b347e19d40ccb7167161c6ead323af34e5ef3f8bb2d1c9b55671466914bd42223b863b2263bf437a3f058ef6ea5554673f3a530353e2601f7f479a3972456b45181175f0310da96fd82d92c7e877d50fbb432cb56f067cdde8550183a890836e6bc1c2d063b7adcfd231f25d5cb45a3fd42468bf463acadea38bd1570aa1d383eaef12355c3e201ea7dafa4a8fc3d7e4440426f4b6fe41e47187da98cd7c72c66e6cdf95d8611d28d92cadc4f18ed2805ef0324ef3f6df30c4f978ba09a8c939e5c26d52c95e6d862c18764c1b7b9a5218cc75d398efbad63c78d041927227484f3b96e050533440889fd165d59c301e8ad54b7f31d2168a8c39db64c1c6f194cb7ca9874b3107d32a27db71fd1ba3c07f2c0bbe4026e7ec231375e7f5bb6d4605fa5ddb44226145bfc8beba7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h54f6afd90c6ac3c5a181a515da20cbad6c435135702bca4bffac8f51a7979a4f78cb0ea1f1ae607d5cfd6af4065bba463c4374343bb51056908e5297b8924cb4cf1b3cb8913184316357ebfd5c258c9c1445176040a131537409ae7561451155b1279d07fe417a63b8e090384df7e873cb95d2482cff262caeaa3080777705d0da0178935d31b4542d9653aec48bbc614e43ab68044638b14cfa9d92abe732b7453d4da349567552f7809bc0d511347e2f9a843325a935d5ca3fc38d8ea199fa4bb4ee1b81eba435de9206fa0a7e480e6c9cb320ccc7767fdc75684cd1af80cf6b1dde879fc94652cd8be72180c788bc695e2a67444f487fb09dbc08b19c2e99915f9851fd7ae48a33bc66f1879c8b94cf7674b740f0534d91489d353bd7e1200174042cc5a584b102cf59625baf39e73321102908bf88a186fc1b5874be9533ca21c6e719a847e7adc4b2c55faf3058edc7bfa17c87eff11b75d3b757aa8ba67af7ff70c54616d7c6eaf1957332cdd09c7d3cc177fade9fe74c47b57098e2731a36102b748c92fa39f328df70a254dca4b92f7584dc0814037250fd8393095449f808670c57835658f18ce13bdccff43303cd76ae424776a4e60ca91029223cd39d3151dda7e8a2679fc8b6539a81084b388d95ab967c739be8f9740d528a2988cc1ecd299a9b07c8eea9666a6f7f7055e34783d04f48856b03063b3e868512776cf68d25f1ded299816b23d2d4dcf819780dfc68d895bb74825422eada62b2fba5a167eefc5be41e7ea502c7edf4f8d02446b788e1072207e35db0010eadd7bd11b65689e470d6b49111b4c24a34a2f4358cf64f91bbf68fec6efb57a0299f4f1f4916fabfbc718accd2f7ce7a1a1470aab697b0a64af8498c2125fef40a757c2639a75a9d771ee8943188c10e84968e79481ae6699952f69df49880aab45292da94a46c5ce1b3189c511b77097b4fbe48f8e20f5e5ec1060bc86e55c19d50985b39b3eb2497ffb5c55fea183aea428314f672e0c20ccad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4b4b3f534be37686ebdef653d1b909baab5a64dc79e65e438101a17cfdd6df7dbc013ff98636e965a07c226363ea02f778d08dc1dcbf5dfa42f7b68765078fa0d5d7cf0334cb9475f893d77de8b37e3d3948889d3fe520d6d253a9bc4c414959b572e53fccff1cbf83b92a74bd7996a52c8d1e9b38b14ae79052a4a85f84046a8084d8abfcd1d41d5b517daadcf46fa8b28c76e645cac232e9ab0262458ef1b0b685e951362dc72ac135c47fa9a53d0222e128bbf19db31d00c4200acf0b7533a0542f8e02a154cdf5a2c7e5b38052ba93e88bdd8cb5d504449e00baeafb63012312bba4dd79ca07e2d779def475826527a555e9f82d1c5b227657088bb94195433903d6d93f6611d35d0c0c0f053471fd4f794ac15943c01007d484618b3e4865eb51f0a951ea33b32157906c5059ea4596d8e721064f9e06b464a3268885f88290d0ca805ae974a0ee0f0b8a4ee9c64441e25dcc337d114b2e673415542b9db6a5ebc57851369abd10fb26a3af15021c03fc9a5a02c77327df671e544e44ad70c192f2b92d5c84872b99cb149e7be0ddddaa5d34a022c5847eeb3f121e0fa979981bc86b899363b02c547bf3e05d698bbd827f4f26df8d9b9c6f0825e5b44af44a428361d58ab9d67ea18038c79da21f36d994c9baeaec123ace56810b09f3e3822f6f7c78c3f453e4923151761e255f56110ccc528213de035de8ed41862ffbb94c4e66753702ac875368799f2258ae1e601904978fec644e54a025c9de64ddc1e0ed0ef618f5321714f0d2b1a1f9dc152761cb1b5e82f4fe109e0ea413f50cd25559346142a77c9d716ec2ecbc471ae56a666bdfd245c61d78ad34dc8d5e169c6924632c18eeba0da68b7c893eaf5bed69a89ccd14837d340019d44036766fe26f4ec13eef15322e452e7252b67b5a4dbf72439e823f1735191b6be67d2ba75cee198899061bcf9afe0173d9203403c335a11df4cc92e2d942ef06c2bcfa14ad2dbcbc95e3a07c4c5eab2ead64bcd2ae5c385d455c8342;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb71cbddf8c3d05ab139390c26286b9505459f22203a84fd9632cb2656cbf78ad6a1188afa6b2afa0d81532615d60c0161a3cd2e34d0e13392d9c9aa5c90a2ed413a94a46fd54195344a1cb6b3ceea01b095798089c17f46450771c16fe2039ed42955c32690e214af305adccd8a06475d9610f0c050f175f6d516c99891c2a071a5c354973ffc162dec1ba10d9b9c8000f81d8c2df04ef36f730b7d22f758dac05ba0788e6eca55f5a5311982d882646fd011c24a698c72b69de0244d138ef87bddc15c9867af423e1b7191f9639d714e91459173187059cbecc9b8e89cc04dffcc7ddbde2c3a9a78c7fc8adf328cec9107f48892f5cd920e55600b5e0277c3ab7b0096a516c963e018ba36b3b9efbaf4fc08127587b54db6b69553a365a3f5362344713fd1baea69bb20f1e213997c61514ac3f70b055d1b0292fa5802d26c1b4f3a47d01408a27eda87b3345eafc80e3189e9b3c57588614f8964eddad9d521fdb67185ad9a3c421c65cbbd922145902270b5aa2c5fb3be8c87d2b3f6ca1cf537baf60398a5e2ba6ba70cf080931fe7e26e93b786cd53588aea297b64f783920e78eff75c18a20beb1f35c1f8397f188720fa0a88c90d74a5b352563c8e98a56c9ce5573ca51428df7b81aa23beca45b5ea79bd87a07b59912b1d2744331214cc562e1e884a8be6677bdef3d7d4df06c148623272e872309c6f78a77b2ff4b238228c33cc1f19419f1a079a59c48b08ef4c1364a46b681d9d507eb75e15f6a3688dc2bce1d5c3e8a1e62a617e387e9f2fc6d604c6351e02082b2b8ce32f14d4697f7b976816f7a89a64dad9ea1e914d3e268eaf409d2093f19fbbb749967f62809aac2e5c3e3359506607952d568224e92f0f9b0990db56236df22e86ba71249733a1752961ec5d77ad2c5235775fd6d6c6a8e7a1d226b7110d6b238cc1b51eb05ff6f98936b4de3e9270b2b6137bbf0efa73d7343b9561d94bd0b6b1db27fc933d4c7fa7697327fe57775dbad1e593a3a38911823e6c9e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7b3c9e1ed3c91a21be3fa4cd7a1d47045d6dc75a6484732c9858e1ab7b6760638091595b7c193c2c4fe75a1aeacd12e13a01caa7e8bb2350f062cf5c3318cbbe698407f6bb06ea238c55f5f10f9bfac9dd36119e510fbe61fba4f714c0ded459e5c59e6f2fda81607fe9c8eff7e6ad6b800282a61883776b502aa9f67ee96cf288d7ef0e5376562dfe98b05d79d47fe1bd425c8b601a6c4cd85941cefa57aec4ed56d823657615eef225121d8ae5680976c6de3fad989091f4172ba0f6670850fd58d57c2fad4a09a8b7e03d356c2d914ff177ba12d36346a42dd3f7baf597c3ae93f3fba8ac00b6c79b3a65d718fb5c8a6bb0e9a2b78d3eeaba7c6dc7bf9cb7d03e7f79b648dab4cbe2d14c9214bed792f109be4e70755749a0a8f1f6b7e691cf5cef8f4c5056ac57fb157e8c9c93f6749bbcbbea14e143ae469d1e89fadb1b1e14ea42763020f2631c1a04afde5104147a821735f632b258b8d4111c829d3a3f3a1c1a85b18d0365cb4915708366a66a6fde651100f969b636f3a7aa54ffbb6b97a31859f8062259a0a3d9eba899687492a181089df8c1788d9e3151e52e5329e76e4ea047bfc4e8e2adfcc42cf4b7063fa56131f51224e67daf1ef1c817dd446710fa050759d28c1ad8d3338fd24adebcdbdeac64260c19b724b03c12cb62b1d0dca8bea20d4e49666d9502ffbd1a32c9cb09e2d00adac1323801da6483e3dd36ae4a6835cde8814c10bddd63d38b3ec93f550897efc0604950e7cfabb2026447a293b15963cf2dae2f063a4ed4ea4add7fd36ad13d4c15d6d09799f548a8d71ea0b386c0ffb44d8262f5d88153d0c56b7589e751c8397dd7c27b90e467ff3fe7490ea75503b5f8d5481ab8f6d46e805fec18ac9a710342765e8edde3d999c905168ab5e3ea0df8f6452b15686e585a188ab0f64550667f75a57cc76bcf0dd7e6218536a38cb37be8a1cfbb1e49ba90c4d1e8362deb48da8b23674b163f6193a4b6e7c81a02362dc7e0e5fddb663044653f45723b116958;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha912f1afe7d908edc9023418340df3a6e9ffa116df08094628717e5b699d901c3bec94538a2e5d74aa1c939ff8c830f649af779f2b73fcc3157553a386ccbe946b86aea027364a47acccacafac2328f05e017e742f27e39b9e5df9e38f6379beef0c762283f6eaf94df676bab1d5ee8d511e9f467fe99a4e04747a56c639f41bd95d81de3174f7a83263c265d9f09957f18f2719bc9e40b1e60bcbc86ce666a5aa8cacd288474be0b0507df8f08b7bf49e5d47e19665e065a7f0792ef661d6358f80cf40c057b93bac8f5f450100909679ec6ee92779ce8110419271730f2c3e1f930c32c1d15101ab44e91fa840f3d5f8abcbdb92b08f761ec8a662d467a25c4836ecddd87a90e02d8d84d576cfcdf5443fd3c1a03cf43be3f4f15eb055a422645d9908ea00195e52843615d1739f0459fc46cf782477d0c6854c093885fe78302ae6ac0e0d1d2b1dc57fe308965778bb8e48517a9e6a6cc9a00d5cdcfe4612e57f06b40b115bc4f9d8402c06bc74d795f0a57778187641c012a23cada9bf15426d8686beed6016199b0ee299a899eaa9c571899c437e41b233e661a522dfae9f0b13560252465a5b4aa3d231188fe168ca8f0ea7406ed1d56cbd87d51be2c73d93f9a901e6516bce4692fd657f2c11e211c76ea42391a07dc780c38d8f7d6d1beb5bf57d7fe58a0089cd17f2bc566e1401085f1c4be3e2833a324dae33f0b9def502008da6c4408abc312e5e5d7b747e01aabd80d5300cf825d6e585ad448728c0e0fb2f5ad17d0b7b0938c064c1ab4f16cdfd72b4695bbd2d5a95fe5967f241eae6b5e099973bcc4941c81685af74563f80f21a780ef087f5d761417e0d87069ee35d685b4102559f99ae246aab622c7960d0f23872064a4827bd5b76c33dbeff90d9b85db579651a2a00a3e9785c58af98cbb936f1979b6608954d36a86c83aaf7c5424e2fd6d77e6df1291f20ec1a58b94ecc4a611651974bb4a3171cc335cec8f57db1bddd6cda9fe22f31cbac123b3a51a9a8e98fdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5ed0fc1ec3327373461ff2f00b066ee21e93ebc1fc7a971dac8c89ccf9f1289cc6bad5bcc0c6b60140fdb56411ec27adc2df706f97f2107b0171adca573c3e26a1510c71cc1fa34d8c931ce17c46e0633b487043cdb39b984922bc3c6ddfd9311b6485c001d4f9cf4a557929f8b97b0765c6223d26ca8308050b5f2f58a84c730091bab41b570eaab53cdfd5cac307dd37d8c2d9f0213305dceaa8a33b38c33b9cf73eb9abc701c2a627753fedef9de14c0faa6604515ad26c51148a86685438b4111a8e9322d2eb40f49abd72bdb5f5e95d0ffcde81b15b936173365c816b54f9885d6fae36c0624236c1e74c43ac915cec5d4e536da61a9cb44385445ed13d4618b4cdeda2a981f04c650091cf7cc26aa393bb65dfcc92b9ec570cefc5749ffbb58756bc36fe81572dbe8dfa7a5cab71ee4405d0c6c17a6bea5a21413c582acdbbee17357aec33947ac53adccd620b1c02207b5442686ef7d275cdf6b210c71121ec16080c3b5fba369fc7f18329a38c53844a3ebf16439e924bcb747452089cd19b659e152f3f8adeed6cd31ba2d5945d38a4b8670b50bbbac0cd9edf13371cdeb3b132ce000d2c415e67820a21ce6baef97590eb4a14b6ea3700aa91a129d637e6eefead3bd8a7ecc4bbc238e4867e49d57f07ad778c09593294759753dcc5ed1fba41cafdea90dd5f4face7f99c31a256a8db7abfdcc5182810259bf6c78339dd6567b1dbfceb2165bbd7ed72f7c1b987d4c3c3e9721f2a86f1110ecbe449c60c829e32e28150b137eb16bd19021f36a55ddf2e62f11a63c412b5289cb87e80a35bf591a2eb288433a86ba014a28fa12effbabe22e75f9dd19e658d5ae6238d7e4eaa760108f4d84449b359eb6a1125e5638016902104b7124745bb49391b95f1324141e1c5313fb7a25a7cc3ccdeaf6e4c1b03681c08f343d4b26265e53cfbeaaf971ffb8222e2001da00bce77dc561b24a83090a8d3e7853ea7b9477816d701cc7fc6003583111aea0617bb2c8dde47b16e98b4be1c;
        #1
        $finish();
    end
endmodule
