module testbench();
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [26:0] srcsum;
    wire [26:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfbbc88c4d09192db7b28bcd483bca2ac3a7029c06eb5f063adccb1fde6b14cf0036642a3ca83c66dc965bd428178cd7cb14046b86d68c252b6e85a8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd26bc9e6d3818e40bb78b3cd76afb91570e5ce4263d945dbb6f3d5f2c394e6bad267efad69b78740f4c772649f91725b5e728b59609327de9b922f530;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d769378e37c667727cdad3d8f6f5f3e4b3680ded4d056cf7ce4ada892d5186ac95ad3e0b7733f5e7e6579709b353e5fb4acc9793f4c986fb44c46291;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3cb4e2f8e6c29c4d5110341e2d0eee6ec459f537b9e76598451583c546d78ebba70a5ef0f290f30f2e7dcf75d947f1da1a6c55e15d303d5f769a8c33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78ac898eb1739b5492044395d8148253fa0171c2765536a64ded1c29cad2c99a072c0811b386c94b257c31646255bf2964eafb4d9829985597be2d444;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94d5527dcd79db14ec79223f224056403d605f0a12e7bd82e18f3dd21850b22150c52e79a8341a3e25965faf1e67bdfcb53a8b67ee16c1f6469736d2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2502dda52fb28d39b4aea300e116d8a750e0c37f11c6b63a504ebf419ad84ccf27b5e0a68fe5c4e5c66181d450cea273c3df9693f88675bd86c991e9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65c6bf6a88829131fb811201d3e0b26e29a25caee2fa0102fdc52788702870fb69f5c052c2238c2e8c25ada918adbd5c2e1579ec9ffa8526f327066f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h169aa6b462a338c2357def29f977142ee9deecec1bd91c1c1c2c2034908442bd50f2cc727d26bf27aaf41f2a3adcd92b7913faeca1969a07778b461f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56907493228df7e6a28d9d653bbce6d1e6c7f538327013aac0c63d965128ceaeb92c34753d5e9679ebddcbe14ac43dd3dc6d94eeee09636c050a6a025;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4151e179e047e8822ac5798fad6a6d08c451d6f2a7802c2ac308ef5d95b1d6f5f554889b93bcf321c9ab0cfa8a548de352ee6847d88b15ede8e67f428;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5b9e35b8e765a9073695132276bc3b5389507d4b111a294ba0b56a97278d0f9975daccd03be779154f4e67d4d464de8a73d1cc9a4c4f0e2bc5ffb45b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42b2c623bbf826f8f7276ea0b06d7bf90ef970ba632b3d1d5851a37d802d3e03e33c051cf835c05eaae3cc20e59c2e0557cd25b42f1c5790d8b13e2fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87d9af44525187067fe41fd4d0754ad2794ff82b862ad6dfa9eb4e68a6953dcbca0468495aff0f056b18ef5b23f653929a9bae8b7027950582bb7eead;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ec00c100a9e92deb12de21f9ca9ef4afe91ebe16714b33c9a4b14920dc355e9e2316856c8f37f664ddfdc5b47bb780c0116d4c6aa71f5584475b4f5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5f337a6c77b08a374bac65c38e7e6c677bfc97ab09dd869748bebf4e8aa10a56532eae4ce18f77d2d730e04a92c9f9e363def9040788426cd6873fcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b750a579adeae58e4f5387bd4f54608c846d701f62d25e575e8840d5525cee32d6076d39024418de19aa44d65db3d47b10003d4b6693c98a603715c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafa45919ea3038dc8993357c9f1d4571647dab8033b3c665ba9268aa0ea3310ccc310a3c66510ca9f0d4868ed84d4808da816e63ed81fb3ef668600b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5dbfb67d0ea8af7a8c2aec1752014a1166d8d5d3a23453871bae7581a619dcb92fb0f6a129c7c65808a3aebe6e20cbc155728aa6763e585406767e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82ae7f855125efa67dde73d77d4be826c3e41424ef7b22611701ef56c02d7b8198118eea48a023f9aceb633bfadb18f933def34f60d6badc2258fab12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h337b309718bb4c2d7fe15c04400c9eb7c83e9fde501ce6ab054c7633135c9cbac80046f8c5013b0aa4287a8914bc7aba0e3730a92f71e2c8df5126760;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44bd37ffba9a8c74b710783214234db152fe98aa98fcce9da20e630a7e1651d38596594fb492a2d143da79a53ab2bcb540de8961fdf88d57b85b9398a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1de59b5ee3260f14a0c7d0382599e5ce21e641675d40ba6a201e0909d629dff9b4c8a4c1b45611a5ce6d2a1babf4f795f080e0a3c7c0636afe7098969;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h847883f8724a5ba5771e91d47bcc86100ceae7fa291104ea75d3a5a4f01d834c3760d0a045f21bbd53c9f058a1434b8642131eb042db4bbdd05029b30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdac7c6bdea6d7045933578fa13b66773f85a478a3eea33b650a89d33cb5971b3f368bbebc007b3851cb45e6887c9ca4158a57ec55ebaf40ba15bd85d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff408420a33168185e9ffc5575ace2f69075caf4293e420175af34bf0d92c3e93ca01071845f72ac1c0c55be4a24cbd5c7b20e01b52b616006e2fc7df;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdc0aca0539ba6f457dfdb85b33c2cd9e20e49bf50fe351319a782e2e1bb1c652d8fbd77b2c20f4bf59e028ecc758bb20863c16efe102985016d10eb7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7ec2b9166de6f9380815e5688dec0ad43fafb5fbfd02a5e620a800be22d6ca6cd06cfb9781896d0cddbc9a34e8b6cf7b35740b5257da3e1baadb168d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e5868519b025d84e00feb073d69c65a0f2a06f7235a19ee5247dd04e625e256bd14e5d08aad81b1eb406b48aade38641e1ed4d7526f76867332b6043;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2765459485c0b2a8be368c78dfd305159323d980df9d969863c11c6ce46cb27ae00c6423a99ed2903f6338ccc06ff7227d181c1c0fd4027237b24a95e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7486a577e6326774fd21d4b1b260a0c4b336096e8e2999d39b9afa6157065b9b8619bd3810aae626b036e0533744bf97c62576017d482711bbcd4110a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e4ba385ce8dbfe24c7e5090189646319053820c9360aeb1425af128d2f85afd0f5d58bea4e6e19eeedf1e6bf46dbc725ebd310438cbbf20ce70e7e08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3734946a216275f4f42f64cc609b3386ee8261e5f09eb2907833358e322a864ff12d8f0a34561e6b2bd8c1a10932ca5e72b3f82b6343e4cbcaef9fb87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd525e63dfb6c596f3956276ea0e752ba84739526afc4f28e0a5d8a1af2a093209288f310db43c5682a6d9c06c1ae03a728107a27ddf566a469f7bd0c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h370a943163f0933509114de597e62199b64a3240007fcfb1e58e177f8c9206d3feb9c75e52f0424461c8cf4ac20573b89fbdcac81b776e86beba172d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8a697b8d90ec82d6a97be20e7e0d1c04786b35d940855811e60090c0ab22ba9bfaed7bb17e187743ad05563229b437f0c93828d4e057922648bf1534;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h718201152e3c3b66d266d0f8244d238e3a2d257ba87da87f994e5c12f9f4cc55de8796b9ca013bd6ffc2f4f071a17e06721b6f775694110742e431f33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72da38914264f732b64b2b6ded342558f382252425e6559ea9c6a0d81978004c42e33cb5b84683f3cff6a42366289379d04d4805344317e36a193c76b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a70298c8210df3d03fe68eb5a544666e95a17b9016eacfc0be9bcd037b4f365e17108dbdb973808fc5fcf231f7126da110654fedcee5c80eeaab560a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf788675606f59ea60cd1ec0f900e2d452d1f1d9dff7398297e9b20054e169c71e63a4ab615c523872488624dd9422335e21952e2a50cf38bfca9ba88f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50d26b7db5c3251ebd23ba57cf68f85fe03b43b09593ee8535a864485e9e5959dc6210e4ad9d5f57fd57b7949531f6372944c0531f99b5de888470859;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74f5a9571b1e520e0da7252eeab85cfcf80e59009983469c8a7edde8a84b26466cad6a29d4887a66a16dec41d128942a471b8dd17ebcec2b81c7e24ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h138c03b66d8e386d216610d05d4c6ec1754d4956a67520bb71a656f16564cdb2bcb87dd0f0598803bd1adc7ca2e7329fb29e9d2c30eca40ae19cd1d23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h551a5401519914825dc81d2f1bd47d99cce2cd710ba41ad554aaf20c5c289161cbb2643ea74cb941c03ed69d3bbf786f7f4bcc1833f5ea39cd85cdeba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3874644045fc83cab282c8c39770cef42c497a46da1f31ec6ec4719b0cedbf0c9623bfcabfb9ad9fe4dcd6e4e2c021dbfd4aff350e5183b454dd148b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5801a1c84cb12c8bd8b11910f79cb20650c12fa70ad486d4085f5bdc8ec26b5b0fcbbc80f5033ba11f77d63490ebf046783deb5b5755a9b98f6edb1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78385b8ef007eea5cd1dddd8bb51ee186e8ecbd2dacfe0f2a36a96d69977f65cc8a912f7cdd015dab24c3beeec2846aa29380995a2d41941854d62a6b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64826050f425e3849771e17f001f1bd0ba221156ef91584337255fe509e516680d10fb5c20ecb41617ea1edaa5c1dd5414c8276a02443c091f161d51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2001232f1303abb3c7b6f3345ea5af03c83d9b3b70b5b4e3ae59f3b02243342ba08b76b23f6c4f40681e051ec32efc7b23839c839153832cd9bd16ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h468e9a00160ef77f30c80f8928708909da2c159b0ab8fc7b146d476b0ff7bc2664da8a2f0f65202242d80b6f9872d9b3218fd1e9bde2d8e76f3ac823d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8160f692df2e20e1d6b63964f424c8e992d43687a5244e83a84123cb532aaaca807cb4cf1e174a18b0961fed4e9bd1ba70d4efb4a4c21e22796118b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0cc045a895ac239712798c9626e3e4f4a3161c3109f750d6f00b62d471afe1263d88ec2f741fe06e88a655dec1ed5076a188884caca29a31392a5bee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1db3c8e15a7ac931c36761f1e8ed8adfa040c6835cbdcc7537b81890097be17b8b6d74691ec3aeadf2316985bdd2543c2f72551fc4f32cc89c8bb2f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15e216c70d4ae68d06b2c16aa989fa4acacdfa68fa807470589ccfafe0ea005a028b450a69571e006cc643f9789dbbe96a7e8438decca8170c791b0ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cf5d603b1e28210747a02221e80e1f41d31a89a1248d0c10f1ea96c9929d67f06bb009352958ef3109c670dc5bd34ec0f338faf022cdadf40339fd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5749733830cfe0b36ab6bf3b45807e96aa6041e51ad5cd092f100e55d4fbac82efa1e98d8adc3bb605732aa1eb9090cd1aa13dc43b73f7a74dbf34c8e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h136edb4b8adfcc9741c01b72f71f9cff1061431beba8c7283484c724fdc9fb129aac1719a410ec86e5d98ab93f938ffdded29b2a7f7bf85cc4339ad6e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdee277b7090118df957d4fcb54e3fba58ca8ef88b4c57970e4bb69f90b10f2958edb3af5c816dec5d366c6472a71bb92106b47085b569d64f75af63af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb25dcf9523f8d392ecb027d7cf448afac87f6d66c5b47ae0220c512bc9195881111b0b8d1f8f38a25f5faec6fb1ae923b05d933ee20a5fc942a90c737;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25c4fab70c08468fe2eecbf07a44ff6d7b2528c1982e93f7367181bbac3b04d5c01f705d83f4fe31972855dfe60545a1343fef425873f577fb167295b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9318b01c4b42c6644d54001536be809d40640061a07804f7767c24214bc8c44aacf0db44a4feded09deb644a5117c97e896d720357cf2659f8e18b565;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc431aab457d438363cd15e277b70cd20fe748637ac17b287b7e18329a79edb10c3821c90be81af5cd6b86482fcb2aad428c6e220de21b5948716b572a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b39c9caf1e83edb3ea383882b785d696360845cb289043221c2dd903392519f5b807ffe053bcf3f2c557050b91c9101e986846398f00fa005e5e2d75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d272ec8e88c195450f05a8d4e16474c8d44e2514ce9a08d36d66e7808a5f22fce0532d0372f13e4c6399cd1612444c238b52c2478d8144215383e7e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bb2474578a88eeadd4626f951d1197ae65ab0bad9344a0d9f6ce173c2d2d36aaf5f0b729b87e7f8acdcf2a30f8817fefeeebd8f496a95e5a81e8b8dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47f6b6e9de09c0c58b20aa24f8f92d1df0ccf99ce15103ede3453d242a38e7317aac7b4150faadc76d21d97582808a565b59ab110c8dc57f4eaf181af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54d7546e822a48737fb31527bbd88791ea64f3508edf82aab4c478f0ccaad2f5a4f35134899a63ad1c9ae5f89fd04658d676d7de254ca4412c2284ba4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bdd3fe8d21baf513839e51fef5148de755a02860c84814a8f3d1c4cf11d7704de1dd08291a79cc8a78972e29843c86e7e95446bad44e7af8b3b0ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc328e00b5e94c8c61370ee9fa87ba8d1ede30d0d277080754430ca7b8fdbf33f836fada68c1d2f6555cb0d6fc45a0134256e334b24db44caff4e09132;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h360b2ad0b7e80988b178483a7902db348b3e86142a134b4a3ef1f55471885ca47ca669ee12b1859a8469ceb6c2140748a7f210b62022e8d2081c03cf9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4e463f6b0890b17e2fa3027dab275dd5e39c20845d5aecc57141b33e8e5fddb69b24203ce22b15ae6bf50d84cc49571f818fab406d22411907dd5992;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h903b1c856602909c5dbb7e9b807c35357350d3c5eb7dd9446e195a7f7d97d6c19bd2e7d239d3ebe80d58190622c5a21b7d7bb374a2aaaa6a7e338499e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9a7fe0c32edb410a69180836f4a41568d2ea53451003383849ad4d8ff80571be5924de84f26c76eb3ccaab59bf47bb517baefcf8d629ef9cde71412;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d5336f1e38749a181c7392f3803cefc507f7550ae1c7d3c355a416cd8082569065c2713b41ca837859e7dccad3727215e2430654923b9740875fc9d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9007e9c21e9db3b3779b28cc2dd67f211481dc767209f00ca8b6e36001f02800bc38ae213196f5679dc36bb8911b2654e356d4968049d1da0bcb07;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3afe5afa0a3288a5c7294b8820d3a5a62cbad4f1e292f39c3c1b6fb73fa2dc4807d0930e328377f113f191b798f38cc8a068cd52d7d0864aaaccb1297;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59dcdd3a765dee7f2a8897cffe4e64adda8790cfe36bb986b20c713f0ed1b623633d056c0468d6fdb8e97aee5ef14b2621c6565e3062770d313d3139;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd4653a4f38c1dca41224c7deb11f7a5b6bac5ababf762e78b8e3de26b4707fb8ebff7f440b3735edff4936002f356b63d2edd5c843ec4e3bf58018c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8bd38a64a9fe4a1e92067d4e2cb9287d390a7d87aac779e68903325c5134b1eb051b700cc0d465e4490ce037a834ea0ddb7f26f94bacfde21ccf666b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13aec79c2912b74cae057a4a2c7bd2651f4248c16024b89c2a1ee5602a8b46cafe164115495743595c4b4f14052ce45dbbc5548b1b9f905249640b2fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bad1f3eb5d9e593b86890ff28f8e4b5a2da0ab136266d8f8840b3889127b776717fe0c2f87c7267078e32204b2f2bf3998655d0cedc6b4f4c5a16f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4470b7728a5e1c78e235d89eee9277f7d190c4cb0da6c6bd4cdf48720d0e9d850c603d43dd74630bb70260cd06eb87f74e6d6bc1e69cacf087325dfb7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0762e5396d216aa9d8ea9bb98c49db05f7a0f9b0214ad44e2c307e2fc1838b8b4052740b188c4deafb6d402724a02ca9929875d083bc91e49c975e76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfad205f86d11040290101ac33ea819c75aef437a8c84c7167c6b49ab50493025be36a2ffa72d9a0a618d6334b6da8c3fce80ae017da8d02ec57ea15ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdeb705792aebfd8c40635a2e9e2f43a563622d4aed17691ebb22804a1c73879532b6ee7878591c7db0c2d23e7b4dd3e2930b6c18ad46bb8e468bd65f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12ec11fd1a98117bedf6d340747934466d7bfcd766dcf07fe75e7e01a4635d6ab457c88067c36ae7fd730dbd369decfe73ed81dec9426588ece1ffc74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34d1ab1d1cea9965bed48eb53e69089e47f328a6160c5d45b373ce8caef2e9bb89d80544ba5c673b663638608fce89cd4353ee6b17804d47e1aed0aff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33495db2b604c7b6d075bd1cb01470b488490e55af910d3374688e2279a50c00f8cf7738cc0d99dc3a471782df60e523dd933b0d3622bde2400aad20f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4737d83c7c12868c2ddbbb9c37ac48a0ea4d1c9700bfa5c6da11f97dcb7860a9a2989bf2aa596874c61d478501f6432d6b52c5ff3721f8f0e87bb5cd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56cec3759d19f162587ed03fbee931c24da7ae35dd51fcecd5545296f0240e92c88062d7a660d02c9e961fb648014e1ba5f7f24cf977434abebab0f40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24f81d756bfa87952c1e9760da9de8dc1ccf291d5def6f54e1f5184c6770dfd941e61758e75ac8d80cef81e798d7a0ba2fb69b88dd158b3401f91102f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f244db0cbfa7a128232f4bb3ecb7e13c03a065d8ee8b0d49fcb9b7923f893339a8a245d5b1fbf5cfc904f51137cc402c7a67820e600b73b905364a08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h773a737478f98d333299729426fb5d18195628cbd60fa7f0134dc91270202702f2d29a8b895b7921e37aa133b66be6e44c5493d106f7b7281629adda2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haec5374b99fe0fc1e9d4dc471efa78a638d6752b089803bb2378b75d97972e7f7a23acdd2b3232b19d9c913b8d5d86234fc2e24eb002a81102e231543;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e81a90ac52438ee3829bddd85041effb91f92dedbc38ef5184436b1b7915b028a79e951a38f5865341f46b43e4001fc3c4edecf3dea67b1bb41d00a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ce31c83e4972f8ae556dbd8be2da5369641fec8fd88666cbb1dcfba76cf7388c7d9cdfa98321751e03d5c4de7623a973a5aedd2a36014a17b066925c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h553d7493020530389aba8a8b9eb0611429c8c2cb565c4f50d2e0de3219137ef9ff87814712652b6650fd1b5ca4cd7fc2325a817391574b7b1c93155fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7945b8973747ca82b3b58079ffb4b337b4b564f3b78dd71b482af9da6907c0ccad58289600b12c85e4046be2a49e3c871d1f551e1cdf52713d976147;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd21610730f7487de33ffc3164a4d609e7b71e213cd096337a0d5d068d8808685c9a908561c93246fe47c2d1aaf48d125c55d00fe24f6083b4a1546929;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e9c5324b20c8385e30da2ce6fe3c1da882c2521a69dba965375922d169637b8f64f3b6e6261efd49c53747710b588087a14cc1b3de12b2fc09dc76f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54311a19d221de6a73d3c598b32338bee23f48f7c0360e46918266f2932b06d10b9280eb5a64eddfccc11a0ebe0f52201e9494cce176bd121b15394b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d30a88868399e9c74936d0559469d48da637ee9dfc2467eba1790cd3d76d0528c1db1b6c8e0f080a31d08ff256dd450c88c0b38b5fe4b146752e90ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bb9b5c6fce3a85b8c6f56067e8a85690e7ad725642b477948860af52d8988a3bbb00cd824dae526b3dfd317f773535d98ea92c8f8bb0c00c01cbe4af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c3d126ecfbcdc55d973a34594fa90cd452b1d129338e2266b3fd8f50048a00f930f5b38eba00917c812071378c601ff568454cf269688f7b7a24bf5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7e14cd0f33e85b7d9b6dab00eb3b09981859307e5516e0e792df88039dcfc814d37bd219cd4de5d8e24b1dda5d4bfdaba4e74903c15e1c0fec8621eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6fc25786c41fdcaace7119db937d6f611b340055e972431eeb87c7d4970e4e22bc5e01f6154ca69c7e8ab04fb4a11eb88f890c8ccfc2b5b8a9dc97ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h184f4d0bc4206e4cfc3c1242e62539a15213eacf2617cc3f36bb3286f5ad65f127c9883faf8ffffe992065ab08ab2be4cc676289a7d9a237554a6664b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he48d3fae2d58f7f51d5ffa99d7872a3e47d849a969205d872f1776feea39741f8288633031aea45e2dfa0fa1687fde80ebaed7c38daa4545013f2ad67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfa3a7858a8f586632c7d406f88868508605dc2b8e5e6a0aea8447d5372a8636a25a3bf694ec6310c69fa5d11ed5e64c975f6c1ed480f0f4e145be448;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a7dfc3aab1011091367353358841697f13f433cd9547b1e25ae2c7595507d8c4f909bbb2d9b880851d18fb3841bacef9b3e1d778afb6482561ddb30c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36ae23b95af3dd25d6336664a480089a510a0501d66a6e230e3cc29f1d24f3b577763b730201fc45bdf77e8a7f03eb81d5fb89afd441250dd1a56775e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc67c4ec756f193d840e402f7cdcfe692ca67fe10c0931c3671ea53be06d63a3793f5d6cde263ce09bc00b05bbe19aae197a7f8193371790e52b425f2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h771bcced9a7780dbb5191df9ed8b2b94ff1037a67d8f8028d6585a3729df8cd8ce9d1964549ce3a15b71eda69c2cf127e84edb8cc83fa64d51a0d4522;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb77f5d0e1bdfac3961cac6642af63cd87ee76504076edbe89a171cebf007b3c0c278752a96a0862c9d1bd9548f676f7c5fdc5088227f028123aabe0ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h111f0c135c5eb6ee61643d3113c65a8b3f1bbb403bb78540096683217d12c6c5cd113aa32e2eb54bbd4c6fa5362dca907692c113a0625de10adda3ac7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f2048140dfd7b94a59a6264dfb60974845bd69f1ccef533a654b65cc366ef6b8750152840f5c2dff41a04549302e5a96c4b88e554a2115536faafc9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h385cf9321f5d229dad9ed563865487fc0220501b38c96558a00d686d13c4add04a6b5e88df0f5ea10cdc65baa54787650a4a58ef4391c60efbf7b3d9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd35d259f9987caf8b2994c8f56b39b8e18263c333026b3f5b4b4181241a809d83bab1fdadbdcdb9c3c8ee263241b8fb9091228ee0ba141cab28767db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4573d846a98fda43b359eab56c4b87e796b8bb83e16623c1c57e338b6397e8e74965343466e61fe15e3851230f616c78dc4f8f8a488db6e686bbccc91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6802d5fadfea08847d502c2b91138521beffb349d0d8fe447012358bf93b02c3aff8ef4294ff8c17eab6c111ff8e4ace992f065b7cdd557899746cd75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5599d5cfcd055266d8146a93a08592bdef38a9bc1ade2a6f9c933e156dda33f967c945dea363c37c336366f94e1e2464b9f9a66ec5e355b758b862570;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h607c1d3ae37a5977435148eb1456a647352cec115efb769d73573525ccdf81aa67dd76b326b8793054acad1aa31f0fdae0a28bbdf16614766466b1416;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4514f02d91bfba0482734097bd44c920196f8f0271e1840cb220822f185e9e2293080d1a58ce13e7847c86c1c8ab57e3a7202dfb88824b91499c17f69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87883da503ff8db858dd488bb50adfb38172615f0769da1127847fef230a1e2d07274fb1da681a905b1f4233b77dbabd8fb2fdb472fa01ee79c81eed1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1ea3e59f714cbf5e30dc73b9484fa833b71da1c6d26c5761db7623dbccc01213f8d7e6136b9b5ea131ce67dec8dffcf837a61e3a3917980cceaf658f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5faf8f1c61827db95464e43ca780ed91cfaf2a3d8fc83807ec82539eaaf266d1c8af37e5d39796ecdebf4b3de335778b3f6ecf86932eafe2be54611e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56072f11eb4edf51afd6e6356851132a3a0641573d6e77978517c8f82daa4aeca4e19da8e4d07fc80e30ba744ce3dc54e1e3f3829b0f9c7aeca640da3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h439276c7b4fb811c430c2f16da6711d07d961de0541b0c7b4a4b9b9c06816e19f6a74095fb7a47a16ebd72a5342fcb4cf6fdca6761bac9c3cba4920a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ee759f2556faebf14f1df4fb120421202fe9740782a82b70d83ac988901a1b12b3cd517d23c3381c184f8e4a464d027b646ec2f98fd70c866a030785;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0c7ce5afe90d8d81bce57c406a38d03288309eea02f87df85411a8678f6fd546745ad8c893d001785b261179678834e7472a9e67d0ffb1e12d8c97cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8239a128b3094aacb1c986111b687e3d5ac984da2be80ace03ea9da3476b208ebb1fc8d3ef3595c65904c58124a1ebf68e6aa445722f63781504e3b89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcadee83e965df3269aee275ece13fe64cbb33c77e686ce2fd86ec29512e1c2565bcf69ca93f48ed514e6bde1b9f811b3eee31c92c8f4f578c89514a9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6efe1df89423436d006282cb3e6db222eb49a00b3b0696a24c59792a61f4051616d8ae8183659ec75f0ec9d6b6e43c2117952f444ff7eb86e9bce8a90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4459355a8b2f62e601c50a4265b69c87084c3749d02121a7213cd59f0a576b9d4c9028da5a6decbc96bc84cf49c18d1c658402abf1d9575423b04c08c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2d47574343364f821d7cceb69eb448314cd6e6882877c978d7b0e3e788e3ad6ccf3f22dec6a76b30d4edf2e8267ae4a2e8b6287b3107c05d0aa26250;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf4181a60468a464afc489677fe243b9de0f1fc9e516655b0826cf49c27132cef03950e326405dc3067bb90b3e4e8f887740ea27c1eb3cd208fb1c019;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43786cc458bf007762df7646b3aca158e346482b341c2c42883bdfdb92cf1eec82872451ffa55a9a388aa0bec7b71014b5b5345b99aa76f7f8983e0a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5d8009693acb026abd57e6bfea6a17ae681398c795734e5d67356bfda7414bc81657a03d33c6f3d3de6fb9ab212ab279105329435ba833e32fb4d121;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h675178fa6790fbd4361a08f79725c0b2753f82784e33fdcabfb60573a00feab33b12844e4995794e2e86d2c5363ddbaff66773b4b97cffc5634364856;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d1e30254a30199cbbb3274cf2acafacc994bca174d18124c38540967d5be90c9322a41d63a7345a962e4465bfbee51bdc6e7e0fd3406946ca1723f02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58100f7ebba68a6c2293b1ceb31502a440c3eea79f89570feaacd450933ee9f4d65de74112bdd015a801aac43ad625a30b62371da93fca08b2400b521;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbca3a119468bd0f722d9ebfc9687c4d6f28e015ee23837f7002e58a47c6768ee8db0bab51f96a7971eee308f23bfdc3976720fffeb6b20f25c6810145;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f54ba2054f3f878a12c74e5df6c0a6f2a2e7d74593b1bca010260ec1e9061791cbd7337892c16d7d5e3420631ff1f4f1158ab7e4b6c67235563d6e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1134a7e690683dbf6e345f03417a942f373f855b2a924617bad88fb6a7ca8763d7abd4781219676da74fff9be1080a4bc969023d068025c87c4a98941;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2156e5289cb7841be3e00c5d080757e21c2e1c5e758250a36e9a71053aceb0a50f5bb8b5176c3ebf7c9a859116557e09fe1d5a0885b1dbeca2a34f89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he761efbd1a5321a6a23542bd8df3fa9136df718ef3a29e28349463b3f946284f4a5802c688ae670959849705279b1d1f5380140bcac239b4092970c98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ec7b5ed06087f842f5e44a57d2b0a0a9a8fadb3b9ca7b5a34b7cf5c4e5d2f5dc50208506edca472189e578d624c14da32142fc0c26907f70ad1f6627;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96251ba65b52b069d814046d9074e5122789f71613e73d43a4aabe3a12d5a20b2dadd8f2e488185db0e3c53efc2dfae11d24c67def31c4778dbaded22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e43be92438936de88cee93afe5616906c0c6496e7ff20138b860e0c003d1bead5b8e3ce3dfce3e9cdc3a3cb93a7935ec8927edd760b0b359fdf55fdb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ed3530cefaa853e87993319aa39109cb58d929139d88a1656b9bb0b78fbf7b1fd3718711747ef0eee54f364013fe00e11fe178b5c6b032cad2a7546f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h876b0682a90e81432170301a5ffe61f6a55cb294ae5978604d58ea862aa89c29c3d6f156035297828b1cf1015d70a64cf65812bf9b471537f1a74acd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17b3faedeeca6461359a0e2e407161a5f85cb67169c47b93496f64aa27679a319ff9f3151f95e18c331452306be1a5ce4614865667bb44594b2495a7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf96e4eed43c90b1f13aaa936634745d945ebb66793b042dfb0b86a93f4c09600911295027c9fb6b3bfeda61fe7604dc2096eea9ad56cd6b1103e95543;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd86c5360bdfa16fb17e51613b91e2a75a6690aad58b2a396e0a411f8761dcb5552f4a9fc7a4d734e0d69a97b829db7466579e4e9d8e55eebf9b71dbcc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha22401d40633c7428a1c1ebd0664e7fd3db86763a97ab25d2d2490a37a816db56764e45914c2c2ae7bc20e5d97ee0ba0e338118b6f2f38c297b0b8bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47f3003f2278da10da8dda573921b10df1bc3df717da1a51cbfe0cda5ec7fa99041ad3f9f19d0d43d99498cf5af54051efe5fec6c6a290c35ae4254ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcc3b72cca46ec982c048fc70fa9e3edbf13a1a6867942691251fa1a075c28b750bccf2e312308d7a28850e26712e2c09fff16ea9868d3200569d6e20;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha52b4575d1a2c7dece5f0eb11dbd5a635808e78eb4cf61b2d70e5295eea3e8c99be9b90b1ba94badbf6505e6489f34a88040cf4a8db6051b089107af0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8593342fb26ab97211fbd2fc1e8263ed301ac40ebd852d234242afe2d66d95efd23426fa19f8b2182aab489de421316539a6c3ff194e3be804eb9d77c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc478c8ef98bb3d5a6fa70a43928a0f6626b7e2664f673b5089c82e62631785f7a87b121ea0b1fd204b1cf81749f0eec1886a65b77f837397ce005545;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h284f57e41fa301b39ac59ea3f751084ea4fa2ca4b268a0b22193628bba7dbe8a38cb3526f9c3862fe45b465d740f0231cebe80477df01ae948ce580f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3e3f647f1cb8f5ad59ecd770c008c7d059d19eb916db4e88b7fdd2d7e3ef8295d629e9f594213bf403db42793d97aa130982ee80de7471206a775620;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h433905de522ff517032cd20c09226722407b0be66e431f0f111f304f5802f8875c25b11def2ec32709e1721b4054d274e68b515e1d25a8c75643829ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb34e43f084d76d836d2956ddbe4d97b096c7f7dcd1c8f7e38d82cf157485035336fb1c35f6d9b93ed52f5a5156eb702a0edf27ff0df2760893af95a07;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda69471309ad0e142dca85360f1da2f9dfb2611477678940af5e7014f2d39e299615c5a7ca502898093bf8959d8ee216881c5eb3469f8b00fef1526b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf50782825c8706dbd8a66c0f5b11abf055b61bb6ae52ca8f09a449e8cc21dd567d1a97e1d6d252221492855dcbde7b6b6173aa68f3d20329e6ecec9e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e4ec6c56c75d6573bc00df9dc79b58537e9f2fdfa68434f20fc18c9db3c4d2cd5950822d2df7eb4b1d84834ced5b579134490ff92fece274d846f289;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7858c44b0faa9c63b4422b2676259762a5839723a2b44822bff94157ba8adc6f472ae766235392c23fb3069ddc380deb5ecb4bed1ae4fc4aa6e5f6e39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f744a987f402d10e906fed32d795333e4ed446e9a1d13397056a05f4800a34647d4513c2bcd5893f01a4338640c9a0fa5f4bae20df0e58eb569c5823;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d95f9ea9ec0bb8e7f00a5b0b64a232c3c2f8a3b79268b627e8eca9c2d96acc99ce66793c5a8ee70cf2da5b727d42018c662dd2dfdc5f44b8490ac112;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97b2330d1fb0a05872c94fc66dc099e22e1e733385d69bde79294aa91db97a9606033d985a2bf58e8aaa31decc3f0dae70f71766a5a733e93cf7a0475;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5f0bd73bff670934f220e1eba9c934079407b3c5661f02658e3dc31f0607afa96711cdbb2fdd46928c2c34cf7efaf80166fdf935cdd17c052cf5f559;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4287e646b86f78c36da94213cda5223ec1a38171cbb06a92384f75d4d4d2c64352653ebcd05b6c2ae5da6f0fbdda87de02581a02dd2945982810b8ac6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3fba0b550d3c55f48391cdec113a2ce2847f89331c1015452be51a1e96697dbea788c8a828660e32c166c53da718b1a2211290ac690adbe5def9613a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f7c9835130be851131a91e3b6eaac5384a6568f900e8dde68264c1f7c5cbc51cf568f3b06d7e4994a81143ea8d5c6b3f1097ef28d03b497f6a3395ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17bd242c812150290a7d6a91a160a8029cfded4ac435c76a409174ac425ae9121f6a284346fce0317241bd8427d450625623df8d1fc38cf0b5707e09d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b9135eab3e071fa21b8134de37415870a81817220dab1fa845b2adeefdea9181d6239bc9c2f2f2d43891c368c85cc3b86241abdba1386e6f55722a64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd597c01adaf67f7c3483e999ca8aec6b8b1b91243794f2a31ae1d83c050eae3fc2b11599768c824a5c2f88d529bc418b0bd8ea7e6fdebcda36c7937c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbaee693842a41cdc25ac035cd2c0acd005d994bd7a2c4d347152bd73bcf2c7b9c3c140f1205b16bc651fa6495d9409e48c5b441282abdaa56f14f5fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb56e22ab4d1a226c644b9b033d4b463eb3da3f6aea45a8a46fa74c2e8c4cc689b45230cea8361f40b5f5ebdc248be2cead38fc134b675bc4ce8a1152;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he986b0d9c97fb7c5d3caf4964b009bb54e0b71be0478759f2170683b3fac67d2daf0b27f3919b8eda9ebdca9eb7b04e348dca03da82653a24b50c371b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa0b1c5fd73d4af6d46ecb5e688fac315fd1c1109158b1eae80c49ae5dcd5e94f2f48870de3ec0009c014ff0a42b0ea204660bb8025c708147941d1b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bfa3e5411282def5cccb0108423c87f2750d7c3a8de374459889c8a26c2002894605b77800c20b12f869e52f5ae49c213fa1022bbea867ef1e59ca19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccefde2f07e329b4c893d8d622b8a879b83bed25732ba1ee694c7ffd0bb4b3e202452d31ab9e5decc068bccf493ec4134ac8495a6a1dd47c1e2e72de0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62999867426da7243f39e3371970a2d2069c5b3bff5f014e6a7aee6ae7324a74cae9de331850351dc65b7775b39242cad714f84be40d87a25a35b3ca2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc43e957a3570becd7290bd9c11cc14d472d973fefddd0c20551e0bfb0e2b5a4c7ce5c593aff3720ad1ce00c22ae85bd195141fc6f2440894344541ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61e1c22625e7d799a9783c361cba842fccc86932168aebc2792fd9e1b6c9d91d6ff83b9f2944190d96e489a4450c75437da238c3b2ac0746a2cd85067;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5a8313416c25fb03734f84778f00d9d67743383c1f1c45fa5b2e0a31b43b6923123940d4d0dced82cc3d797dbd6d956473a3540863120391d4424919;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86ea44bb405d8d4de58f9c6382c93e6cc5d38f7c89f78f5eba69f40e8095cb7c6e736e15d610db19c9b2b7ed63c3f4cea0e20458797a892e405aebd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h959e30169a9efaecf8c07c02db99e6dbb4d6996e9dd030029e14e0b5cd96e9e7676645f5c9313297033f2855dcda394493c57935d8dd3019b08fa9eb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h432b92214e192e6404316d33be89db5f65f5309941ac2d97ef6a52b4edc628f3a8e5a3fd5d59853a570d907154eabb551f093c94adc772a3df2b9b10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbd26f55bd31583bcee81c02cd93b1e580cb6dc07f1eb3d2047fc196341185a80766fa42f8e5aff10a3ae93deda9e187ecca53a43edc754d985524821;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h801ff6559b7f8aee0582ec304b5481b08d650b57078809f5ff6ab879a50eee4a4716dd5b119ed85062d0395a10664e36a9d05a6d1a55d688d6dd224ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8dc01c4c1752f58752c99ea4159fb994be57c4e92c062dd8d114f66019be3a5f10ccea1dd5e26d224b8dc9da4e6b85c53f5be9b13384d8c8f730db89b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h747db340747f748ee0ce321588edd3d49fe06576c66f362bb3a297db0fa350eb1555bc71305ed35651f2406daf27f197b7ad213083ca8c1713eb61385;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e5bb27acd9355eb1202a9b30e55268ae63e7c47c9af3d92f7045dbcd9380fa0ce55e3ad70dc9f4db9db18fbf6acf7419e050aa95a7c9dc0d4b0cf686;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9b3529a10ee56e774641ae9f67a857a0c7d861d9f4b0ba48a9caacc94ee9cc7fd093c76bc8321a8344dd5b7e042dd7f294fa5b4a9e4a1de618b47f1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a6f0846f8a436c73da3d685d56b1b9adbafbb42a81763676c5c09b2d562ef53db2cdc6acf1aa2c8fb959f69ea530c96bf1a532339e6189450c8e4c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51c419d2850e1b929bdf43cfbbc6bdeee572d9342d15a886cc1099814d55906fc1ebe76c1cf9ea5c7d060335117bdfc86b76f582fe3dec68236bccca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1f48047d74ba4111c1b8767ceb265d0615c2b89e35383b21aa19dc89c97ca6bed0397b9cf4a9e421b84608f82015f571df0ce8a5d44635f33d34a541;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c6a0886a6cf85edc83ed78411de87e7028f3ee2c169a86331d14e9c84b404f337f96c5b6f482c326deb9e2028f29a1ed3a3c64fcf545936a97e173f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99d5e81aa8ed6dd41262e346e0f2dccc189ee513ffb5bc8c622b95012da957c1b923317a83f39f436bf1688f482704ebcec29b84e995f2b766ffde5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha92d653a31f55ac0f76b7fd654f494a5776d4a3042a088d94a60f96e7c4f40c52c3ace70c925b0c40ad8aa7687c1aee7d90a7826ed22f3e86433dc685;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h528f61e8df1bc7fbc7c0fb87f61882642cc4142ecc3e5c3476cefc051f7d46acb7f01590766e28ffe04212689460d28388988fd0c9018aede3859dc4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1983b0442727a7c37620e9b4147b492e378dba7d984fd5f6656aee0f9baadf77872c114c83c2a1a981072746ffec9448e83a1d572385ac0ad9e88b178;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfd47a2aeb6dcf589e91d95c521b98eb37caa308e15648d6d9097dbc5598e710ae55c45f0b4ee48494dd9d13bf3324c20497edcfb72cc45bd9ada083c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4efca4cb8d21dcd69ace1a922e11836a18403467c552c03cefb21047e4dc394cfaa92e6f144d1df6993c8818638b74348abd6d8cf6aa818f23e477867;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb921b447f4abb85c9252e15f8e4eb7e05a9faedb8d4235ffb2aa1784bc77675567406c06911c8f44d72db5fc510218bf1139ff9fd29aac8ede28cd5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h376a9c594e1c4280a297bfca6cf3c667268e0085d2beebe47a962d216be456185c145d3a009a1ab615f9b281a381b9741aeee21211971fca3b3732792;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bfd49358303cf07e9e10c904e1cc548156299695d622f0af5e59de97109ece8b67f2d79d2047a59b59ab680d9127380e09f654052a10000440ccb769;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a6becd1a656589b2fe0669d180664173b783ca6ba29d8632f9f1fe9c25e68122b02775b42bc4e58a20ecbec8b2a1f89b96a7c8156dee64afae58c861;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64fcb10a4b9f76312750eac7e973fa6931397472cf6364a3ec320c5d753cd5fe3f175908d24eb50ebaa986b575b9ff666620a26420b4dd049b4e6386;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf302a93f7cfbd031aff489b7c36330a3b9adc8274f9c6a58129d18897e3f43102c80eaff5cdd125ab3faf236bb1af46114b9d1652241e2f42bcdc793;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94d7851be3cc447420c4309472438688639122fd8a02d0c0f394ee5a44fcc051899414171590a386e3605245ac4e52d9b98ccffbe3f4e7801f67bbe0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc982a63aa166c9515ef9fa099598be361fd8a46e0832400913d100bf314e71285ba95080f53149332bdab883aab2a6cf633d22a6b92c7f3091b201b82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f682e612c708b5788cfab7861bf80de2dd53748a38f90cf19e786081003eea72ad70b7ef5fd9fbc9f1dd43f08376dcc7e1be1585f807f94de667590;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf49e352006a2e67a6149fb47425e9b9dde5c85c71ea42d505974aabae36ea6e656733c91863184f91c2fae3a9b5199fbd74861eed0b66bfad1e7f0f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdc0a70ff9c04fba15e0cb312e14d2f5abf711ede79f0b9cb7d002d4cb64cc72ba81f4ff8911945e1a8fcac7d5529bbdf89fe958682fb492f91c96e7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb566d842f151d85f1d142c63515a113aa63060d567c811ad2fb1cbf9ea498218f96c852e560b4fad9c9d7d1407b85ee5f65ff3d7b9b8ae24fdaa678c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h908323d53470b6636577dfc032f546597244dba8bf7aeeceb92b40bf55b9aa028627ef906368a3abe6c5ffd1717c9ec81a571b1c777feccb6970c8c98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5bb5994dc38d219c8bd8eedcf63f746e387363753d8f71259e18dc46ebe375cb1aab867864121b53ad2762b36160f82536b552921d25fe7f6e712fd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4d64f4596788484d1756f22bf9998381e6e5300f89fb0e0da73fcda29b701c723eac1da69119c104b16d5aafb0342eda74668a262e404036ce85b5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf43f02cb67a154497a0f19bbc6c908344ea80104081a150d80000b310e25f4c3a7e9faed13691ec3ec2740b35f332448379319693855040486f405b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49267b922a531957e186af7efe39bf317b35b112e1a15778d288d5a2da450c97cf7d04d4f1dde00b70797736cbb8ab377f2fd6ee669d5aa40c598f59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heacc897d90e04c2a6904269bc3ef34c8c5776caaadb5011cf7be8fb3d680b6c9dcbda80766ef2bed485a28ac5d7cc73af3e252f088cb8b5c67bf30bd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8293a4ed908ef0fcff9eb6a0d2d3f34d3ccea4e0ed5e23a5f4d3d2e514eb045776a7aa8bbeb9ff116a126fe279652563c4d8a8cff655cf662ebc46d44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc73bde0eb08b865c00b0f17d4ceca76ec6046b1595a5ed342ec1438223fdf466b9f8b9f502f50306958b5e6399c3495545f1197a992f65f59673c335;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c66e05d1472dd322d95c911f95c4cc5d02ed3bbbe70e9d4624332b962c34488898c8dea0e75296094aa4641e314e73c1ffbd223eef4d560607b735d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd037da4d7b02b67aa4d610685b0604e6b9a33786933c548d7079086a65f02e41b7935dabd490fdc6eb3930595a79794a03eeb3795af79c61c4766dda5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h549ff5d4df16632a5a3df9b918cbf6b747ef80036035a92559ed1e2ea9644bc0cabb9cd11e0e8248fc5b2bfdd8ab150dd191505409df7927ef9207726;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9a86aa00bce091a095911262b633005de11559c91f8e3e089134a4b57316c89012986911c7e23d19b361de4ac11653e864a39eabccaa11d93ac6f694;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26ae7fbd5ff67f932ed14d6190c8cd58bbabb51646fc66428a58781db4c17716fd9fb9189faa27027e0e7779322899979f3f8a7732f7b4831a390fdc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1144b795a9d78f3f928d5741d70d68c5e74c9f819ca73315c51af24690b49c6ada20df6e280c8ce8722a6f019285bff7a80819fcc9f0f75f0995e9bea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd560922420fc0f9e44ca14274359c921c56451c51dc4309800e039a7b46a62b7945ff3ea23676e9f571ed117a7e7cb98c9d0947c837e85526c0e74b75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h143eed194a6c1cc08b528ff45e7bdeb94c87aa6f5997742a3336db9372c8401c4ebf5c994be5a44afe8bc59cdb39ce5bd6fe2dba49240e28d391663ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf49ee0062595bc33df0db3188a311690391709b88d23bc48788118a1c1103c532b7423d2dc591c1bc6b313a055b9fb3444cdc30e55b219fe2be25c1ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf19792b2b5f8b37b9bdcd2d05319add2cdbbc2ef02252c12ce72d3cb4021231f3dd28061acc19e4164b8c063236ef472f1e8c905b1409914a2aa99796;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbd5de165e0726a9ad6255e4715a04e1bb65c92b609c169f352be4c9c7e8d6dc2a18b8cbf4303e61e82608bd8da30e9c3e23c3023149ce764b87f0ea9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72e5f3fb17d4d016ff27c20787bfc27a7cf8d00ae59519e670b906fa68487bafac3f224e856948c15eaf7a7abb2cc48f10645b7fbd22bd8bebaf4a976;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6afd3b34f2b09403979773dab14395b99a67bc4186221dd54b44bb84dc8a8c77a02f3ebc06f9f85ab5d4ca4c2622b7d4a67849628a7d258ad8192e3f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdc0baeaccc81927072f0748d0111db413ab44e8a86ac76ab8b32381ceddb8c4e044c8f562ee3ac47ef5ade1ce44635afcb66dc7f09a6c09a00ea47c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1f14465e55252aeaab26b3ef4c3db58a586baee9161a46d037bb0d5784c6d2f3951cd616078ed06a8d802311f88ecc63c1a2c90370bcbe7776aa08d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha94ec9fd8bb863008981688ff9a40c894bef708343ce69e2b4b3b134e4ebb2059ee5928873757a2bcab451a4397705840dedb4c77c2addb649188335d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cfc71cca697fdc40190f561a8f96124b8d59fb03f1f3c3f92a3dd8f17c1f4e4e437a09d9716b53ace174df2276c5e0ac6f2daf5b88da6e8b9858d7a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eda45093415ee9365ccf3b20880410869071ddbf0881d5efd76db24e1a0bd021a467323525a153fa65674f8e78e03984a4b320f1e5e24fb5b58260a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67efdd59ffe122374357acefe8699c81cd1e0912937bf4840749fc0829f7ca7984758e740665f517d176277e152c4c38c381c174fe665df468bf67cec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb0aaf60e33d4933e292aa47eab23e6f54c0a99acfd306c8942e5e444dc20b246176569e562db7b901c88c77feecd4adbaa9e0b3610b49377ec909275;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fe67edda90ac0ead64876d7fb606ecb1b590c0ff181391bfe11188c053ebb5144e0fc3cf8d171201e84fbf16de3ad19c2b4b9f37b9c4aacd5a9ccf1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2b3f031b5b379badccb73c4e69c9ba556d9d004a2ff4691d7a557884babaac1115f785ade9d9e9ebfc077fb4f202209bde644cb182e51e09279de7be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2f237ad99650372e471a293e8bf4f0128592672a05bea0ce9a5be0cc7be52a4816cd2b81523ab36cd0b141fb3842dd83211aa543dccb2d8258746a43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58b4a81bc75d7d774ee0bad73ad843da34c424485c6a99b3694b76a6b2066297435b17f14bf49a1cbb6598f6eb3d268104496d810ef35d336f5efc9a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h297f5de4dcddb15f950f4d6bf43520e0d18688b6583093cb3b22909fced629eb03544e441f4fa6d3f913d272438e47b500899b94f00a27d0f1dd2f1bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb811dff06a685ba0d760382b08b9c4664011718bfd01d84180c4b7490960f031c0fa693b619a014ab8d9a4b93c70dcfc3937fe8c4eae7f7d5ece5bd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5755bcd198673be3849fc615e49953110254ca92b4d8361e16f89cbcca72f62aaa830b0a08fc36f2336853a50e195d19fc635dbe489e761ff17e310f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea2b104fedf86afb864e0e2d425419c57ab510f7679028be89db54e64341dc0807fc6ee2bc5481151b3d31975e3bd64e1609121449770471d60c93480;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4604c345b545dde50d2c6968302cae7d8d2cf88d8a7c40d6d443138cc5967109a0d360165f2cabcd1836231bd38fdf1a2ff80aa0b22a320cf84f8a7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c5e860ec4382811964f157978f2d90c02011965242a531f986fef09d2c9bf8ce31c9ca20a2d1e93dcc8a0b26bb9a7680a709ff40294a1b7e1add4df3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3c9fdae75536b45f9864adec99825d63ba94a30e569b0ea945184acd1d0132a0ae10d6cc98f97e41ca5d552ea5f3adddb970e9cb3d93c8a8a5148db2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7a96da878aeb65b71da4c267b1b8353d7e9ddc5f3b2bb721cd8d0967078d9ee34db539106ed20fac820b856aafff5ffd6178d8153dfe7511e767055a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h798ded15efaa95e098bf3f5f1d174e1db36d3a6f0770e0cffb247e2f3f11dca7ffb268123f5eb5d06bc9564e4135f42c56b215ae92b434e51a0136ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h719d8523e2ad32af970713fd1b2c3863a37c64f624050a0b01a9ded3021b2c13059b1f7d15773bd27a96e1c8e0e88519ce3e281d59794cf228c506119;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd900be134efaf755e593aca94c94c66393fb740fe58010c4af91e6b5df4a0a722285891ab58640f4e4f739c321076d0defccb80cbb77fdc4dd4ca47b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a13611fa830ac95d1d514a8caf23b0f28912e07650bf0c90fd7e909fb4e8ffbd2819d85e334d0f268da82882b9aa65baa2134710febb412cee54e467;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f5637253b0746c9ec41acfa6e49ed2785a260c5d499997532440e61a8717695b50ac6c3c3161d118de5fb5b1364a626b7ed65f069f32577b4e65c96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e4ad3e33839f1ced0e876cfd9637ee15366119ceac3f12815288f286468120c338baee445e9872116bdc95305586f55828507d37647a077fe37fd169;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd056ffb24dcec9fd8606b2188896354806ff1c24212bf48800331460c10fb01fe2a8522037fad785a9f97019870b4db5bca5e5372bb2dac1296140dd6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3e77be7498e05b5891545378b36122d5b0fdddf8c5b9b3831bf6500f82cb746f57b271adb68b08f1d952251b8eebcf227f848e07f2311352fed43924;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1443e231fd590ac1b16226673cfd5241219f0ac83076526a530899fc2969d80e67cc21cdc83d9ee783ca7937a0483efe5402871b364ec69663dd89af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62cf6909d20323bd469194900f1ff6cce587d3d4bf9c408ffb39f2662fb8ea243773a1a81237c9323c3dd37b295e25790bf8818901f20fa0fbf21ad32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dee2ba7c3afcd23ac2f050aadd6a8d0264c3da8cf778b0e6f876db7bbe88e64efd593b57dd4debb2fb352dce0d4d9ddf572cd8ad1e0809f7d246a91f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eab577c995a9b7e5c51e921734a2085a8774236e8f6f812f50199146c1d04a6488d02ffcfb04e287d6128f369e2d3ccadd08f20a8bb7ae21b4be7c04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32ebb227ccc090b5404f4cd2af0d22f58518c3c652742d9cdf92fe449f521c73a380e569362a60b13b7a62b7544e02e745561051715f809a3aafc89cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0967f669b3cf8b845af12b03f90737fb86f2dfb828bfa4bb68c0e2918a1347c20f72d9d7780514b3dbb9b7cec9c505ef8ec0145f2165e22ad456087;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4affbcb03fb3e5aa79e73f30531473f09237229bc5d034b382150c61e49f9908b858707b40947cb7eb3eed6c0902a0c2f3e72938ae1c8bf806b1bc60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf42b2d7d0114c759420e64f520cffea3153074c46df86e7ff107c978e8b6f0f0190a9af99310a0581bbb274f09ad5313cbf8e0b3aaba44a2216a66e69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbd0787a58ee985c53c6beccea9433d0464f5c926d9ef2d57e042a2882649b899edb070b26c3b80ed464a669f5cffc2ce17bd2fbbe6698f667b39585d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h847c9e879c51554083907cae01d2572dea050be6adff6608fa4f0fe2e29b6f9a90bb2691d7f6e2d744f1f6ad77fad74d3fa6f81b71747b1c41372953f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haae1191f31de5de22688cd4c149d9b71fc78389838634383b3c6e1be04ff975a108f634a37122375ab9b9fba7fa9547e052d7d5f943aaa1271f359aed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23a157e343dcc642d9d90dabc4baa86ae31653253b6ae6cc37932d3aecb039e950a8457db1dfa0703b98bd23cc9729632aa142609f8be5b73aa5cda53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha207418d6bbb0c77c16f7a6bf8de8a1c73b1f505aa65412826650a6a386c9a4e4bd270b0ed94925b78a79046430446feb0d4855764cfd4364a8e90644;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h200b23f306963310d1519648613e08c8c76eec2f7ee1ba1eb560bf9d128b535fb76b7f5d456b15fc1517d37341226b804164d6a8652374526e93b8573;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27d40db15087519505705448ce6106c2becedb77c8d6d1db439351e4d8e1ca3d78ef4adeb4e88edb3249b2c722c603ebf5084de1ab09c146d0363ed5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27e83145ef693054c5ffc4ffe9bb595b419590e1d3d5390c27515a7f1cc5b6286f3d44fa40838f3f8686718844996361bf91914a50fc7e3b48033f396;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56b080348dd5557f0f594cf65badb24f6159261aeccf974daf8770877af2a1f649218bdb152ab75f722340e88f6f0f4af26a163a037d66399ddbabeca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38ba1c37c51e4b1a358f05d168fcb1386fc2260620eaade477199dba9c8ff1037e964b75484bd3c3c09ba8946560298e692206e43f714f0aa2e7ef343;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7319c8fce9b0e41677eecb083b92c7f94ae53d1315368f31f2347393020d1196569b821baf1e3e9a68b8e39c966b16cee00d15c4906e8f07fabcc00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcceaf13056d3b1b479b371e41a7fd08789d4adad28c4debce82de5c06cd636f7df06d9eee5bd45e719ad9ec1440162a41f6bfe543d10e39fb3123d07b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcde930ea4eb75c8e6db438a52bf645bddaddab6a58107ae3ae475aa31d5b9a0c3a4f572a86b3d12d7ac661fdea81dc53374712226a27f434bb7ae009;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h224051755bfded6858ea38076f77ff0125fc25aa4e5458a56de66c7671bf47595b54c49b440412a32403435103f746bd37a6c951d8e06e7e6cc541280;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b0183f07f330dede527c8919b8c4c038d39d3a90d43c0d94103b1787f2b7d948e26f9ad53429a5b1903cd7f2cfd13bb6c70775ad9067ee49defbb8e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef90c864150e623602a7f595c0fd7a6beeb3336c456f7c1fbac49bbbfcfec68294fb9b848711f9816ac7ae183caacc695c90626a1caa42422fd70c0d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58184e55d9e17f87e55f16fe8abf438194fe993e20416ea25d21717275d967643a2bbc6f41114e113aca250a08cc15799cc79ea5300c2e788c44eb46c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h898d9c3a3d3fd005513cb7556ca123dd8968b344e8bef385223bd363b3c436bc4077027837c9a3c4e38f8a9e64b86b0c40ed45ff0273cc926d3aa2817;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3aff38027dc5836d1eba598b2b79618f6fa103d7197b9253ca9a8728cc9e71416ec1ef12ddaeb2a007430d2d2aa81ee5f2c0ee1da5c3687098569c53d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h388672f16ddbd10abba0e1d8cde23c3d99f6dc41de68021e9e5171f950902ae4a41905d631ecaa3186f73f769c5b7ebe1f7345600bcad1f72fd67d70c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h593aea4222abe6778fa9b0e029ed7d4b73b56958a6981154ed4d5ec8c926f6fe8ec4eb0e706d47e598fa515f0304559cac8823a972f32e41fad8eef3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1cc02c27e58513c0226a505fac6e7fc256739cf05cf278f0b4b4c063e535e36cadd0677a4f9e78c88bf7fc39d19cb0738c79eec1be5ca25086398a82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd626ad1de6123636f1199c6ee5c25aa2e4d12467665cc346f4576e67c359a8f2301a1ebedb1bdaeaae9a95f9270b7cddb1154c9250dd827a0c67d1912;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b920a0765c0846a2628ec73595193f3c4fca681e502886e050367cd7461851d92d3d37338af907fc3163660cb5724e21b9dc654aa5a20cbe47a98697;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ce0d587a40dbc17bf92ac72d6ce5816b14ebd45278e675f0f049a97350f8eabc0bcfe9c25cde4b6313121fea4fcc40d1848acc535b7af7fc8d0cffe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h759113e4a1b391ed1b0b0f532cdd820a194319f90fb6d8ee66854712134191d17b4d53ef488b0e47766103077a0d62ea75286a86588adf5e8f220c352;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b92d6b12ca64f707a0c032717592ff412504344ae6f8b8f68c4137dd65693604734dd227355781f7d8d57ac8b5edf63f692a545ee82def0fed729b34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e8eabbcbff84387fd0ea888dd5f2e0da2f3063c1ff77fa98bcd674964e2cce42736f61e24e593d9463223f82ce467d55bdf4f87e1f1652321bf7e05b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb08da8eb6a541700c32e422be8caeccf2bae9185455c57e8cf25ad09931be03490add1bdc506f80dd5b1c961c88fe0f6a5c39308eaf1da6dad36c890b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60d6068f6985033a5af6220a90f5c99e35865c42ff9fd778666ec7981ba34f95234df988cee4a046da9d8e4e99c9dd77793e68429273dc23465642c8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h113639835ce2a9ac7dd28dd0bb94e192c012d28ca822169b5b4b6d4ff46218bc46d109246602b8d095c175e0909a9daa8feac7e967bd29ffa569bfeb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c85bddba0efb14cc1bb2e10b821ef51b84106511a485ded451c0c01ce8ba6262acdf1a51b8707c5222f4fd60211087a11e3f6da9185ba5ada243c183;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9665c5c798ac7688b0fa7220fd785767dfadbcff11a1122439491f999ea81d737135bcb2d7bb8c829a1d4961d8430eb912a1963bcaf734ef2e19fced8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d0354c1e94eb19c10b7dedfb6c56329362841e0df6502d2b113e785a4ed1d8057104a65679e4b28fe37b045d5ccf3abd077c85b331e971626fcb55aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h666cdd11b2df886bb2ae600ad00abef24b34586b8f506dbd6dbbde217a54a2f48be05fb68916d13c416d7a842450f99439458a1a4ac3b18db773db8b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h285a3263a3e81124936f829d962ba57a97b174ee84a532b8eada45a16095fa34f85af11372e1f9dfbb195bc2dab68d7f446874f81b6a0bf6cca186d92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16b061ce677602005972977a1ab4dd24012651fa3670b779fbcbc50f1d12d1d35c1c89d4042133968dddfb0df99bce48aac393c38591d1fbb58d56f95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65e79561f386a847db62133fc81a8366f1e698ab1ad4488c1df886ee0a6a960f59234a26a0170323255d095bd3f6f96b550d3de13c94de1167feedaa8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he68a237f9921e7f79a51a0f53b4b4617f492f67f17b5bd82030571d00c66aeb5afb9242948d693fd9ac99c3fc63ce4d2ba56e9a26cb76596492737645;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc0c95bcb6dc3f068c92cb61a3d31ed7121f78e346b6f6c769064bac1828bb8cea26c8a6c4fd109bbe2a0becda86455b2a9bb1b2ecce4b38069b4b9ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb024736d14ef6356bc70b74e2a68c2c1d19a3d9c3e2b42d74fe2de8d1a51d76f0ad9c23e88ad26e7dc796dbea1b2bc835f4d4b3127592486cadca2686;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12d476164de89bd0ca63679e8ea04017ba10919189884f43c926f4bd57eb3cf34ad039b8ad54bf0be762c641924e15afd0d107aaa155739c234156a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h766d69c5868511c7999e35f77a9a5aa52e093e524b243119223c197df4968f6ecdb285c03b51a0e48ec40c42e1736f432053f89115855c8eb39762f11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h161dc988000360a5c9b8ade767d29e4a25e23d0744ad9018f0b166cd8a4a02a3338972cfc8b9a936eb61ab331bc3f6df8caaa89f0b7ef84e634444ee4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fa884c79f8ed31506779b710533bfd141356e9aa2b9f43b8f5209978c3616f4167bf54bf86eb828f363f620d92da8aeab8af354f2cd5191ad800ebea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7310159e9d79959ddbf277c1d25b8a5cc850a93bd9129e53ddca5decafc02a41c5ee34828136263ef1ed1fc12ba8e44e53f591449262c8376c790997e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd37de6b4f7ba3d86f20acd749c6dc5329f0952d2b706b46a32e5ae4873e9df1584eeb1510226e3532ad4f294e554d2ba1a585eb4b492c505864a79c3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c75f5a4a84f535cc856baf5e8273ec28d750d23190b35ba3a300982c42d18a9ba3ad32f92b99852d603b5171ad2749204e811bbf1745b97a514c5d3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5eff8b4d42fea3f449ef7a474924bc52581c5604328776f663b94b1d7a1e672fbadc76912e65636de5b198efe09226c49e12c86ed4f5dc21263479ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd21e9a8187859845a01b0b5a877b51320afe9ba44aa8b1ca4afdab7d7a236bfa0c79b5516777375bda556f38f1d9bf2935898271aa9a9b849bd0609dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e25d0bbcee3665fbd12884bbce96741f1e37aef1bdb2c0cb1d3e4cc4ff66d2d594591010fc0405598d33ca802dca82354069d1d54b6fb4a5f68f943c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5720f5bce4d7a8c0bc561f4ccf1465512e907f9c310536dc35213d3d332caa78016307f025eff5eafd593854b6bdad2575f8164dab0e73a8afeba5cb1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79d5c514b3c0a0bfa83cea43ee0cde1dcd46a827610864e8a8d821bcbb00e52142a7d45849e397acf97b0f9450841c28fb00c5213f3cd258efd13e12b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d7e70489bcb2d13f3f22556571399570ffefab5a7df89146a6ee0bd55e602a85025c551bbb6e0b3ef039c3b852e56006bcc74ecabad51a5d3c373b91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ac237acecff5ac6bc94bb3aaa7847859bc89c6a0e003d708104f479aee4784c398f20d09cadecf76bb089934e25df66951feac62621b536af95cd68e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26e09cc8cfd480389f99be992721af3a7b0bb3dd289512e580b3deeb4d5a34e73846a6dcc1f57efa8dbe04949f78e2e36a386d2b24f138861b382eadb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2c8a11d17dac83de46eb57a737be0117453c034851885a78c5b23efca93a7aca06d9599e9632bef060096b822ff8270c8ee1b1baf4fc84c7b1d62edb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h707df73331467517af0b30584769439f10c514fc6e0dc41ad7d97888efc2d62eeeffa7b764b41969b733984fca8b889dcfff5a0b4c05f27c2f6331a66;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha02cc96a0a01ceebf5a666c1691bd3985d441cfd676d039864d1d83759bb91b62608520e91c48c629939fb11366be87751a4ce1718e99803a2d9ae5f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5f1ce419439518381b0dfeb35ffd21fcf51cdc815bcb4c220c440a3742fb7d7392af571f7040fa2e94aa64f2fb55052fb96f725c448e3f95f30cd7fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf04f39c8dadbd5672a1a717ddf5dbbc3963422cda0e1fa56f2aff48058f8a7271279c7d275023ec017df1423a79c985d5906643bd2d01b5fce4e3a495;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd95734f005af1349aa4a2abbc5ccd95cc30a12428fe560fe1dacb04940140e2d51b3b22a77b424047ba82c0a37a87ddaeeb3953a001618ab2b5ebb9ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57678e0127d08231aa88544d90a3c5198d2b710860d58d4f8da2273b564a40b4f56d6111ac49758b29dc53556e0b68646a116956ccc4b23d5418787ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29ca977321bfc2182cb3a67b0c8e279bf007686db659e499b2c3d28cfa00ceceb9cacb60e40c75841135f1f3ca103f28631f800bcf12fbf244095d77c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e9465454f8d1775844ac3736386a2974900ca3d86a8b29a617556db1c6c20deed2888439580918177d90e9fa4a08377e296bdb345dc10c9044cccd99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93da6dc0ba60102d6331f48ac3a4cae51f489787ebd9792a2b8a8773f79ed85bc1d4fab0232e3c0c99794cdcde6d90055649c0f521bae1ca0ccd8eb6b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78fa0787922cf0b97d38d170ceeb3cf0d45ca9cde33fa52a7d1b992c22570311ecccbf83619ad31b9d302d6bf991f17123186764d8897f4a370d8f2c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3576f93e5bf8c7d2a1141703c054a6aef7e4025168a337ba493448e3d2e9bb09ebfc83cab56ec74c0e45e44240fc9e367bc6b79d756a4237deb1a15f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc70f2c58d9787bb73542ddc8eb1406e7efd05f8b92a5aea812a234583c3bfd86b6a657a0758cb8acb518946319065f0e10e43da2dd71d12183380f03d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc47161b53447a2ce398bde9b7eaa3afb73d540a30248d8a95ec6cc8e839e6c5ff6713ef05a7b13d3ef661b77cadaec3c5ab10dac93c5ad46f27297faa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h300280221d890f336eeb7cc0f2fad5eca1dabb8a5e8ca1cf89f8753bef53c1b30bba277976c475f52a8b3f20860f74833e56804f953b8262dc9798bfc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h130e5d952cbf573f48f7d2e519557f9566f4db7fe36f0aaacc77e4ab5bee273f974c09d5aed745a012707edb80bc48cacaa10779fcfdffbd776854457;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54402a65e49304baf4441e035974d8068fa77d2f4719c70f96adc91b85e698c779b1595b710c79115bd70f60954c7ed15ca0eded66200e9990c80a78f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbd2f137ee97aa9cf5966876049af88e5b2d4a797807eb06799274e7699318f3adc60e58c32f27eb47ef693d1e3e4c97bb3cd37519bb85836b30e641c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd663c1b060447f22a25e3c6a67894d76335d357a23771bd89629ed77498e0abb43d05ae7783d36a858aca0cfad683d480f0a08ea6280a2d9a0df850;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf52aaed02d0f5e4481ad9ab1419ccad523a7ec0b810463ef0406cad876be7775a7822358bfdb10cc4b73de44d0ef746aaf9a65c505e7b01c6a4869f17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94518cbfe316cbc063940051c9b8b3f3dddf7e3be1ebaecab3a2ecc8d4b41410d6148dcf9207365a07f0344cdf5adfe559d27d5a2e1a577ec1e8a36f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h477153bf335b9ba7feb03d9bf8182cd8ced8f279028939f0735bf193a7b53c4e10947de62e82ace118a41abbcc8b75044cf5519031b75c3a4367066bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39d2480c92b4e607f08181ba51aa4c9ddca420f6360eff7507e02c082958b6b1f1c411078cc606f715112c360a9ec3ea8607a946d482b4aa117566938;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffbee1fb1aeff4d5668b87883fca07e06c39aad58d8fabb6ba09b204458d283037331ab64fb0d02f39872bf09941f1d00039bb99425f55961b8c22916;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h138f9bdc38759c346b9b952625ab7a17e05a59b6e73465866f16c98ce98d32ef274ae3fd32b81477cae1bc59cb07d81dbc79c0b34b7b27515900f134f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2dbb81cc39c83f9c2fbede0ddda6f6ad83bfdc6ab14ef0ca3809191ba18a78ea38f06027717246b968226234fece70e5de4f31e2c4ba1270d5ca43ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf282e0f1c77491809062e3030f3c11ed0828092119738ed513a021908c2dbfc39410f82bb4a3d6273188cc17e1de225ed45ede9dfd43eea92438bee4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7505d723a0ca6192b458251af41d666a2ad38cca21f3799500a3a51e2f94434d64fcd8734aa6d368283ba82cfe318c6257daffb5e011f0b8ce214df59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h132ced0e6f3916516eb54b8f3f743018aba2aa2641b7bc12f19710630519a85436c1b8365ba89030a3b3d255481549b424f891e00b6ce6ffb8cf4b495;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5ab4c6b275407ea616c098f1be1af883638bc895b7440ff2ae171c5ddce43bbf43acc73bef0f71a6e3fca0f340e1f62301b4927df20aa95f13357dcb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70d33811ff5a52d5ddf1f38ffdfaaeaefca50dba1b6c4d504ee5f2528a538fd4340a7890e0feadf67b330380758400713e831a7987d2bd548cb4b1306;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58dddfc2373d69220a30bf548a6f3d1b4fafa693990d641cff5d22f6cc1159a83bfa28842f3e10f702cb8af0c46a18be389166f1b3339289e73c7995c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6db703046a24027fcc20c06710d1f0900601183a331d4ba791513775785bf4f64d4c26006db8fbaa2810a821718ef2d9c48734713c7e2a828f0963620;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fcc24798dfdad7ecd7e280dedc90be7597a0fa1e7d6af34a6be3dda82d9290e0473580a79fdbd4ae92be855facaaa8757727819ba66e213a59e0901c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h975f2242e41de85f228e49bbdbd45aab742f2299f9890b21b8899ed079ddf8aeeecab8cd80acb519e99f0407748051230366cc2bf6169017392862001;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92fb475b6d79977e476b6ff4ab44d28c52e321c8217a6f82634c48595e799c4df2a8527939e2b3866d83a13346a8d78902cd2d66e138892fa90cc91d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb57c015de746c58c16e06d29c47dd2f6a0a2fef80a9ded5e3475f364cc16851e64ecd666e63de17b2ccbaf8a69af18964ac959c2397653c2c17697990;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc3811f5727ce8680968b46d48fba3ae50ffc856d3781c34c130e8db234b441ffd7eee04d331fd9803e9db2ea494a9c16af3ec7bfcf5640a427994561;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf39b831729ac4604414f22318cf17e0da3b791a0f5b48083ef4cc48196af8e25ced9c53ab408ac26e19dc31058d9c098eb69dde9110f6a160393c84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he512e9559371a8c2b467368a2c0710c418e61bb7ab72d1e4c38fe86dbd794c9001e95ea5cd26af399ec70f7c27344a3ba3d2990257b5026d08e6b2ed8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha30d0b1b903e1353e9e705ab388b546abbe4349e6bc38602340e6de748a5952800b29d3854a22f42f685fe597cd739d984ebe6d54fbd76283d3be8da3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h323af99e5428833c00d5a8d11823e3887c62911c713cc9b939c5265e099e1b215e2db429403e88dab13048a4a4c545f62c5bd48e95c88c07fd3c9b9a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h815e07ab05b5ba501a15b7dc6059ee7edbc3c5b2c48f8f296928c9af7202197718ab84da003f1bc95f50865b4cbda49dc6f95cdea1ac39b28a7b20d56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6606150bacf34c6aa5ba638ba99bdf29f1d0716f87bc1a298d93e45b61605ebd4b80b6fcb1da7c3201f5b60efb43d3f654d669faebba52ca9dd938dd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e81133d641dd68ffd4d25beb66a55e8c7ba06d6c8a1bf7dc0939782ae59f024008f0f5ace533a16babd1c9d7373f900a3ed142bd239415cd9e9b8bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6792a1e5ae759322c2d679caadf2e413e2faf0c85509825ea01dec209d8c18647eaa92ae0a8cefd719c396ca50c02e372f2b8709e98d794e43964101;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he94870352f996fbc5be7d225a9afa223fd217f74ce8ed36de08b1b2093054f9e78b2153e7f68704e602835f2a36cca87697ea0fc236528cdc499ab4a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ca0c00618194fb22ad63adc883edce18821ee8d1faf492066f277e22af9a1e6f3c065fa8499606a076fc35933de1e21a898c13c91e6f24fb171377cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c6ffa4b4d2f06752e3d386ea1c694bfe2c7d2085f164020dfbad0dcd9dd23702d2cfd85c19be6232b9be45975d1582dcea4cc8c9c23c916543b35b8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1131edaaa2dc58b2e6af0536b1376e938a877ae6998960a39bb2e7129eca5244337a1a5639335da3eb1e65a8b862663a898a0bfb3e184126edc2cc91e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h424a8337d62b2271c8e0ca51b6357dc8f879b8543b9c7addc3e48b2567d862b3cf4f9df9e5f0fb3416210e7a2c5a9347ce818a17d25adb6da23d720a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b48fbbf2abea26c726068394ba25d86145b4f839ef1a99f19af127fdb91d9c7bffab81415e9c81f22ed6d3fa111fdd99bf4d0b462394213002e5b8f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb59252a4117a03362c54ded310c784cd0e972b7fb09391e603c24133a3f7fbb1a145ba575a8560a5a9e65c8e7736b6842b2a030b522a79036266d7097;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2f52beb7477d4feca25ffda6e60eba6d014e48e8c4b9a2df43b4689a43e3d2c79610899fd9fe98e2d387a022dfc7977f3956a868a18367370e28e7eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a54138c88329c7822cd88e3e8884dd8ef7772becb3038669aa28cd33d104934850590c4f080f66bdb3d81bf3cfcc9156d4e44c895513327b5c206e62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29d99303ce231b31193e22d1d7a787415f3ff14354bba4b8c791d0cf4a4efe95e09dac82401910c03a3130c4e0f3d2c313da6309ee7831df4e37fbc2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f9e024c205cfcb6a357013706e134b3209c51eb5085f911421e69683c38feadbf4065710fa2e4baa25dd8379f8263df451bb6b4b4219330040c8593d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd6212c4dd88b2701e8dd7ffcacb970b03caece256a3f7208b03444a41facf69446ea735e8ee375210d6f4b21aa01113d9e0bfb80f2c8a886e6b6d19e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c3a1867e718fd1cf66754c5bbfd7e106d9bf009f1ae446c7b88bf222db3f812ef9813924fdd1e77150bb083c4b59141a6e584ab4929e31eb0ca0ebef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h692f2b4f294ab0e10268c4065a8086a649bc439a21bb9f712b4669f028fe9953a3806c39ec359525dcf719808a38326869a9b9c0f5781453f7644b7ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc468d85e1da9b5f60fc3c144e9e180f7852818f6fbd45f53d5c9b6afea2d05f6f5d816299fa866a518b1d01dbda01a8fb9520b0211038d4551b664ec6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92843515702dc572b8d63b14b1e5d7851ce01aa5656169bb26ab0e10cff76e9a3357ce8b54013de34a9aca80890a242f5f7641a76a8d345aea4cafbd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20317623dd27d9d5ee076b77eadb4c05bfa687c28337173866eacf940c072c7050cfbea361658adde7b262db4c8b2358318c9a8e68ee9f4f9ab1ec837;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88174e39606ff53c5ee66bd628808e713d5a522450c4978e47dcc8c2695e525e8a05b0191bbe815137a13d7f340dc5b808853a09e33f6198e12ca0572;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5727626b676ce4bcab0944fc97c1a07721aef232bbbc7d1509288fb7145c1ea440b5c1b24047488d71928c62616ce5dbb791695eb5c5d1ebfe91f2b7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9407f1209812b7426abb9ab6fd792f172dcc9764d988aae7369368f816338eb829d215f41077b6bd8ec3c707af42029c7b80c9a89de265dc8551b8bc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf74f83a60e4a0072a93218233a53ead78ac1d0c727a7d1d710454c68b38538b79abf86642a1860a829abfe983f31faa29257200b7df874e779f44ff81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2b16ef8fb642324af0c1e929f31afc8664cf83a6d508449c1cf06af4590747bed782251ce52f163277015344d239be20a04dfcac44660e73e34a8560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he87fa45709fbb9d17b73b7c5d009a872f352b30d413e1cd6dc0c2e53655e9acfcc48720212c73fe2d9a2cdd5e5fdd3ccd586b8ae4bcb9a710710f22b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf736daa6be1323652c176791bd612866fad81eba0880b47eea114a55eb9c17100fcd3fa49828911768b78109c7b02206e3e138742b4f72ae8bf21e032;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9081221750acf350b955ea77319eb0664ca21a7ac634a0e5f03a43fbdcfd96289a34adc93bcef4cc25941610704a0484fdfe26f3ec04f973c4fa125c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41d9f1cab1342403704b825558d2f3ed9015561b377fb9ce4b969d3383a7ddd634aa258cd8ea0b41d4ad469cd7979deef54f7698dbaeefcb60dd1bcad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9707c1d64edd5a07b4f962f943e887f1c90c0efdf76d87feb6d996313f1555f3428cb8151047ca7836d1956d224811aef05ea6bd758ac389eb6cdf8a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2dc5cf5403e06e2511f015517a5437f7870959d8dc2e21ebbc34f419816cc2eeb66f6bf8e3cb5bad5ca73f66475aaad5a6a77c885c3bff8b3cf44181;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22c7273c2d57b964d7613089760e060ae06b30f5e0de902db9e5b658bc4de39030a8c5c1453b8b498f35d612616b50b59b578887cfdb8e63f8f8581e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc856621aefae23db8eb5392d6f695fb0416bf080490c9738a66a35db3ede6108fc717c394b7f17aad800aa6472a99d9646435ee93cb956b7d055413c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b2b660918d29b12d52cbf8c395ccfe03a57ff98cb92eaad4f15620d4a70ff8ee856ec828a7c90f309dc338b71f8519c531bb89993e6bdeb8bcb50546;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e4cabc894154a5e8024719387cc34005c94f205daebf6e321f07ee073cc1c2dc3c54e1c9646e260391c83e4db02af0f6c73c0e7b3503af8ffdc882ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51aa5418e343027dfa6097459b9e93297410029fa95f55b8292782416f887ed6e9674d467b00f4f8239a841937e081774807ec0d688a9c8ec82e3d760;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdb3dbea0e4dd87fcca73e6415b33b61c9933c035ce3008452e303d412736f72c62a7016a99ec2b62f17d51a13b37d698bbb2b47c1ab1b2af778bbd50;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb4555b003356ccc57720e51193fee18c47b55c2d24ae8bc3411d13f0ba5ee9ed3e60e46a385061a30fa363b8f01825f0d8b72316fdb8f4c9f5fd671a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc15aff4f091429274efb91c662012db2e222afa4c6e737d3841f71e2a50bdbe0f226890503db9673b38281a27b49419ba304d660cfd852e043d736cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe6f352fba1e5d22a0d41b5682365ce806b9daee061163932c90e1997355be556314308d9d4d4aadbfdab63cc8c6bf622bbc50aab2578596eb85fc7e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a0a297caa5df3513f008a31e7b8b3fefb0ff2a2fd9129bec25b4529473fa3105759fb44c42b27ce8f5dd1c4c8cd31acea29cc52d8f862904954c96ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46ad79358c422c240491f827891c9f1dc8689aa495909439074c0a2e01b811322857962f14bc530871e9605ca72fbbad93853aa2059b1cedcf67b832d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbeb850a4c5d72eafbd4137c6de1c1cd02fa4caf23ed49c9b8aac6334054f55c38c87192fdaa08fca75f02a073efb2f58ef83e2402884f86fb6776f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ecd9ce0ec0bc73881c58f7a293686bd5865b9681d4e68fc9f8488aa6c99382249ffc83e5ff572cb67d1af1cc78767e55d80a6dda87e8bfdb3ef3e564;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5565a5b28fa0d18249ab3c2e950d1428545fd83b8466b961478aacf8880cf03dd22e8ce26af702d655309a57d029eceaa3c921b146b799a1fc4f089e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h245bb6aa933404fc9ae67ea825c8b7c7363d3e626c15b68a5b28dc909449c40ccde602ccdb0eb902f2a4d0dcb8258390e80c6e9c46858d7b336ff1bd5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdf3c1a37b0a19e6e119760edecfecc17628ccc520f34558d35f07d65dd561222285ef086d03ef4a55314f8001e65919b16a7f38c8ccf35e5077887ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h339af4570e99ea5eaf75f38477dc745186474dea461d4875b50ff4f7eebf551a0ffe7030602ba3bf37e835a28e8af5bee2f5c1ffb6e45183525696bea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26793a6536290c318084b15068a2cea2c02262ef52f6a62a356af6a5b95e470f0e9bd1e030f811472e2065d89977410e7b0a425b8c78646f2566f40c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23501075151ff7392338377827c5cb62cfa9de6d05ea21a28f0df87bbaafcf9676ecd588a7a186ea41bc1549d3546e3a0b96dc7852ddf612d9828a1b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf976b3ed7a679e6f13d9b400a44fd6c820be6d922beb78119eeab4a1b3eca2ee3ba2a5143eeed604fe8735279380ebd06e15fc5de5e5b1c7aaeba8daa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h402cda4335770f376815db49564bfe28ddcbc5bb798f97b172062e3f0e98a8a03ad7dac0661ccdb8ff64c655e5e0e7a2418248c69b3067911cfc788cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12ea1f6578816ed0446cc04dabfba4a979a04e09581adfa64a7b51f9509fbd31b5c043128c3a4272da3749c2986ebd08c65ff97f8786615ce5cb7a8fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99d1e053b92855a7045277ab5d27aa13e47de19571770f1818a9d064f2e7c92dcc26009ce20ecd9c3c8567a8be1c63ab01ea77fc843bfaf0ead35b1f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61ba6c22533ca99aeb90218aeb1a7e93d0bca40a524e4cb8bd4a5844503269182874e27cd415ded1bb6b46adf9c780034c58f26a329ee06c2cf6115d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1d7db67a4ee0e0e6299154097eec95c24c4834f025beb12a7ab1c61c7181a67f4f124b7f6d161d0dd37e867f062651afa62bc0fa4a924a6e7c551f5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a9365c9400ef3d1b79fe59e1356dd3534a719abfde613f61d76536c300fe78e18c97fb0eed8ba0fbb016e6d77330dc0d6d3c99eaae44bde32fea8983;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha82b26c7ab77648f21aea0ded601fda3f358e19a03e4cf926e052c59ed3fd4ecb16c1f9b4b0f8c242b9ee452a9b0d5de623c2845a8b0eab0d45946a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9df9fd6ee88904f7d0c6de98eb1d4d47fd6a6fb9e471761cf4baa501b7768ad4bc502f590b0368f4a18f09f6261e116ed8fb18463e3396cadb89c6ef7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcad19710c9ea106d588e0e1e839edfcfe812fb26c5e0b2043d6d4ced3df5efebca3dc2d4232ebe406d55639add51c8a87adfefb948c75c7a63b0902de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb08560f78d6aeb8527af4a5d5e4ac724c61c666308260d619d6684059e595173c6cdd1ae156b25846ab91dc9bea1f4ead1411681e1515a2dde32af4f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb369fbcd91e3a7d8d260a5e7c32b32c243769cee54ec6bae195613beae316ce4cc6bbc947332ba048f6e7f90c97a8d3122dd07f3e1480822ca734c698;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5387ada40ab825a78433baf6bcfebd8e27185f22e10679ec521a8f1a01c83616eda94002b9ccf513c54cc815007f5fae096b9a510b2556426321a801;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51fed610f261162f1d25fa8d91cb4769f3f140588fbb0b9f1769e786ef86f01df07a7cb08b3aad74f41c45ee1d972fb2da283585f1a8c797b176b55d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5421a2255dfaf6040f64c9e948d6cc15cd16f902c4cdababedcc89a428500a976080341b5eb22497cbfd042f1478f14a36a698fb1c93f311bceea5d24;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34d3b86e063976938fb399c7cd9c5c1a11f15e80d53d62db8d8ea1931bd6c89c8f41681f9ca4eee954a4b785c4d857a5d7aed2cd8a0f44aa2c194706c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h178d4985a846af36c03a9a1d7ace9b24678b8c14b97dd5c6758f36fadfa28d7fed20476e91e2dee80d7a0168ae297a612c2d83f9a58849e31a27823f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h208adae1207060d5ca620f7d9310f1a76c47be270f1a4e32d0778900c891299d706b34c3926df0e6ac53c9c41984e5a627150569e22ad28e4a18b41d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he815671fede86eb799e63270af2a001c2530e601d21a16b1ccb586809fbca638a309864c322e7d1a5072100aa883c89f0b8fb2f62053f0e5820e7cae3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h454fd78663857fc3cb9b1f2e419918a7c88e502218bca767e37fae20a287c3444a9fb348ec6e3a1be4ed981a70263ae39b3790ebf1ad2fe7d855c2e82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h224ca7b80d4727668c0b633bbf964ceba7be0faed59217e372b1c20260e9db94c7623e8167efe935a1c8760db0510a88a8f1407b7fc1551a30cc3a436;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13d2a5442497193e66d7cd9a42c516b025b889580228e88cac2a0cdbf40af0a9a4ed02716a0588ca8a37cf7b895d0e3c525a75bd109dd3a63c976d714;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27f4cd6bf960dee8384637dcaac85a820b191539d3f1e3ff3f623c03a3fae49d23110d4929a9fd5e7bd463867371d4a4794c8cb55bc8bfa86a7f9b58a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e2510ad9c2d277ef7ca9aa72db53443719a4a6cacb6d78bda3afcbb54aae5826338936dc6ab2167afc110cd2933d7d55fbc6c21d843f90641be51c0a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2285e071744a6b965cc66294ec0ac6b222c457d07206260aad6495ea741c4026421bba448dd6e525d7e68e61ff268f7237fb5cb961ef939514ceac34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb256abc56bf58fe64613152d39945c6e08396c64cbd42e721232b0e1cc8f2c8e7c5f6e6ffcb8443b0f9269ae9caa093d9eef21b419802db3a0f2ba1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8247c8afcda7a4c915b090ab705168b1de16b10c8f09b7597bccb2b1514c76acdac17072c75aea3f59f07768226ba68910caef7c0e7ffd5bc9fe5cdb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86a54f511a2932536c9a33831a219dc58dea19d3ba6ac1f1ba3b59f5fcff832987aefd780c7d618ed6aee35e26d896cc0f6f06ee627874a05083c3318;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b2e772bb2afd157f88fd686da894826befa57a10090f8156bda0a949637531cdee7efb2331fe2fcdb5d282849044948de2640a1bd8dbb74824d440c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cb52c14ccd3c29a38440597777455368678c384739a7ee70b48553f4bc87a981f00905f8e561eb3ee2924660a4d9991e2dc7e2ad5cc0b77a13990405;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7715ef7a87a796676ce875263755466105eaddd339081cd0817d9fb3cec11e32c2090bb35f1f38eeab7f5ba03f16388b1313b8b940a8e9b7dde50a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c788a6d33b99080ede589da76acd28557791c7192db3d7cf4bc1eeeb4ba3de114b3bf746fcc77c16b4e27adfa5bdd246df68d05190c1771207eeb13f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4d14b4abb23148874f1ab8b852fdb932887da50eec7d13eeab8f2de9ec9a2099d85cad2cd513adafa29b0ed0f2299eda6d745c8ab1961c8dd836a7fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he12f6c50a9488d682f8bde47a7e2ae09062f502ec5a517a9f5b6f5f8b3a4090810f1ef4cd24c8b53022cc2fc0048b38e263f039b82adceca0c3fd509;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h281c8ea0f71a3dcf25dfaa503ef6bda96c4cca1e44befab619aa0396b9be6afc5c63c2756c65d1290ff41c529ed1d1d546008aeabc4727f69d20bd8d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bf45c262519769d8bd8718be45a9fe7091a6163769c69d25039443a69c8ebd42ec44451145972c9d5d1adf0a14bbbf34f376298fcb960670296b9e0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32780b56820b565c2b840fb57cd192e835f08e6036870fcfa8a1c8b6111f496b743654e7f1a503c52d4d8a8688cb51500c4d560c23263d75e95e057e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1c23c6eb7461e715e6e3f71e010a5570ddd8fb24e879c08cef8aef723996e2b56bbd67f9a2409e7cffabf50eb08794905cabd81294b5f6af7176dece;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbdb08ec2308573627a3e064bfee0f5301c5d6407218026eab2ec7bf3a57bda876a92e5c559d88a4f60a2012d8898371122abd72d0982e27de27805aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2de2c7f27adb2e33e03c4f45eac588bbd6152acc11d5e4116ae408af7d18eb003db8e992087ac1d86b213ab1166c68f330bee851e7a68d4ce34ffbc98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9330bbc737ce0b9e58c1cea5af8a63de68401abe2f170aff96beccfcfad7f81d061c78db4267dbeec1335f1d0bcf09feccdcda4183256534b5b7a18c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78a3ae94c505ec16224682d4d077b8698407c039a7c14cd5de38c2e5d98a34ab20d18f62aa51c076f0e7600eb78de3bc8036edfb323fcff042cd0f635;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb12bc07d90954ac5108352b749594511623d5949a15105bcf710779d2a71dac87c22f2d122a747f0b8e37ac71e7eb9b4b130c8779572187c19f0984f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe71c3f4d1db14f80615c19d86fdc0327898b5eae1143b539fa4a156630a1adccf928f134fb390fd30cec90bba2f534515770f5b51826540b4baf447;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6aeb590a148677f0f446cca9dfc68d62a22d91f17e4e43d7caa709bca1f516945aa6dbe5c45ab48ef177de632fbbb3d1c751aade2e28a4c1f20d820ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1c25385a2e706cc4c09c355069b5de1ae636aa862abe1ca73c166f15294a552aa8bd607b2a9ebb34594c7e8c5f19806474e34c59b937ed563f07632a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14fc3187023d1f0051622f06fa272f97983f2817c9c8b97aa3bc02e1d0474c4d4086a772c782756eb41b433155fa7178c2a6618b4ab70462d90994f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc4e46249b3bf658653cf651fc5ab5532c1a980436f468ad4d68060c2c72ca6c65dd22bde2dc3c10f2e3b04dc650ca1f834d9f4dbf69fdd6fef47fe38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4e72848ffc6bd2c7dbf66d9a9d7c4085654bc40be8be6e14d2307476075172f68f678ed6b301d2b83d4a17b906515bd3b50d8ec62826255d6b4b09e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef5996f0659e173deb665e2db239f23faa8114c1a87056beac5dc0865f7eb00588f8ea4d0eaebcb677b1beac2c2fedec5bed64d789272b05d0bcb6f79;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8381e8bcf847985dcf1c0ba5eb93b9fedd17d5b45f905fa9820491d3e144787d88a48c5e640e14487a71ac53936e3168f1be3f8a704ce5c739ac07ffe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15ec4a0d6fc9fb17c2355f883649019cc173c863529e7cfb8e3a118b7093911c8610812ca141d4992d10fea59fc713c5f49b0d2d30792845ea757654c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3410d27812d3fda0abb7b44788f3c60a30fc6a48a528e60810a034fb3c442d7df3e591fe14af5dd1b19cf0e9927cf5431fd50fff6fe01b9ce296beff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca37bce969ac53f1bf603ddd74f9653361a35d561a242a16ec808ad8a1a2bbb099960a336ddbea92b63f38e26268f6028d02ef6a65e023b53ffe377b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h149fe1e7a903c6aa3faa5e7b0d7a2cf83d8a9c38ea65dc62d218f6be2b68ba5221c4520701c7f8c73782999af0a5bd7f05df776dc3972500f431edb2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he27e149d9b06b34df2e583cb5c37ebd848cecf50d0f8e94829ed2714de35dc9ccb4d13e8a0c91a0e5ce33c5c8aacbc29112c9fb770a0524e11afea0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48dbbe763d34c5d6666a312e7f44e73fab33f59a8f1b44e3a5aa0a03e4af8b7fc45851e857b2408b6a297cb9509a29c03be87c91dac85b46da4f75f00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8019cf29f30fb6c36d0d9e0960701c6ca60e842c162ba2786251de8cf0e266d1d940a0cf7a3d7bb2d03717d91809064b310b58eed8c21977d908843f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7c80c22fa385389292056eea30ef08ce0989798eb011890ad837a8c5f52ed0c901e7f8df958aba73c7d171125aae225dc3add40c4c6642138a509f73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h201e3e0002811bad3c3ff3614bbb2acedb2a3906e670644d935c6a11f57d5470bd03ce01a458785855c25f0d9755540df5f7f68b1a4801f9d5e2a3c6e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h801830423deb99e1e865e822a1c82fc68afa76525a8881e1362b3c33ce231e04bec6be3f3c0dec0a26814647e736fc26b641caf201122bc7c84077e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb27bd03789a3ddb32d3bf70e7e7ebd5508f0ed76d35a306235e2015d9c272685e4dda4ca1a300d89feb30f1aa640a17c38d976e725b895991aaa898fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2054250ae40eac3492b98e22230872bfe6a76277e88357a97536d7544f308fb3a89b8c96e77073317b21837bd621803ae88729aba605f4d0f2437aba5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22e4319625a288c5ad5551d799a46b212144b2e5dd177ac66fe62868999a1d2616cff6a1effbb33a6508acc682e5935a44bd6d7bec94403efc57f510d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb926e7860bdd332cf8e9ab330876a6a2ed84ad3030e1dc38ff97197ac85dc436dbf1f6f908cbb46d17c828d6e47400f550e4f1358c21a077004cb1a27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3325dfe01e500a6e2c606afd8efa276f7d9899edd761ce6090eaeea7100ac3a3d1f22e2445cf48a4ccf23cfdaf2c67da09acbf0d1fdc06b7ba4020aec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c586513fbc4a080b8e710881adfb6cbdde10796472258598b4246bf7ee4c6e72258c9fb940f5ff5aee9f89690675a03d46ba1897afe7347a6de54397;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90a890022bfed32f3a1f3bc25ecc0ea7a5288f853e2ba26e86c0331f32432c9f0cf97ba484a09ce0c47f333d92b30d643579f65f419b599b9747d254b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfad08a58c9341d0413a5d2b0881d1b4eaf47c1cc44b06d00f90f89721c5ff8067de89defee189439d37b00123a7ca1af8964fb4d0b57e3cb95f79b2d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5937257968654b768ec414198c02d29f46f45c9d680718c5000509034b063610974cbc742fc1f9c21718c8e6132089beb690c9b58aa8f397bd56725f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35d59ed24118889e88eafcd3f2a4af2974743d32f8f280fcce47891774750eefeee0ac1adcc7b18801758d4c9aeea5a8c2677af6828028a7153099c46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c27270fed0a65a7e3f339f30d4b40cbbc23a1aa9594b0a8e5724e116e37f7ce802ad9f582136f030dfd7d888008a34d6af3f7e2e5cd3dafa13190675;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5948d3d18e97eff43e3d282a940d7c6bebe72b81236d5a096d7a929936e42a503e4c9f6c811223f34ae3a21d88349c7e1ad85413360f727b92b77d14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc09f9a8be07d84edc0119a4c655ffb28405b29183fa669493c68593a03a7fbc8da9b1cd9a322ee1e54b76fc935d1b030d87b2b47719ea6207a06c8104;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h134e33f6659a389d4d25746ae3b6a80d681bb4dde61a98a8a8ace08339a8f6c89532eecc1b92a3499873e65dfd964ae6109875ba5ac025f16f4cf4ee0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedbc6f534155336932c08649ef6e6623b24e7bc28f5865b3d63cd83601d458e1959af5bee53091acf456a62fdc7c249c68d951810c63422ccd23ce4c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b25b72fddce6208f5d81e4b28783825dadc8aec30105aca2a6e0be71a3a60be2e98a42201b0959ffe99da0eaa754733016dfeb3246e9216c0ca04a74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a5eb467754dfedc97507fbf299b648d58062fc17bf9d9786693a188a9afa873541296e07cbddde61c1aa722288bc459bacba33acc2dc93a07ca12519;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae5509e53c0b1e64b7b61e1136aed381e9a6d28715137ec89c0d127683145d7231cff51350a8546f95b04497ea59f72abff8bf399ca65f055c3c71707;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc01f81f3a9d1165c4ada77f0c8ae329384ea5a399664ac5076363c52944d61ece909d9deb7c686e2158b2b1a3be6b1d256983962f408cc67d676f3f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcf193a6132978b4360af29e06abce1a3829043623c6e882f778acd9f4d274d83dc8fbf87e17f44bfebf68403fd3a5e2e21eece29c79ea323b1878818;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee916687b09664b271bfa1cd441a9f0d4903c98730a93a26c536487aff299978acfd4a1e9527f281ce61cd7396f08f7a725601b7ebf996fc7504e698a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32b3e0eaab41d1d4fb30ff94853411e0fd3d288376fe352941ad36c1d558d626f8a337764cf280d9f092971f14688f1123d1b449912c5d5119b846079;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30080d69be6405e012480708d806497e404be87a494d8c505e51a96c35840cef1ec8178c60a1e8c6a4fdc95b71aba845fcb3f371a2205ae4bfbd49b88;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d477b00eaccb305122f96e6dce7c9bb0eab3c969f5386fe5ae6616f583d7df06c4c71a77a6d972d7428ec9194ae3779745498a574a83ead4dd1cb185;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h152b6efdd5641fc20aedad531a290c3f9db14c5f0230d13d7529a76f38a19229a8f734ad2c8b3bceb439414e189a805603d8ce6bf513bfacc540dbb20;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca1b9bc7a2b28109c3ac70b92b2509dd607adbf21407930498b34bf9f02ae179bd6fbe7f91d1f63fd0b85632d540f95982ed7d07d523b0c3a8462f8e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8eb154106b98fa614e541fcf895576343e227bc584df04749e03281d81bfd560ffedabce65a8b20e11787667e0b6b16a1d4051c0241c0e306256c987b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fefb16e567700fdf49153f71417d3af45f49fc8e7362db1bc5ed76d720607a434018b1732d981ff7e87be36408b80825ad57ec4905b09ffbd4a390da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h412f524e34cab22f763edd658a7a221bb57c74fcd5893516b5a3bacd34b83a0480bd5bb90887a415d06bfe345caaeebf0836284c21a11f5ba60cdd780;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7809f6cc62d485073d2a60994f117f3d971a09150f93c52c0f5417fc4dc2ddfce238f1cdc1e24ee8ab9ac909966b9650ae20d7c48b66b361020dc4d2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72a249949f4683458306baab5735be2b71f354bac2c0803bffb0826c9228222e054276dd14129de024d8b170573b8f4236ffcddbaf04d5e050e29b437;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h209557cd841198eaa1512542551352f4fba483043e81ea4ddb0e818ac887e12d1d5b409d43b03678f4f9e369af50066e969630fa6a26fdaebdfe334e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3289c9b14ca02d60abdae58c8457836f7b34ac28bebc891a71b517b040759aa6d3268c528a326bf3a7900141b09fe7bab9d48727cafdb2b0e60a0faad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h381ff60a33bb33fb790de487379cc7db33016ea172c4d101acbe5c7836f308c1e6793c1b2b274bca5c84a76464e9fd25d4582ec506178da8b177a3bd7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0b4acfd8d0b88c54dcdc3d616b357583d2ccbeff38b958c61a8315a5042e7de6410b923a8ae9bed0bbbc89d0ecd46c09dd9d0bba94a9924742bcfa74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cda2b5339a63a67198323c51e32a9a7354471497bb1fcfa8a72f843a06bc1f4c634a1c75970a55a0af79cbae02a2b8cd5c7aedb907d9ccca4eca434b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc94eaf89813fead58905831a6ae7e6c9ec92bd219d029b642f06ae03455e46af9cd4906292b55d75913b681e6989539e37952d6872dac6e8c270b7f05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2bb61077e942d5e2d350d7409847eaf78f016d37bf6336ee9987619f521c37b93fcad686ecf05bb2fb08c06054d208d8c76f2dba319a2135defb2d67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20bc22315305685d1584b1f861bbddbe0dbf94eb266ff9388e726f2e30a99cb3638cc03d7fff667e94dc898f5a2f94c52861dec0686cd50c4f68777a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6813b11636dd15b2f3b6d35ea74729a86efea04b6f0534ce0cf98824baaf2295ef9aa5ca9572a2cd92381ca8c53fb2aaa8e93aea5be31d0344143d041;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84020d98c7050e17f948187d431acc2a097887156f4179929b21c73b80c0e1b3f02416f7af465304fbb4cc213f2a1df837d40fbe026470a85b868289e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae02423d520133f31cb1d603d35f712833abd2ddeee4cc3908df7056dc79b54dceacb0c12efa749df18190b9be06b47fc500517a0e838fce1a0716b3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha107d625d42b6de215f533b59099445c5136bc75135cee631676bcc537c123014e279c763ffe61dbdf92db8e3d1be70392ab619e61bb56152d2c05f5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b750ceee3aabead92f6987a7643909ac228445e64e648a681ab8fdd29e459708f718dcf3e168744ff03d3a0be786c3ec5fc61694d52155154c0c474b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35fdd1fc5d714a11679793648b292871ebf189046d1b84701cceb1a9f905048c8fa857486fa3925f2b83495314aa3aaaaa6ccc83bb0901d0ec2107405;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h253b3aec6b0b2807e8bf31d12c817157f77c69cd08515037aac4b19f66ab9d2ab4f41cfc8acafc16f0a5d2fa3eadedc16f45cb1e378db2fb49138c5bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19f1a11dcec979f070356d5b9f946a0355b999f77667aa6f2927a0d52600bbb971998b4a205e69b3e3fbd76cd6f9014ecc4c7b5b0d02c0ec30477bc05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f24bf0d51f007c71ec2d5cf163bce3db71dfe3657cfd01d7f78699134896c513bdaec20cc611ace0f10efdf63adaed65b88c9d592de6e5a2d1482a92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3d9901053884330ecab0923e188bfc3a10b5dc964e1129665fbf831d130bd4b36b009c149744841c9cbc869022d164ba135c946aa8e9102f12f045c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h262329ca1fd6d8e0468b91a4e4d425fa9ab9bf45963d41a1eaf574c43f249896ff7ac49b57309de28a59f73ef103635fa61281a0be81c472b45d74700;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h654efd56b8e43bbf7223f608ddd2cf5b90d446188934100594e7b8bb599bada70a714a5884aa4a5d6597d243ce4e02de517d8280d73c098d1e99c35c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha199cc41ba6bd3490e53768d8fd969dd28c392324735cad5bef922cc097353a7fd1cae9bfe665d945c42e0363161790571c16a0c28704749cdb800bc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62c7b8a9e892770cbe83e6cd1b14906170ff60a68e3a4f7af37ee48bfd08a40f9de3d2cb8baead692303b31aba8d319771e559ec764ea537a062d48ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe79278c329ed5c541b8c4bc61b04518af82a409003efe4cbfabe41b57437d7fb7b85d9d7da67ce6794e09df5a825b023003b64708039979be784c811;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c87802fde4e0432acf25ba981c8fae87bd90bcfe167a291fe326efa817fe67444e957d07597a596040cffc75439300b06495a695f3d277b85dcbeef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a4495e617b1fdfacf1cda81d4efc8ae154d11585f07222946310157bfb3432c69f1737dafce9d5b673b4388763352d31be8dd02f55ab3efc093ed89d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8e343b6fa043756f6100bd13319f17ade709e6954de1b84bb2d4cafa1fce3a41b0f805566114c7db25affb922d08a00eff3415a9cfa9b430b65f2172;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8742d89171b83a46ecb728e2deb1c158dfd247de7da180a08f59c81859ba84b73b5bc7a4597c55cecda59437af09f3875f780db7c2509bd812b98391f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9881c9851f8d78320a6b107a1e66065fa28edcaf409cd58b2bb3e2f7bb57b87d1ddf39984f237f5d77e9cce90839bf0b1f05a8c61821f3bbc52caaaef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67d51caf59b78691696349e04eb239e4ce17b773843e0f27c414d94a40fb4653d333d78b03db004fa29c322ac4aaa84da04863262ce5e01b6b8cbf3c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d36c22486b3a06c1ef581603e62fb1b00ff77c045e1712389bc2c5dfe3f0ed6f54e10811b9ef3fa4810e9940014786b7bf587a1584fb7c33c120f9c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he592b420a426dcab8a2fa8228a5e6021d34f1b0ee6ed3c92ebfa6439f6872c4fb47ac413d5dac50ee77d38a924aea3e16016dd339ff6c76fd0c5e6a8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he399da761e84edcce3f980e289a65f85aa4e017e02c9447474cd785a25bbeb810e6db478393556be967f1d7e40c04aaff6527404702ed29902126d8e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haca7b7ea048bcf17785e71aabe7d54f489a347707c93e8315a559e77016dc60a474f777cfdac67f797016f7238653bb22d0db1ac8e5c0aac276b13939;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd51a5b690a87809541fa238d4455591eb0a4fda387faeb2c143941917d13a3b078bdfad057560cf381b6299b6fa00a3e3548f010b951ef435d90e118b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f86965c618b7cf96ff0c04f707f4208f379c20d35699a8f95ecaa860ccba1d4a166f2b89664f7f15ab691ea317e0fd3398dcc8796172b2ce8dd7ce75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98a21abdc0e0a2f7aaa8b4c2b6b56fb01c6dac988d6d7d294d3f01594346a15b4d7f8f226fa71ffd3098c3d55d61ebd1f9a48d367e42dfbe3a2544a39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c7649bf783a65dba4436b061f52fc450148e356306f0a79cf23c4f6d918626d296f18541516c4eebb04f33e5de32d399461af08f83804d526302ea71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h757148d43b686319032ab2084f36b289e8cfcc364f50fe6d7f7e9fc5aef6b3bcba076051080a5278b4cfd8c00de0b9c61a4bd6d8032a6b5c458ce682a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62323df07c938dea8c3d5d99c2693bc086583cf5ff7166b009d2ed1802df83227d26e66b9bd73b20baffa706f48ec5ce3a93d996e0296430aee484571;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9815aa732be52f0983494c6ba4555a444eb5603565dd3b6885fa74bdf3471f938b3b2cdb0527768564c6b020933c787411497240a7a3c0b372ff8d501;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a139ef261825d4d0c7c794c3dc8d18c20c53dcbf4036547e014a20f8e3ccc77ef537997cfdcf822c2901fced1313a40b76c8b394aa9ea65298e7193a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd945db3d6e870522568cf79cb63a3d1c3dc57b33fdb0817c6bfc7c693c840781d964966df21546655f2b7ebb5a05904d8173b024066283808b6eb0213;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69005d973724b11b1fd059c76ae095d76d90d71d1293529f61157f3f8a61245361a76e98660f91f9c661b3b112c7bb727a08c67f70e4cf195871e5faf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59d2700a5fae3dc76b36f7c28f54d38b888cde60f5a8ddeea586ae75d32f115ca516afd92c54bcec717534c347c0b84dda5df09324ad023b73b0d075b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd5e7577592af31ef5d16074530b437c438bbe2c8736c816244723379de534778d5a9f84b4bbd3bdd33e810950dabe293524ead09db611d8fd6a191f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f1775346408b2d48cf08e0ec24dd3df59cea39dc378c9ada042e58648f46a9651ec471e84f0eadda7e5b3daf1a576beabccf45ae821db2d97949ded4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he12bf3550ff247f5b710652ae417d08e371d5a5955ee237543ef275b89206c7aa41e830528ab55b885c5d4c2e961a5a54f872f0306562d7b387cbd386;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a26c7cf8209914a1c767cb659af769ca5d1610def8645f6fc4e4362ac5c84c250103be296c6f59f0e5c9bf9786118c44ce09d143ca1e1bff0a401287;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2430622c59f494074af2784d6e4671772385bbd9b76ed14f655b0cb600fecd6d42bc5e67c3859ebb69b7cca581b07dc45884d27a929234d07b9df9381;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4487270e386316cc6a1a13b69c3cd0742d8d9f02d27c6415bb477ca61f64965e9fa81553c9c518a2d67bbb86906a980db8ee20b377872761c4044d847;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45dab576b57289ffa775ea755c47e658b9ec22e8780e0693d4d728c690984a53195d9b624fac6fd93255a7be8bd9e0b190c3553fafef48b33c56be27a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb164dfcfad537329573188c1a8f75705ef57aae4d76af0c951676e9c77f22269dacf408f260f910f9a2f13024b6d0b0d073154476e4345b0e3c270137;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d1a30702af2f44680eefee5e04f0cc5b61b1624d408764e50338f3764484b6521a21cb1eb1d55080e48e898d836ac0184c7b81dac000b2c462f730c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7caf53006406d31c1aa8f2376dfb3925e3ca4921a875c0863631ffaa9aa5c4e814bac84f643e8c75013768bf3a3fb9a953beefd31b5e888824990c493;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48a4a91b100dfbe1d61f76c64fca664f643c55cae60937a7af16a7295e95028f3024e016c5fbc81dc05e5d4f5b97735d7e1192090ed79099a6161a05f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78922b5dda008b28e92d32677b0c5c2fb7338dcf8314e6fef7b9e3d87075a3469df86bb093a083e7afe7d838e0a03ede436b8dad1e4ae76fa69407f6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h744ddddd62f16ffcd8a16b0d5d012d0ba1b86013b2a79a1da8e51ca381c368d9cbf66162f75aff358d400b251d47b8698c0a39e3b1a55cffd3ad9660a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26d2472527bd859f9d5419bc03204b933ec0302b918c9c85829064d1e55145cfc8401b269d6f31b40e6eca42473710af2bb5eda8d9c94a0531f618cef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ace70cb70075f5c6df79d2088f22a33ca743d156727b5523d28e11f5ae3c18c8fc1dcfd18e6a3dfcae307ed6b0799a034f9bbb3fa3e3d8cc10abdf3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he07c1816684287daaa2bff44ef408199a5db5079783483e11c11d504727b711dba1a63f0d0172ec5574cd24acaaaa4dcaaefd1d254a7fe89b8b0ad44d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcef9ed6c1ce43de95d11fe6a2b923d3d16ff301b35a2e3964c598545a6d868497909a131189ac976db68af983382b4b1f368db2430e03bb050f66ddfa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ccd64089302925b711933072fb79e8fb523eab60996a6f3dabb82804ae03659d95019b49d55fd4b4be9bdc28f3e7e7a3fc6725af54f83b9bf3d8aeb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dfcdccf7d8cb218f629a85c7e330fd8e30e36a8404d4c9a57c004e155e2e7c0dbf9f7e55eed4e993caa419b3deb0823fb03311049d5027acc67981c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f69d68a03d06948f164ea68511b94ad726d811892d2c21f14ba7fe704186db20b81c136ebbac737fc5707a2036cbc9ea2eedefa0756d933878d43f93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h648fbfa8a9f2b31b157ea5fb946865d92a00cd331ad76da15f0fe6b425a1f40923f31a110b03210409726b8481fbe64ec19a72a9984b47d28fa3da514;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfece64830b49ae8c74e8bf65f2eb05f934cb8ba6e66738ca47b89f18f38e121531e4cdbd10f4be66e7452451617db1982ca00078a78b48026dfde6e35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf05929acbaeb62dabf0793293d7da13593d45499478c5b70f249ff3bfea30ae70154ec246dff6120a01a63d9591f5a6f3285522d86a71d068a7a59779;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60c2bd3e13bbe932612ad96b43b8d23b53ddbaccc658b2647d2da284c9e985a8e0ef134d79465031096e4d8dd2d9332cbb7fb332ad14ab04d9ba054c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h919466556dac29bdfa856e20d5d81bbf8376955961cb80691bff804a1c64ab39eb591bd03057584bc8faf3bcfefab20de98ec9d3ef37ac4d0f162ab1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d0ccd4b238385ea2491922ab47315dacb2587a99b08d685beb0984bccf6bffc924d2571b6d72d9d057c1cfa5ae7ae4468df41cbd14ff6577f3d185a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h755889d61c0032873759577d3e1878faa21684979cf7ed336a8134a0fa01649de1ff8865d9721aa840316ff37bbcc011843e89bde01f65e2454ee2211;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he41042dc46a8349a5e738a45f7796ba5c91c68a0cc0d2d0de2d815c547bf02591de61704fd18ce791606cef89a183468bcf90fb3888c2ea16c25b153a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa5b13a471ae6ba470635e5359206cd14970ecf869f1705ecf9c18ffb58f7cbdb3bf625587b4798e3a538f63cfa7fc7f1592eccf2c00a96719728e886;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5f9174851e23ff75ccc384ada7876eab32bc1f8cd20dc58890d90495bc97158ac9d547eb868c81c783ab2b42f00718c646df66280478d996b7a2a795;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha419d72ab6252e3fa21c9d33ac1ad2872b30a3afaf2dd298507638b42779a08350b7fd9b2ea879f72c7feb6b5e1f044467b3996852ca599e357563d2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haeb28b0e69cbdfcf864c048400224635c71e8f532c6f572187565e04f645331e784e41090c0561096e376bdd7332afd5019262fbcd288e26681c62ea4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha18135fc29862a385705c7606d659b3914e0f1c0402e9e8163d2a3d310220cd9aa7c832e0b828adb38db3d649daed071e5f3f4f9631a58ec501eaeb76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6baa79814ea0165801b7243e53da4bf6d1d4d1d206429f3b57025cdf529296766a632a8efb790180d9f18797ad774ab0d666a942e6da2e74c308901e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc08dd1fc0eb7c96953ebbb3f7c8cf3f565408acec3e524c310579170d198685dbeeea498461eebb850d06fcd5a59a22e1bd1d1a83b8ddede115ca3b4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7b28615843c7d7ebd503a3a2fe24ff69f2de1e9010d7e8421b806eeb21aba02c651f2bb405aca08450d95f51e53866e4e5da7a2831aa0954c3fd1b14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h431ead1d66aa6649f538403234d4c36f02dad421776ca5224106e21db65004c4d47ee3ee9e5bbfe2e4e6e8bcc35c5f4ce3917851c3fa7af7f67d82cec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac92499d62984126395ee7c3626303f6c796c6b8e4d0b306df4cd529fedb2a33572af58ef5ef2d5a79cf497fdbd6c9c3aec4147f1cbb5c736f2054549;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h852586a57809a50ffdaa6b7fa7d971534e0e0def266510938ec497961f32de025a2f5857d30853e130c604576315a1008ffb250e069bdd0ab7af2914;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3af2a6d946a9edc842c04709607d62b7b90a545458c2a4f34cec2d96de27cf5d69e45438653632140512888d602ca7e88ceb498f0b03b079d241bb2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h561a2c001692ea7ddde5978e4f1695ec7dfcedd5260affafc5bbfbe56d54d5ce572a46f7dd99ce0d6b7608664c9d571ae426891a8c3c627af4505f43d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98ee18080add6748796e078a5c1bacc4841b0fec4a8af7773b1af7d5c3fe100ee431a4d2fa1c0479b0cee27ce3e7b64f1ded806df1c4c9d5d32d60881;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7afc3c013dc5cecd4b81e19f54d0bc8bb9999803e378778c381810a0828b39b037c5a60ab67a0901292a0ee735e4ebd336c28c4a85200974dd26dddc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4443d20bb55e3def041f742110b68e531f82807bbc0fd1f8dfb1a379878137412178cbdd3e43fa6803873fa9da2b2f11f9bacb140a0b16ca2434d9db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5deed3a1e2747021f1369e98338df8397088a241759da1d92a8c35280748f019e201e5860e1f164dbf85627c22768d8cccdd8968eaf051b25318724d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0d53beadee6f4526ddf395d45532360aaf031f389d7df7d3ff422b94456dd30b83a75ea22bbf04a1cc1c16c19ec3412421b530faa3e7670ee8b5cecc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29be81bf911a4812bb17b37423d39b77838edbb73d33c56a5d3837e6d8e3ff1fcf5d683225983fc8e92fb9f4d30cc55f4fb4b13806671f28f32066ad7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76bc935ab2d2418d53e7b1cb668b974c669b1dfe1f80df4cca22a2e8021a9eb333771ede397c6ee481f602d21135e51a437ff84ac4beb127fdc53b15a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha82fd7c1c6037c1d46f964df9a05c038d0a3dc21f8f40612ada531647e9b562fc821649f681d1e4d0efad4c547457a154a6d8b357e32eca9daa4c18f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29a033ff78d58517cb16f849aecaf4e02c92eea065e96ee111babc9afd1c4dd763144080a53d037a486c4f61555b2854023d90e95765cfa3895c07f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f3abe3cb960917bdc1b593495c970ee61e9f2542c14bf7c640a7c67b7ae6810856df4b18aaf97248e78268ad4501ad8dd1d18b5859318ffdb78f7abb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf70afcc2ac28a4404de6e64534739990b509f87127a52b3e9f306b0069e5474cb1d54f8e07b248ae4d1f9b67c37fb9cd3ec87270cce66bda6963c790c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb0e7ef0d465721a201d2c5f841f1f1677ec2ffd65a8f4fb0c85cce191e3858a86e103c240feb1c7b331867a28a91ebca9b020003f937813f993e01a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91bc719c18914e350328fce4ae0b1eb04f256ab44a2c458092d9ad04f7162bfcb0282bd75e653ac8de209178a6643fe4c7d8cc5efa048cbee156d5529;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h805fb4c4d23266643728c4960036e07f706db8308842f76cf5c347535042ee43c99a14b41b03d357f1cb08f7ec8fd81a727de78005f1dcc59353232c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d728a23788865f93098d2f546a88f12502c6685faef0f69942d46f37c31bc29984ebc2c7d368cc46ddd8d14608ad87453fcb8531388fdee77af9d1d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1da2b32404549e39ed259efb7d6405755b33320534fa47eb5df91eeb76b8086add8924f7830d572f400178153d8190129ddfbd4be326d18ed64f6344b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1267ec22022b719f7790289fff400eae36dafac8f69210b5e41a7aa5b3121fe320fc39341cf41c36054fd7e5e856e8ece70e6613e157d2387fec11c86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e291203834ac332f28269a55206a36edaad01d1f94bc1db6993740712dacd114f8c4db022e15653645e8a738ebadc28c63cd6ef7cb9a97f307df998b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2028c0be88e2ed4746fe166082ccc63d696c5176c50a2d2db390f5d507fcd7b8698b0c0c3e79d7ff0ad46f5c47755beb4c5afc71672cff4311db48c5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48bae171debb5c42054192305ad668cc856c21315833fd8c0cd73c2bf8e0015e4f1a5646c8df57c4bb413970bcf8aeecb624d02f0c6d4fb8c22d04337;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96129cd67836a9252136bc6fd539006477e87740990234fc6ddf2c096c13a2011582abcea4d5097ae50d78ba108547130704efe65be0468cfd9785604;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf72f8b3c836ad1f3307d06d622e536dd4efb1ac4082aa0d340daed31031ca57f13e70d7c8d3f3ccd7b0ddde3d91cd5f005fa95398dd047462d529e98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he95a0074ff9dda779c012cfb422b70fe3fc879a01d428489df930b601a4d4f2ccc8cd2615bd339a825191af64d1286b0d4c707ff744634a48b42d5e7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4384f8729b1bbc3a95ab51c0d9e0a121370dc5c8de96f08fb4a42336a782c7e57457a60da854d7a4133853a58f1994f75aaef1f1394ba5a8b4856b9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7925d344a0a63344d496575e5ece3be3cb6169a95d035aca1ac6fdda4b4dad5d91f5d549e275488d8b1f6136fe3be66b5bb8f2424be2cb642b3af35ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h623fd03a7083d46fe09112c69f7321d9c671ce0e4515ae907fd87385c34c1271d98c009f8010a7b5d6fdd1ba3c0cb570ea1e738329c6d0f087eed257a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac36238b3e544c42c3596ac7df06735142bf7be08cb08ee6682293523707d4c6fdb8614fd0e49dad49a7e39e357970744eb24af5e452563a8172367f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha05a5f5409c210531901d342f8133c78fc08ab199d09323a18f963bf8c262fd058a528c0eaf6c4a7360a5034e7758143073e07e383d0a3da3c6f633a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc364b5683aa31fdd4e3b6f7d66f98d82b2ee7ac5754e9ce31585e82c85af1bea0b1dd01345232436079cec6d2162dd719e8c3ca7024d5169e32ba6ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h893c3c0806b25a7b168395e94582b17613c312443117744cf34004e76b961584fb73f341d3eeca06033ccaba777beee00e5013bfb358571b81ba065ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha66c67009df19f6f60a1685f3eeaf33a3f405b7e1b6c9ff3f26724b0d26b320b88c8082533ee9acba807e398a76d11353013a7160a3c91134a7005bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he112545c4e5573017b8f3d27b6049adb23ec579b41ce0bc4df10162da6869bc3bb1f99102b91454d63cae145847d7e2da038e6123538e6b13a5113bc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d166e3ff94faa2bd87f30a7e59201ac90a76a90c8249c5c720fb64560f9fd3d875031c552075d79463c61d6aafe07565251bdaa0a6a1414f13a192f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c3b65b1011d772331d8b6c323fb5df53b507f42d4ed53c0727e55edad2784783ac91ff687a0f7540a366f1e8057903b5dbdfbc21d02d98058066db7e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h292bebc174a9d4d9efe525bd65fa0d184d1725291dd88da6c3a018c577effcca54896e9e121d82e4f3042eee35f68bd4984a6ed7ef4613839ac8cf807;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h719243f075636ca6046512db15b2ef2109f5ef6a1923cdfb4228c7a086bf7ace4196e423bf3cbc50b1044ea76271e579e6611f1c4983a9a9787871f12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33607f26badae6ca29c7727987810c4f7a5703a5eabb18b9875f87bfbd0e10fb505b2ca51c23b28b71089d8e668d7d797890d9e2f7d82982635f565ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d66e1dd17396f8bbc6f7fd0bdee05701a563c401f9c9e4977618a5aa1def0a3eb1383fa44b0b40040d7fbf82928ec81bb12fbd54f308b6e2980e50be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf26e40ddd5772718e834bdf81333dbc1a250dabc40e929dcd6e3e48da095c5a656d25bde3f4a3b7b1a5be74afbc2ebe83a5f6dff5c1f471348b8b39f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ed7a76eb827303eca3eda78f23a7bca69aa8a05dcd8310420071b1428d81125a6004239910e34021c831ceaebf85cd93ba4221258628a66ee0cd661b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3151215c081a895f715d86e80e4d69e9b6d011cf59fc1506d765a7359dcc129972f3538a289df9d54d113e5780480116da03f0c6ac79daa76c2d6e3b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f8693ca59ce79a16ecec8c374e6a84a9ef170ab01d1cdeec28b1073e8259af05e71f7efcee6491882b8dee0349ee2e3a925397c26ecba549dda919b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25fa2e60f535282133364a1d08aa141045053acacf72375a1ef72e81ab6190019e7de7d0066237d66750ca929b58394f53dc549c2e5c051a3bef0aef0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc23d1e452185a438be794e1d5bca4817f2941304c155b13bfaec9f7ec0bb8dd5fbd080a46748acc3ed276cd26039e17d7d4eb23279869a6a6f56d9091;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfeddf65dee0b653404406bf240bfea079b013cf1935e7ac71ab17c09e789297e0d6f1e67277f24493d5ffccb559b0008d6ddf1295d2ae1e7a98ddbbcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44d4e69bdedf72fcbc7d4493c70844d32d4e169aa71839f3c18668a6d4fe5327de48688233f85bbe712315ef49ea7ac494d07476200d172f85ce3c3cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d8bfe41bbc205984d3363226eb7bcaa714657143acacb2bae05eb17e2a05c7e2a073cbb4ad94fdfbe68d373176172c87ad07e3c215b906b154caa92d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99aaa60b5ee7a58f7fe785744f30698f7aed7147d0ceba43bbf1867f04ee520359561d4848dd96ce66494b6c9927cb396eaf50c06e860a9e7c5c2e6c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7521629bb5a7fc1764f048e3cb7a4b6b38f024b3b6d1ccc0b24a76d49467a81a0c76127bfcbce646e88e9410c7d17bd3493e4c3eb0e5256f65e0d2da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5ea0b2cc303566fc22ea174cbb9f23a7a05aec1187e0bc975bafb7c53d83e1ccbcbc0b52f3720f74466879536b0cc7a3aa4581a5bb2157c7913b222b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91e415c2f6c3f993fe8a7b6591165150b1485c4037d8774ee83d767d9e9fb1b364f172f3093c696bc65eb4b95f5c382b29fe7173d1f6883f88bb56ea1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96efa586f907f070735f32c9e84f09502cf3b137425575ed2c6bb0bad3d46086c27204c6225a379ce93f9e1e2af07e7c1ba1c24602f0410520a0a1115;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d2bf485ce18e8f034cafae7be42c068a643954672c85b2b64bdd3a45a0329673ec921fddbaeb52c333694b38872febfb85ae3fe3d20daa91790d78f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fc9bbdb8ee12dae1402eecbd5da2affda8ed1b297929cfb7ce0ea99524839009dc96e00b407ebf1ae1bb7acad561343d7deea0d343fd6dd13adf8847;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51d1d717cac800461d38ae585c4f8e9d9bb389c33bf49b923444029b6f91325db94db4540cc90e7045dd986b9983afabd09a955ef35a1715d930b0298;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf5a00c69def1428f2d025d54845e6f5f9d36a996cc1665b631df9c9f32d3235ef4e510ca128c6faf425efe3d35d2f82e4883b7a8fe39e829b3bc6321;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48274fdf6cafd4bd36c402e89327bf952ea8f1ac749a16771b2e8ad40da70e4c08f6d6cd285c831817c9fa0b5a45325bac300aac4591214999b9c676a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb35e8fc2f7c63216e3de0cd2599d624d772af5eca935797944ed9336a51a1921239c53d5a2006e6b5b4775315cf5c5227a4af26267a2a5e77db28d8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54b0add7d2365b15d4fcae35393062514cf02921395f30d3117f91be2baf9fbbc078e30758154147a415a073605090384411bb2f3eff5282848d36242;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb169dc9c3787cc277e77cc23b7d8d5b37a4ca8968132700b76a0ef6a4766eadd3df0636e7c48e45e15583e9ec9c03e235bb18e223fe03e0da1bda53c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34dd8617002ea610b1e3a545a8a0a7495a083d36eba46404e49b51f32fe63b65d6dd09db60ac9486307f0d3e9821a19fd29e740f10e5dcf2a61231d58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h535043193d2aeb6fec6a0639c46e0503dfde7afa0f493604440d1faf3f27793210be90685884f2e6e17b2dcb394fc8d7002f9b2961c8fecf58fa4f7e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h413b5b2c5615ce98dbca7fdeb0238ad502de14024cee42330d2a4b0f4a803cea8ee90c6c81ea385ad89b1fb32b2050979994b413682bf6fb73a5a8f8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34836c05e8972782e4e7a7001dada6f0955e99f1cd24b6e6924267d525a416cd3b828ef6e7baa0bf18f56d62577bf9f9e1b7d21e18ef4df6ace381771;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcea368060eae808206c188fdc5682e7c69aac9833d5a102a3c8e47c078bae17b4bda807daf39c6f3274f78cfde2b09f7832e433cfda00a81429ece227;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd95874dc9010a8aa221eac9839c3ebb493592b06847a6b7f9e19efdfc845275fd34f316dda18f56fd99958e33a8ec6ec131db734c55a197a400121e57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9d77ff38636ec372a676a30690db9694aa4a3214adde5a71e8751fcdba48d0f8bc269dd145cacdacf9db1e4fbe8a13f19f2ddad168baf3a96886d730;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd17d13a3503d728682d532109aac4baa72145b12b45aad969045b5c11cb6b92eb7cdd9dcaf1f7f2b12d15ae662c37742852f900b3d2356ecd6cc6bad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd216028b97168948a7842560e53b012e158e3d4293563c6ce5cd8a4fd6f7e8bbbb7012f86217c48b3237188ae8242843b013e5c51ab55befd71d4ab6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cce04fff2575723f93a4f74884b01fa33537159d68c0618f02daf46aff6ef87b2b8b02c9b56e2f30cb9781bd56d869bbcdbfbb411cbfe035bd76a52d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90da7365afcee45e1b5dbe1443a74d91b65c2719b3b35fae1cb2a0571d2c6702d44f6901147f9548de2a4943ab0b1f02a940f78fcfcaa8a7ab38f3fd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6fdf8f7879800256eab62cea7522a42ff79f7dec4b7ff9623b1524a9f222ac617f840c63c45b3a1bd6d72269fe7b817c0d25d8428d15de6cddc36102;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ce641782a91b3cdf52cac051f65c7cd45ad0e19a75ff05ce6e7a212f8ff702522c51f1d8ba6576de3788a55a9658a770b64d9f0b6b8af1f8a0a8755b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3578c4219b1b58158f51aab909b8f34fc757a31fe6c54386398fcdb84c915de07f424bd0f97df29c25b290a4c7b68186e05606a3797662a748da6c9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h154c5dfd85d07d552a3da090e55c3dbe6458ef1f5c0f3ef5e47698f416eb496f5a723e20cf00da6fe2dab653ad8cf1a194862bb5d8dcd5c15c5f13b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3f4e09be27d21090d6d43e6093d0083557d29b260c1f93818801743cbacf65355178a0d0eb0912ec7c1db43ce5bb2ea1116759f7cb9dea9698bbb8c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d0b8c77f94c4d13bf6c034cd43d28b82cbfa0dd697ae6407efcf1c4b02d35517d125bd4bbf1c7058cd83fd3b5b66eea53d11d195995bb8255972da9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h756f22f972e97603ee0042651aa1937613a27e117271454f58e0e314be55e734f813c0ff4b2324729faba5e4c0fa7bd90c147fdf3114a40df53b9d13a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd76d3151af3a1eeb683e378dae1938848e2046e37c80b5e593fb391d5bb690af9a3a25a448d96b7d1562fded033e0a9e7857bb62a6e533b00415390d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3422b081fb8ed12d3dc615a889c7b730661252e5b5658ccf237342486ae43fa8e94f161e4a254b34e5ab06ea76860710f8f06895a3952045d50f3e3fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd23b38a8581739a178bdec6998fb9e19771c4abe03bd167e944d2ca14c757d9cd0ed478b246c430a4a4c8ae4a599655e25c7958e92bd0bf3e2f28d7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27affd5e3487e883d14e69ad9602fc242cc2de796e915d731c3d3e88e8d40c0b29a9cb5013ddd450b1b04fc8af08e4bcf70fe7381e0e0c41faf32483b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9bf8cebb15b72f3813309a78af395c9adf0e52d1ef38c61508c97d08c4e4fe70d9cd62eb7626c4dc65e7abcb60c563f92d7bfebe4d9385500e30f8fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff21da1fb4a9bb1da0eb13f30fa31f0c13ab8d1e7dfd0743957631d4fd990de32fe602099cec238d1427314202d48d3711121362832a6ae30eace4c6b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5aa86dce661d735810a2b0ac417c694123e9cbe7140febc36eb94073833b1ecf1c1a3a1f05f72cd35aab3c80cd01ca7f370fd0dcf0f90171c2abc9206;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8c35b5ee1bc128b4fe01fe52e52e4ad93cab64a39d1167183672345ef285eca78c9681d528e9c50141227d45042a86e651bdd61c4f0f55daf3de3001;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h137b7040ec675bc336fd8f1762ea776904a9af99831aafc82cb1355d14bbc682dc896dfdcf07efb7ca898c7172331d1be89a44935e51aa313363d5bd8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4113b294bfe52a9c0f8eb7bdae08500d8b4c30d534a1a3414f0fe6ceb5f59c4de9d87bceef038ebbc44bf97bb2c6df23ee809db298f6a20f3e379b684;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44f8fd414937e02dd355655371a400b6a7f753a8e3dcb8b9c0ba0be5fe183238d66fc9660143d436e9833864f8f237af0d95eca891770578e37340c9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab68678d3de12c462b5b44a19cd6dd7fde51dac74805bddc5c8275cfcfecdce0a8528f6ec1db01757d2901c8401d49d50c82d7f93f315d924b09b5642;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed3a17b92dd5427d391ec0a138a83a223f51fe8e150e3cfde713cdfd53ba94b35cb6729fa804bad3fec77718f06ec0103740392b3a379332c12143a1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cfdbfdd980f0eb4e1e19bd6963aa1b1595754bb44bab353b6e4296350450e26da16f7a484daee2e7b489f01ad759a660a73b8a817b6e09c749218b92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf952bfa18779ccaf3915cd44a134ecd5e45e2acbe5eb7bb18c365e3ff855272123933455483499e312fbb9326151dd51312dad5b767ac993baf40f32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8993db1406bca6b87018a3fddfac577bc0d29fa1cb675701a47af0797534d01879eaa3ff7c01d526495cd8c3bc75ac5d7b3bde12e8faba2279c47528;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86b3b0299101dd8eeb615062fb794e5b06190d2e5345a1696077e43dd85104c2eed88303bbb2015329ed0e7513b25e92f9bb484c3e55a21f81e7820a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24601e4d2ea7509024b2f4def32f3c71ed5b25f9553e1ae95ed9770b975cb0f9f6c37f5273bcb34e6e37c1dcc0a1a873c68bb56de2ec01fa882bda938;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb5e4c71b39ffce80cc3031daf265a22c4fa9c298af5322146b337aafa19742dcdb5ceefead664426c75f9b25245b5af4caee0925db496429e3f6431c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4fb2450aed30f23ca580a78ea7a6409d0df389803cf6471259af33e26c5857530997e7061971dda84b79ee120789674344099b3be95d7964a1d2fe7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e2a330cc38fa773b8a30a7fb7d543d6330b8f2f0459ab64a5929d9adfc72b10774a4f410790f7c93629ef6ed8aec60b600fd259a0b0bcc73c91156d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf3c7cb3310a31a7f255c8cf3db2bf9bf47548e6d612b729c722626857e25d5e4244cd41146d899588c79f4e54ad6339341e8408c2ad8328fdbde4bf8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6847b3917528b1dd140d6b0a323469d4d4d2483eabeca202f50a744002e401e952e03412c8e628e7480e22626a1accc54f4175f7e3231707e8661c065;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff797b6b3b74984ed4cc5e2a66aea3782a07b1fe6a0daea75610eb7359a9076dfad654a82401e13fcfe72375364dd7e8a07eeb09804752cf39c8fa7f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf3f7c0cfd1d06ede3c1eb4edd9f1162420918be47fdb62a65075d08376ea2e420aea27f1617e343d66ee18ffe357ea31a49b7455a9a651e9a6d048b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h475e8ace7fb0412cf9101129332f0fc2ed4f8f1b54d41e29ed385ab1a4f22b7504f322294de06c1f888a49e88a6310f45ebc77fe323ab918d57ca9c17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13bb8ef5e8206496d13a7c837edef1d78a9be2949d91f5db7a6ad8686d3c7a35108757b872e81f4bb1b2595dc09722c265f5e4b6e79cfe9532840e8cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88602b19f09d83bb2729b0dddb717be3034a2337238f51ae26cac85e5822c73ffb5376de4b18bb815631fc9320cce238edc4a656d51c68fcb516ca8c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf17ee77004041f4866d927fe3aab256196702f2844d9c7433e2192babf748468fb922606360d16b30526ce7c30627d038837bafa4eec210c1db0a33fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb530a8ed8b454e18443e96f6a92ac8de46a552f97e362232ec0337fb00471ab3bb6b5d7f588b81e58549a2e7154086aa1255b0cd289298fa42bb17bf5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80d77cf46437dd0e53dc9465225d37cf2476314d665d4d05f4770f0a79da832cf50de0f478479c93366bae65091d297a1d4d6e6261cbe527090ecf66e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h173b9c214907d3ae2ad01ff76e008503755422f00f89ec9b1b206a880f5c1349b06b9ea1f035e03efd19aa8415f326947506a82cf286cca32c26b65e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6ac1d43698e25c8821a13f6e45fcba3590e32f9403d4d7c40d320ec2ecac015814c4220771fe4b424e2ac4d461b4a420de4e2680b2004e14acab9960;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc70e5ffc0d297655ac4895d8896ae3cdec30777f611812cc1d72526e0116ec23349f4288c114bbe6ced43501749d36a5eb16af5df4d04e65e596bfdb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e694f7569d2ca368ecf15852daac9a1d3d39db85e75aa6f06ba168f6300419cc85ffa3e10f55bc33f9c767733fcd60daec85c7f40bf2891f171e1872;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b93eeead06d2f17df016cbe25904bed697533c9ae6bb776d043ec6c56cde7c05b1c25e62d995af544422f54fd9ae8bc8ec2042d80aa1644d3b05a9d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14f363f8e502123943a80106da190c3d05240bb42eb03e0efbbb700c6a5148f52477128ff7d95aa5956893b962d1960d767b5ecf99d27312069b896ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h541dc0993d21946304aa139a2da0770f9055d62ae6453fbc0be40fb04dfef8c69fdb1d2af22d13d34b4b2736675b1e8632541cb56c15f386fcba00fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ecb517035fe37f479d61c684018200b9629dcf188b7e8d9640fdd9bbbb7c8c99b638f20ec4c5733f1155ce3c4b0afc27b72b711523153fd9ba1382e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc37578004399f85ae9421c27311e12fbd1cc557a4846e438362334bb1d8abe21af725d46062aad20abdf0199eaeb6b73c2bb4f6550ef324668f009429;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h946f424108fdad0f13732d88f8302a1bc84de50b8fc34260ed6fb776a7f2a78ca668605e83acad3054e99ecfa796268bddd988561e85d03b765713e65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e22b990a2d047916ae7bd055c61da8086611a9aff8cfdeab566425268ab05bed3ba7c949eae08d3c3bd60607afc6e03637f6b0e78b6ac4a934a97659;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he09d21a7814f4a9d6c38438b8fb0e3f208c914909a9ea4c93a25e2078f54167f8e503a04ef243784f96e3b61a544e6cc6e5c55dbeab17e9525888f829;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22858e460415a9eb2155b9cb22fb1a795d82f04259937cefef40a73b4719b4ba2fdb537f4267841014d4c8b1ef9077eb076a2bf90fe6a7e751d2c75e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a3321fe30d5ca8feb6580d1c9645dc14cab40ee6be55ed645414581b582ed207a8b6a53485158f2a2c8df50b1a6fa7df4d3b0ced02c010f2b74d8aee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9432a45fe634496b5ed5c4f64d66db52f7f33032c538aca1af7484e2d60714e5a33c464a328fa6234b4f9936bcf060bfc85983d3dd7d25c63b282e0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9201ff787dfbf5ce704faa2ade1771ec2ae7f63276f8c361e310dc197a7eefd90182aa45f9e4fa0947c45aa59e62bebb9f4cdc668d31c3df9d04edb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he245825b91f50cb5e5581a709b1188d9c54bf2ce3f7002cf7d3be136ab4a3721777da5a5e4a261e26296367f95953436dd8bf18f755cf9af3d5b6cc90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e25aa8445846d0ed2ec5781e6d901355d54fe47fd2b6c37a34cc79ed10bd68486df40a6043bdcc22abaf63a47a41170247cf5c7aa34cc98bd18820a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4e23fb9d439530bf24676c008fcafefdf74a6475e4b4d4ed46b3433b6aa2906f81c3a69cf3da03618b6eedee7686cb65fc88068ca94398347458de0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc747e1a17f92167ec7bf614340ca6f3d467a04d70a166af280bd91f03dc256968bd536b58aedcb836bffae5f1fcf64b55d82d622f7d915f8d10e12c15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc33e54c0d5225fba8c60fe888f33e2a268e970d6c451be5e42763868b3a95beb6f861514f2cce2b27199778411e2ff18d282d8e4886de1fb2f9d7774;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8db3c9a129525ce466fa5fce298e62e74927e0e9ae96d8630ac7cc37a8110676da29ff2164fadb9e6fdb1d7e0ca96fa2dcfe03d5e1bb58af7e831c0cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1f7e0e075c6592119fb4bbb74527e2ecd058a08fd102f1d043bbbfa4a61a7f777424f940f31e124ee9015caf056e0cd41b15a302ca2e621029e5a89d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h755c09989ea1b31de40608d8d620529db25cf8d8e682f4dc7121e7099dec928b300c46f2d53fc3e3c465b3e4c72b6cf05fd756848e8c4ee92e55f4e47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fca2faae0a2643cfcf4f94a2c2299945fa980f41169c42c4847851c633b7ff8643a2525a5ad726de265e7ea8ed9c9eed46c4229c3cc2740b68deb45d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbbc74de90a95f6a5c3141f2a35f5ca2503477d5c3e99c7beca8e406a54d678922f0a13f8c3a44a82e3c79bf8a5e93dfa94e6cb99b18e4bf250e943eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h921d04fe52eca6d4b031bb43807e073f69f491e7478e41a670b6f61e319e41bd11396380f514a9946545be37e6f641f3cddb078206a9ae701b1cb2354;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f8a966c7528d6f169cdc9995ff343cf3d6a7fc0f56231051223a62ddddeed291d7cf26994cbcdfba3ceb0b5818cf3038cba2dfe8234047307a48ed04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaa035d3fc23fda45d555be7924d29eece10d18c8ce52b7acfaa5c96ea6ddb0b8d93ddb16ab40ff7f085eeef23549c486b7afc729f035271d1f363f92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h271fc6d984af64cb82d23cfd07a28e129cc6a75d21963b49e59993190e4865ee7efd34ac7449924d2f1a9fe623e8fe88fd5ad1e859ed1e6bbefe7d68e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha04e9b41a11f064a71a63036c51c179fb5e7d449a738c604d073f596fd15b8c513ad653d7f5fe3c194319e9125526e7b407073593522848799b806964;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb948dc98f277aae5b233f8e53da3daccab4d77e5e96bc37cc0098b451cd18dc821a8219839eb133a0aa50eb26b57d6df26c496e6e0de2220b0a902865;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaf43bd5e0f82578e6bcc8432a797f418df6d9cfe034567fffe3cdba8bd96988c5fc6fe9b06086c36a7a36811c35c730d38e10d1534b43ddc24d9d362;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4196533ccaf8a91941aec71968354332b405b4c7367b106b8070d0ad4dcfd8f6809a00960924d0a02dd3844a737f6f3d1a455fd50906b81fa4b6751c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcff593646e6fe767bdf6e3556e44bbce0cee416119b7499e9e8c80dfa0efeaf11839cb293c13f9871d5883f7e951e7cc2df962b8f8c29f9e1526e9b01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb612fe9dda968d47dc48bc5e63735e047a88cb029382ba86d53dca3042e1738d51710ca6e00591aa8a41a943a8bd71cebe931da048f184bb11a4189ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96c3ef5cf3d8b17b91244172b4340cd97ef85f01e6389bb20bb8f199f3e32b35bf50f87a79178e8da08419910961e582befeb9b2ce9114c4b8a07497e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4e91af4e08a19ba6f46d936b8561ee8b2033404e6e281a4c74524f86ddd25079d4a9e1287c1fd389d362f1814740cc93897e33f1158f3a591dfc3e64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58050997e4c619139753a8b8078277cb2148930e8d2dc4e8708e910d60df46e44e370f99be731b6c65fe06c809717d0974191fd069d7f35972a7d09b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c457b51177d6908988db480ebb3d4a3198dc0c9271d00a6a3bc36baf20ed6ff365b4c4fd3ca77bb36b80345f15b4f850de432dda89f60ff912b0e700;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h183e98640db3d5c075ccebbeacabfd1d795238a21df34f4c1a1b2c715fa9758d75e6347b11a0f952bb1459de3590ca466c55a2ec283b9c4b352c21caa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h245839245aa8a26cf8bd210d4a2f1d943c168e3253e2b212b190a2f408c900623c6c09133427fc486e3f5a4ccec92615e805f77038d97946a7cfe207d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3b2da94dcc01677f2dd9ff2df280462960db4ff2b01050cd79b01f021e15013fbb0e0ecc7f3ab9d47b841ad98a1a948727c3c8913167a27dfe321697;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb2f7943a51341e2d2baae6f417bdfbce2abc0f825ba434ff4d4a528d4a7715068124a267779fd2797d6e372a1beb5492be9764306e3628fe7d1aeaef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9af73f024069bca83bc5f739edc9afed2fb30cbc6f301b28efc4f0d5cbdeb680e8caee475252c2877094e3445e970e07b053439e82c0b2ce993d74bd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fe18cc0883a3b44e9b38f98b7c86c9d91802d5028cf74b7cb0daeff8e6c821d323537a2435ee2c5e303637783a75b83585db594b4d0e410cfb2a1116;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9e35a6020bb68e9bb7aacd10ad60928978446e48b6af5ad3a79308342ab1cfc95f09826c1881fbaa8ec3b3dab4682cd3b32f30c192ae87e98425cff7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f476b0750b9be0801f309bddb2075e28c77654a5e0c1fbd116afa1b5ca2804eca41275a1233b44f552bc15e254610465df16e814e14fabd5d2c3ab4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3406fd7174403c661f22f4451609b2e719940e1b51b5f9bbb49a067c8db3793a4da66241a47a539997dedc06b1834a509bfd81b00914139d4d5e3c8e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fbd1b1440eb93302e8e79b845ecb83225686ac438c66dbe3c40aec06e8327999efd8c300f6742232fbd90153294e2abdc94e36b727b36d967ed86b35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98f21854419438d703dd8b8cdcd1a175e8a0ecccfdb497e6789f8568f4706812d14d9fd7693d37af3e74b975ba40e1c1ed68b79cf8b7c04227360eabe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84f1ecefbe99f9bef32f9f147896597a6c4dbf5844de80d6f95363d37c00fa665e13daa2703012548fd64e79fc63e578091e9814755e0d78f3a811858;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57743d4e2480e666fc6afaf83be40a1ee9a5e5e6f5eaabd28f9f9f2ec0586217da10ba61eaefe26d63fc3fefe0dcb8c301a1f3d0a8c5d5cee4eacd142;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd720b3f84da4aae03bbaf5b48d4b7c2e15b84e8dcc1043e6393acfeca663f56f79b62044a68f811e0b606ad693e9b74c49fc8501ebd626df596138a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec889f4ac88f8afcb6bfd4a456fa4ac1587f32f09fe8a4f199ae6ce32d8e94c84ea2a5af217eeb66c8ab9ed5395b48bb33dfb15e3b026047ebbb9e675;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c7ec4e2e776351cf948b6ac4c840ac8efeed0fe3cfceefb7da1590deb9ef4165aceae3440c0e4d01f14d9e859d4571c815ad289a8054102664d73bbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8452071ef98b177ecd5211883c8c5b4ea84224bc5258ba9027543b9e866e9e2a0df90404e978f63a6224dc6601e57ba91b5dfd48d9b4526caaa611acf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6f7149d78ffe86dcb4b9e4fe2a7ed8cd1adca7a58e26cc3ba9da9df73babadce29b03433c77d7fb8c2c0f8dc3bdc6e5c4593cb2ef6f1aaa826854470;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3232d57aac8eb48645a9e08467a84aa9998300c25c6acd8e104319ee876a5b73c6e7b42152efc675630b849812fb0f2512c42e939f8db5f3da4538854;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4968d5d770c68846e43986ed43318d551452f4fe5a1841f948059d55da13f8d6fbf1e48fb092431641d0c9d9581ba2e8fee2cb5e30b08b9756ccf5842;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb63cdbd5ac608a7e25017ac9e8a8745c5b3972742766e9d2dc0108c32aaa7e2c1aea9aa588b07fd28b5d6b3100fdfd03bd39e7dff7020e0f9a65eedcb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd7d2fa4648258cb3f4287dc62624d081e8268f9f0cb11536d7ed2beefdcd214fd6a17e37d6460f5578c9b83843847949351358f5f30e7aa82a41782c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87ba0afac3216a01539531128452daa5be3bfc7faaa8bdf2032660a06038d0a78e4b9c948959017ce0cab917c76089405098bc58f724c37d1fa83af35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ae73fbc7b7c664b737a40c54fe1a37f11e1db90082d2e881c6d2cb11515b300e35e923e22ad145cbe0ed6a51199a9184234913349f698cf234d7137b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37efdf2f425872974398d6f234f5c3de20c15a889159e375428b6a3f65d22ee856a3a349e23d1a4a050fb1d6fc2937889696941d1cd46ea2c6cca22d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab50e85bc04be413530b0d36a8affbdbcb08c381786aefd62f9c361a41eb64af462e714ebc7014df38c53127e951fc299cc99e71b5aa7a729dd95e578;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h813e067213072b382cdf92179b0a252c1a05dfb8c6404032c01da48c3084badff46d6a2fd63588636f6cde13746118f6ac7f4606309145d6a996c9ba4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d5b23d28a833432f4212fb1d5cd8612d0bdfec3b2b1adad4f32c2e063fe02473190b590a62ecf813e401f97b02c5bc64616b82def14b0a7c92c31567;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71b0486bd18c4b9c8ac65609d522851177601ec98e09c132461cd6903a3ccea78ae0aff6e9dea4fa54cd9662d8ecfb0f733e0ba7eba89e4e8c8bfdbb5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he83d66e55dcbe086a9bbbc140b41a7db7fe8d10de0858fb0a4a5d4efe29ecc8e691885eda0144b9270bc9f6fd590e30117f8ef0ac66a5ad3069a7851c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha566a8114564a1607a70038c576dca631da6d95e98c2cd82e5356cd4003d61e24ced56e964fdc4f1b993c548f66454c3ec9e13d48c553215e5848fcd7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h285542e17c5b3cca628a3c55bd1bf22493c8fcd49184ec686e59126d8a59ee28bb0ce84dbcd7d81e41012b2f045c40cc173d299dd9aa95566e373c76e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93e0e29b60aacd044a83e757d345df5f35cc110686cb2d9a1d83baf344bc3393b5e87d7f606145e96d174e2b4c3f3bf032f62eb6c76b33c8f23d0ef89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h831df8283a5909e2405317e9ab0d1c6ac234a9c04c9c0ff76c9389e2b26c78b31ca7e54ce5bf1a9f0bffd929c1a400c377a6015008053d32e938583ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h195037c3e77aa8a6a04677ab5aee216180a225dc9caac7f3c6e273b56dfb1cfa7501e000c834f65fff9d81dc15c998bc861b71bf83d3dad24d691495;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62d9e0edb5995308d823ea3232cb7b82490a2b0bfe800d3b8b351b56773d2df1d150d9344742f4788fcc5db4ff19abeeb03a63cbc9cdd5ee9b3fc0243;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8639ad83efcc1277b53dd9cabb0d18cbbceb79183ddd16f76c9d6e9460e335e075449eda8c3aae5f8c0c9fa30ddc601c736fb0ac80a44652532f42e42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he09747c0f0a1f917b5cda6829d37451b9085b95ccc80c4527604e5852c24e0467e8b3f2b061f1aaf78e776f5db969abe1ee7c4807b4ac0c6053dba012;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d2ea5b1928ea5fc2cb1d69fdf3cf44305043f0d047e5504ba6671b33f2f87915e287be6dac176c66447bd57350caa178a17512952c00bef44ad7aa5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82a8706a4fbd2f876872545c79d788f3ffdc5e9ad79e6a09d78479989b0d942d08f06b09cfa5d0acdba10b87c57fde1fc27af3bc620f8528f10e46d3e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he09e4fe87845ed309af0dd9366b0dbbd8322978ee930dd7d89d563b7cc78fc8018661e976f825b2641ebf0b911d2e61a92eb9a4543f9fa141f7d9acc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6193c232c26295f523b638e02ed3499e06addf220ca107b02f1b018aee69f52f8e35c5df68017b67d451c284b62153aeb64cd66057c73beb8404b79eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha03779cd0c48c8473bfafdabb4d5748a1a956e9f1dd9b95749f36ffb603c38cb5831a398114b41fad35b987cf66ff10efe6519281279ec445321742e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c6655288079d616cde13727a753d768843175c34da6b46f493a0d553af133f1937c1e36085320f5a2122761688cc508f5eddb091d85b236d0f3977f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h403f37510f15c34302a49e1e16296a2f220ba0575c1411bccc5af814cb62013f30084856f6369bd4e87ce3556cbcfa192390f03a7b8d08d05979f8194;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ace551a367ba16d74dbfd7c45bba6ebff49b1f004472e7eaba3cc26df111cd95a6573109ac0a064a8d5293b2f1e62ed7b7c7258a2a9d6d1325ff2364;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bf8502bde4173abca007099a37386d455144b86d1e512c962c2c70a2e0587ac5951fc77f6a4bb6a306ce1fd1fcf78896d7a311df56d636e789a28b23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2927a2aa35bf7b8801dc99a8b03d553c25936cbb71a30249c1636b06eca047d82275ade732e5bb530cd5a9ccb7b545422d719bb4c8816684cabc5b560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7788fdf445f77449e79692be70771a019a476b52b8f146f02d24526f3a39e52e1aca2580906317deb74050a7e95c2dd22bc0d023955c66587a0926be0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ed9d88642f72247ac43ce63db17e17f1049bd838865833e2d4cc4e71793f7d7d9dd902170d5d2da09151fe5008bad8b68f64633a507ffd19c1c67413;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f5ffe43ffca27029db956820a5c6a08636dbcc243830d67db3994210e10065ac5ce590b585555e6a97bc22542817dd2a52a8067e67aded3924635ca3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h955a9af7e276ce17c3072c8f1ff0928b954decec1d50da2b5a87ab71248e7cd4fae264f1361e86bf86c454f5c91650902d41b23c83431ddad981d38b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ece276e70578f1164526181fc9c10b4a2b4d1572bda2f53232b27f5555731b2427c8119675a08e789eb48d5fbf6a7809751ec96bfec93984e389277d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb57e1dc481068b5b6105e0f24c44862d429c60c37c5b526559381143bae7eeffbc62ff0e21e488cff220e1982621dd2b9f85a85d963ea538bb41fbc15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcec3d1ee1d31352619122b4d0eff3868c52ffbd506a582e6e0b207b4f1af054945f6c997462206b3cdc608d22b8df5bfd1e4d530fe4aa2e668df24b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a550d20e727b6dbcde73d8374ca73cba66f1f2390dfdd527219553d933e495642d2ffef5ad42884530544ca8abe239ead92daabef4d4b1fb5a9197f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb12f64b5060a9231641c84811b8b7e72ca6c44f7d0513135fae9733290e6d22bc8bba9148b4f667acaa53a12ada139d023e6d4647962699d6b9e84063;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f49fdb1188b270af0fd4e47b82e0c873d410df31344d78d1b83ab282c1197b59aa1691b2977a0a0fb42cf833d91f0bd05f11eb50cc017eb84e4e49c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a1734ae62a1910de90f2faf1120c67180765a628b74df941acf036fd034af6a38353e86fd13690e394c870aca1978b93b92ce29770a30d4124781f6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb19375d8d925d18188f9d32938bb238e68694dfb9cdc858d10e398f63a13bd72f5436dd02445b78eb2ff50e2c2c72bf469a30ea44d243df24ebb75ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d83e9127e73ce04cddfa0d6e0aed29bfb5da3f0828cfcf5cbfbb2d7272af3195f6569a40c7889a53776ab53475b0fd1f2707a5d98c8ce43d28fa7d50;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7289d59bdc9a585b2b0c322292bf9ba27cf818439bc2ac5bb2e0aad4ba051b9b8be6dc6f7c551ea545a9e275198f574c42cdc3a8d8837732017b84a0a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8949173252db8fbff83c7ad1648d183041734395c26dcd98fe003fab2d9b35d328d48fe253db29346a62299bcdd9e11bdf251a24b387598b42a07e6ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c8fffb776c510a8297a3679bbed152b549cbb5cfb1806a4bae1482d29480f2bfd2c3fe445f286eec4af26a54c12af213463983e7456415f1522f5871;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf97c300ca720c216bf26e730c40c68ce1465b8eaf598f58c211dbbdb19408cf34ac8b95eaef9fd0dca70fdaf3756b6e15b603991f8f6506a6c2919bf8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he09bab42ed3502f0f9caf5cf0ffeda1e2e735ded0319f1f7c152b593ff80a06a7f544cfde39e59e2cdf7f9e97a47b6c3c054c6815e6f74a46d7c15f72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc8a41924a3c984358d3e47963dc38d2c948e71a423bda5ef317a37e9752a5ff4c11866f345a530ebab925b030cfdb6f2ac530190ac803ebfc4008b06;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a4156461ffd7a275452199eda0e730f67945b066e08cb0d2e6cb415708d53bd6f56d802f78c50ec99b4eb2d8ab4c01a509490f0507d955da17ad2036;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dec239226ea0c0797aff5f14fd68be8a29823ad27040893a20e7124a50a248ff1fbea80fd220efc28cfef8a9d82b95ec887289f9fa637448e5f855fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bbadeed2147bf4bd25a002388e85f0490545bc607440b2dbeb1140650fd891155bf42b62e0db93def5cb36b43042237e2471c4aae56b83e347a8bd91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffb2186b256a7bf57be6d1423d72b32e27ccfea987afc1179b66c378fea644df70bae7289255158b94df84e976a04cd1da9acc9541c45d446f0c7e26c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd526c8369abc6b74ea1d68776ec7d4e9466dc5876bbc5d62845662a8e0ff9a7dca78958327931b3842f7e857111d70ebb0a2be89b4e3088cc012029e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h258a55adaff74adea09366df3bb3d1a304e7e4ebc04f72d7f8dc401ad1dc4882b6e777ac6de6ee4fca9fd15e8c3a215080b5b9ce5d9c7f22b808339f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85eecea2234e9702af542291c2d83e97ed45ca99d2354936ad715e8a97a1ca2f83c60adf48e79ed27d8bf95a9da457a5440b32f984760af4e14b872f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde168394f1f5c1e48d932863eb50c8825b288763515dd1e15e475c8327b13058ce0de925fc8b7dbde967f5b859378b009d3f479552a134193327933b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9de54cf9317e018951e60d24b59e9734e0cf1be6a2bc0c65fc0395ec2dd429507848abc67803d661ad47bfdcf8686c051d3719d55dac5ad63c2fb447e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc69f7aa6b91ef123e95b314941167dcfd991cb1aa524bf4fc8dd5a5f43fa330acf5ea814155e5a62e1dc0b1f6a129cedf87c56046723dd565e978de9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha65a1c6369511b17c2cf6bb5609879f8e9056bb691b6418f1e03f500f70aa41a7bf5c9ce9e8efa5b17c87219c325a75f6ca3e66b75561af4d7d002b97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f39cbc51e49ed634df39e09c30916645565587f4edf917c4ba51969ef0a3c725159dc5aa7f1dc2a80d711835ad8af956dd738dbb3987ce68e796f3b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3b70850df84ede07b90903160e4364f9a6b7ece2ce623c15ebc3366aa398dff8df99da276551e9ec4e8484dc40a59cff2889f30b16f63e3f5ed1367f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf687f417d4fce349a61eb15221644fbd5cc9491dbf4cb4e4d0688dccd14b9fafefc898f5229c76de7ea7dd4d5d2806ecde3a9a908c36f0cd7f07be72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac5034c06a8ca6843012dba13318c70a2f498a434ef142ffab7ec91e646576eff1fc6ece907ce359eb03cb63599566cee01ff8f61a92ac1c089362aa9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc78b5a49350ec0a1edb25b21a97aa8168504724c60492e88762dfd9621bbc541a230ae0b12bc02198939cc6afc7331fd579dce78ed98694f0fc40ba2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e6f08516c734383fb9950f816db33d1013bfad31f175eacff522a5c1a506c0fbed93f49bdd0893f8709527ad09b7a7902aff94f9b7db08debfd61c3e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29c34f5045009de7fdd092460518a112980098bf39096da81655e3eb87188e4f695e7e53edffa95f2346352e20a7ee38a4e77a1bdc665e7dad4bfd3c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33717e75c5f5230c433e012e80837f72882170126b66af373ebcf47f695de6adabc514fed0f2acf4a0768b923b45e630625ddf161bd125f870b0e2d49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39bbb66036f3c32253f05bb037fd05b4b65b4850517547f86425ec9422a11b266e67469d51fe4e0e7c94cbeb99318e37283cd943684d1fbcb6c0157e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h344b963076c864382101c9db10981e0d0dfe0742c2dd29184003e05a4ba48b8f0757066473384ebf9fffdd9b7acf86c86de112127538abc5fb7d1b48d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf04142825b43f5c2cb02ef72f2dec5b30869af291b5e7295d7dbddfce5b4cbb6ae5725c07135929a8985077c0416ad21b81966c0be9abb6a5960cacef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ba80e08a7db4d56d767f958b7c68aaecb95ac3de9852b159270cd3b25f07536e15ffd18d02ad6b600f42d312bb56757f09924e1216cbc4ebd2c13626;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h370c5864216bf5cbe18a11bc4ff06bb2709e185803d0a6e81092e50e6bab0994900b36e5d431b1e43179223d335e940259a0678e8ac8977fab042ff51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb886300812deb89d4bf12c91b9bd92736f1b39e853bbbc4df09a3bb639a43deb62430a137cf8a1c9e6d5386223104dbb105bf51ed7af97569249751b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6a75f9f7cb36d24e53b114b27ca9cabfae92b8cdcdbf3240782c0df1bfbf53b1ff7daf668d6c2d239002f4d6b98fe5f02713c1ccc5c5485e7446878a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0c0fec75e8bc9cbbb58868b1c52f4bd2326f180accef79087d2e772d16ccaac804c914b976c26d12ea81f6ae47ce36463ed5022b16cad56dfb98d591;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89009f4a78ecab6d6987cb1a82ad7afd6412126c910bb36405346c8ee47c5e231c2bd22a36ab1a6b4c56ee42be2650eb04d4ade3594eecdb769fedcd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h835375a0187f3d5a22f02e35fef88d362b31c6da52c1c067982a75d92a940e42bd3d17ed07a49b10ce05fcd84f4356f542a14b9424aea87ff370f35ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f09143c9fc56c5f147910f1f48941552db6e21e739e8e659bd6a9c0e38d3b3c0e5f27ff8c8796ab949ccf76eee95667a73892b7eb5775b20f7bc37e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7d718109e1873e269abb30f30373e7f5032b3f11de14d063e58aa1eb6942037a5fa8140fc7bf46ba2b4f92e06b305fc9c22de2fe48baa62502d84756;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h299911968f1fbcce54ec60c3d561c8084d5ad62cba5d0c4cbabaa20c0ba8db01c1576b4761bb65614821a72fcb37d5aaf293e8b9dd1508b40cd1f2650;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d01f86cf1c24453165a99b52b3c34b5bb3d1cd54a493312352e850bc76e697bab2a90d0f956b6612b83ee5444c3b54b2c9ce73204d1105644b36804c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he46819a1095796bd17be28f6a745ab77de4cccdc0d49a98d36a5c85469d0754ca43c8c61bd8f7c514241969a2990b12b2200a00cfc14e8c3c1ba772fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea80a7abbff17a5795d12acaea57291e576e6a34bd051d7e77ee5ceda659fc43521ead1c39084240f5742201a567464a9a4992256d8691260bc71af8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h665fb90761fa631ddbadba7000faa2dec1dc03398f52538e578c4fbc41bcbe02d2635aca0f1a1daa8cc6b7a98c93b422a3ba0c4792f2d7afb50f65b0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5ffab2aa6ce61e8804f5fba318a582c54f29f189f815e0a0c8f7b7fe15113370edc19940a670ca6559cc810ee137eb796fabc9bf098a868e612c0155;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd06cb323642124c91ed000416b7233eb2ecbe49a23324e7698ea1f8266e703ab92c047f6c0f579d1b55f4dd843e5ebe93e89acd9d5e45703af48c9a60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7a7714d295484292871e1686efc65124a493ecdc18d6c8fd170fbb4cb17d9071f61e0bcb86d2ffd6c0ef7914b5c1b74366c28bb36b9758af6ea03f2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h733a64669cbd241d806963cb457b592d052298fe5e6e3d5f27ae48e91bfb13e811c2746a28f1c45b5747dec2545674abd37fc8035669d104a25018edf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ca9fc5cb292a857f8518e08196ca213dc8cf5db63305a7ebadbe18e04b74a375e86a0efb6897ed750f1144ec72545b7506371f2a5ad08560d3700751;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h353e62669e2ace46c45c88b028030052fc114edb5cc81bca54bc1836c1b311f0024acc8751c44d1283bbc21b776e27b91711650f8a2a19dbc33718366;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16f7683d9743d4b324afd31d7fec213c8f4bdb2b0c1e8fbebb32ad22513daec19d70f8675fd4d4390d6f4015d49075e90a626de78cb7380fcf48ca2fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39b7eb13568ddfe8cc8d5909ea39b29d5a70f7ac7c92476aa4b343c588cadb9ebf94400cf8eae408eb9994c8c56a44149774270d40f4a2746ca0017ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b950b796298aad40eec277b783e8e37dcb1ff25e6322fd24637180a0cbf755f96a4f0b1badc0b4261e53efb0c2448e65416268ed692140dc35f244c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h846550ba65d48c16d953f830eb58e0770efd8dd3253c5c33636fbe098d43cc28b407461e2c7554d3de5c6b8592ba0b0efb4d95cd69943301c7ca58a96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa688845fe1d3f098401b4c37b010462bfa8b046f7beacc6733d273f49d3b84e03fd2cc59642b920b6e6120a863bbb2d298ba5f8c329c0239351787a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3e7e26a3c36e0bed0a773bff9fcf6d2c1e24142edf6076845c41be628bb4f9ca3537e5d08136c8c9eb7654c8ac43faab7f25b5961b318fdd9f6559f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb82b9af5371d200742d991841df1a1594936f7185665fd4567866918b9f1d6880447075a7d12ba7214897e7ca25b20c60f3f64ab053e55011ce485f43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a46a130e945996b86143a8adbc9cd3c7ec175c8664f3c5a7d3f640158a2148a0946b875da2f9d1efd408d953e3ffe978a5054e67d8dcdcdceda6159c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c03d458c04a2f9b70cceb2677fe93a16bf15df9fb95c390ad34c419d0739ced12c3b9b09793374bfd362f00dfe4d702ff8ff3ec932cbf1bb3183bee5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3304b524b0d85501886012e1497385f979b94a46e4674a8706231a7716ac4e17d6c51d27ba7932cb5bba168b098b8e3a0f002c71d67c46a03745b7a8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4edf5b99a3fa17734d0d64019c0f22cbe84be22b38b579f793a8494e39a4a004efe5b57a34519ca3624e39b4ddc2dcc70d766c13b037f7e45ba16594;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he40a474a9749fb43f03665c29e63861bb95ba1546b86b785d9445b591fbd86636ba8b2340e34f2788717b86b4c54760a76820fe3d68af71b78af556d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h753234a0f478bd83e8753b4b6bfe22c70b98376db4528956bdb09ced69a92ce38a5acab7e9a191cc08c3b438b215c66f4e4e3c96693f1665afe969f39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdbe5e1ab3d4c83c126b27722483c348b6007db08a25a6506bbb79561f6182aea16a3fb07ff9ebd676fa9c83aab9f24e379a3b9a648e9b1a8fcd91391;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7187823355bb3956b456a217707ca510317339a16e497224850dd708dd3ce1ccb7e8241c077f335a91e58bdef8c34299feb91460207d0611303454fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0a77548a666e77aaba5fc20bfb8a8276cc7ef1feb76fa42983b485e996aa9c3338a51ccad05bc7b8af3cde33de94512a68f228d9f603387bf92e3131;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1996412d3c40ed711482f84cdf1c07a83152b09037264d76cf3e4d6b960e13cf4d59129d9b80a72a0f25ec8a98b0d699ddf8e2ee47483849e96e5045a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a41a1d80bab9efa7691042c6765e4f32e67089fb368d39ef1e90c9bb459c2d5adf381e230b5af3648ead74c5f949069a8dee2cee97830056c063bd47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h700a199f12f34366ab6da261215a8dcaf75bdb567f513eb9d1725f276f480be79ff51544874da9f6bcdaf63f7fef1418ea0fe58a7011929030893fcb2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0c43c2df518937df284334946fc57b8fd6413c30459a7314bf34b22fd2ffd59f60bab35382655326e28470a2216c7dd788f9303286e654b61d23743b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a9d0889f6698a9d220a2764ec910ab83475e74bf3e6a4e6cb59c147a55afc92789f8f3dce72f38d015b6cd2452191218eb84c77b44b500d9b93df00b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8bddc7e042435670d6e417d48a2be2884a854fb522c800848f98fd78bb55a66d5557d303f3cca72b8ebb1ce009cd83f75b6b11760ab57ec1a80fe81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7da863e880acb6a0720fb8be303e81bbb8fa4e2cc67f8742fd3b98c82abcb08550303d7c2cb25d1e2fb23a5c44bfb8103c9ead59355afcf165e113f26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1214c4cd48ab02855960f73d77b48bd50e1c8afce01bcb8d96e1eed5db50e0fbdd916258c9fadc65f2e3ab817de07c913dcc67f207f0ff8f31bc7ac9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fdd35401c504b89fc996c6e6f05e1d0f176b1bb618163ce1e2b1a28366a92e106998ea307da988cf1a5a2e1538dafd9fa42d6bad48022aae3a93b9c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ae372364d3c54ec0ea220751013f98db1c819f598c76311901f725d6082a850212cb87697b3c33f9068f1c55f5855f579ee7197664d15accc9898d7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h688316ebafa6c175cdd23ee2563c7e2fb39bad43831a6ea33c81ad6d492ed64b1a9ba597e2d5a05fe348df453b14da2059dbbe6c96918118a55d10cfb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc24ef71a0ec1ea67e4ed5cca975e2cea8834d69e6d1e76449c71cfc8a5ecf19375efe0b94683fbac234833f665862bc65debc7b4375875bee308c06b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b672e378d78d73b46ef177ceb13e84b7b9b6cae4f947bf4a4bd8d7e946feafbcd0a997c58d22da90ff142ef69db1f728746978261f591d608fcc6552;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6ff4e15a4ee46edbdb1fc766782f3761c9e3a844d60b1721c188dbf4e8e5f00437846322b74030a90c784f4b42178ca927f48071659022b82cb54525;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7689f4fa8639097e4e5a1540c678643477259375dde89a1258d14c5d8c6abfd51b3056693ef36941a5265ed4518d599bb420c2b6eb88f9b8844a7c09f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28b4ce9e943742af678eaf80af9c0238b7f2e1a98d30a321ed904cdd1cac5defac1e6a09dab76a54d7df5a81fd331e7f0290e2c217de6717701d5083d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bcdad65e298cabfac118e801c4d3c7f8d92436728f7dd6b2520b3ffa4c78801658029e027fa14eff211cb75eec6cc0d7c33ef1f512e037feb0eb97b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7cbc948dc859f94993ed54547d6f41e9d222e369c8c48b151954d44d378600cac61ec7dfaa4c7bc5b4b603acc9123e9abda4263b65bcc1db0b999a18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63944a790dbf7032c5ba1db0e1c7fdbd3b8d8eb27e24bbe47d884f750d847e72cd8f57dba36e4b07a430dea97edf0e032d573afe7067698503881f9da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d72cf23995130507451b749fb37e3295406ae9cc76a5fba9a914d87c72e7c5da80952178fb2f9f02867c1751468cbbd8805955cacc47cf7a463cf8ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aa63f0d17b18704321f993c41ec8326d8e391c7a7a639db4e6312e9bbd5c68a65f39e467273d769ad048c10158ae696843097d11cc8c9b044b548f94;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h829c1a9aa4d244af90b6639ce63d0fd2919c20cb94533f5d5a8ed787723c2dfabec0cdc343022378e551de8d98325280f5cff1bf08d1c3a5cc5ad262c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91a9e46759ec913ff0e9320978a4ac463bf68fe23fa80267a52962e1104829c3c30648e3f002f3be28bb77333deef16c9d662c3de0bcab239fe38f05b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9598115da2104616176d5d988da5a15ec2bdaea1f5e6e3eafc26249b81862757a412d9819afc7e41b4b4ccb61109d8b746561879074a2d051d57b776;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3ed94747e295134966a52f1ed1685a4778ae46525322de32e47c3b71267f267756b6cb36adabb184a43d2294e06770a6af49944652f499fa4f437de4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6080cdf1574da65c1f2d62717c51a607bea65a74b093e3e51a557a7ad3762c2d33426dd7af4e0a7fa06cd1f9ae91b79bb79d9b2fd09b153767a190d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ff75819678bc3b3318a2afd090eb41971a2fd2a48d4b44e1209a581ca016feef8ff6e2725fb2fe414dbe777d90ed22c5d895e32bf8e6080c0041e3a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h809ca04d1e0e02b98a4b1131a615e4ea7bf25c091d15d1b6521f715804128f5267f352d54b078eacce9e1de432ef9cf30081692777cde2638a263d8a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66df98caf1c9a364bccc3f032c04da80f399b5fb14153687a1951e38f140b847b189a18844a92bae9954bc7b60546a91fbd88b0bde702216f28b98d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h308ee50e92cb521ae51ddcddca68aaaff81295970e570bbf712ffa614f23e1b32c5578408542911c9c5101261b9c4db502b0731ad3231eec966e10e8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc98273ffeb74f513618b1194ea4fd812bf3c381ff59c442885b7794c75e03c2114df238f84f0bff28445216f6f167df1bfb240244dd088ddea954993b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82b0bda73ff3f2921101b14be6aeab6e7ba39b1265968e0c2fea4ac266bee18e438ba61f858cd79efea465e0467f1b7dc30ff575de6a1e436aeb29626;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79467121a3dd9dcd408778dc4b246bb095c66c574eb0349b9a38cd5a07e6b87a1d5d608064500d35cfe7c48c59fac3c2ea611d193a0e9d5825fcc372e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc450a53c0083fec6fc87b3422873dc4a1c77779123091bc161199da724e5f794eb830c572e88355d728c355e01e8385a1039546806a915f1f8e97009;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h182e05fc9ec4d9ca515d68bb3095a1b3681e631f9458dae309964e44d8ad845be7570f37156793ba52b3c6a6d89d865d4a42b2f43079ff247376d66db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb992c9f428778289a493bceb28bf1c66de72e28ec296ce457081a858e771a9ff6a03f829c2943dbd4c7fc34e2f24828441078f04d108c5f71a1a74470;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a30766d267da2df1181bf12cc491765853dfedadbcce1cec18906c694c6c745037e3aae2b931c9aa4c2d99bcb2db22b9a8047407ceec397f2a802182;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12e3c53db5262eba4d9df00280a949b38aea5e502545f1bd4dd49e0dc0c75cc0267b56c7d13aa93d124055cdba7a2cb7cfea3eaa6e1086d930dee54cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2f72967cadd220b8ea38444e42341493536eadaed572dc98ca43382a661e3c167a1724593866a731f3e224d15a0abf68c45110a5f0c6be9ab5208f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fd8595fce23a823253c7725a26206ac5a498c82e06eeeb2e08eacfc582b58945eee642a100f970ff0dbe97903bae6a3f6fab5b9d6c8610e6cdbad199;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4e44b64634929fef9a75f4e95a1f61e874bf3fcb121158f7a723a26096cb28ea0108877c336cf4d44d6ffcef57f2d0d47e67470f7a3dbdc7eeb6b898;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9123b12de604181b5e8d92107b5c1b6e410fa2121523787391a822a6cdaf0287032b728b2a9346da7bcdd05c17a4d0ec1b3ee8c601b75cd3f591988c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h657d2572a9eef60a77c2d2c0d69369a604a6870627badb9db5292535daabd42e6f45d6ddaa6f4069547bb916c7d61927fcedabcb46e3dcf8aa397bde3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc07c36accf0a66eae0ee8dc6e268308837b53274e767b700e9356033d1c5f10d692c6901914433e4beb2f98e6aa545c05541fcf20cd4ccee9f3bc9c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85d3c4ca4e369e5e1b9046f533063344fe932deca82c05d8355487190daa737b6f3f414df81f0e62924d19dc1945131bffee997f327f2bd6d6892e983;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h784af08b6f247a236dfab5bf59532b3d3012040d9cb50b8d44c924495e678963d3066af674c7ab55fd0685c3809e24f35c6064c0c1fd7ea795e0f87a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h166d1b6a380db224a03f7ea6ccdbe8828e601f52c1b2ac1e28b2399dbdb9ca1f9e4a6f9988833fd99faf15529c7058cc447f5cfa6762852b5ab91010f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3394a81b0b57f4164ddae750adbeca0313b297fedad75c777cc2cd04f0923c730647456a9d043139fb36dde0d5fdfbd9859b1099690f751d5bb921bd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde926d1efccad357db069767c01bc3d7005a43727be50a1390f48b2c50e42c3ff52c9cf772377f096a02302250e8e0437a41eb393e03b51a512cfe50d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf7c0fb5bfa997ecfe99a22a3de966e83f3a092bea8619394cab82deaae209efd726a6e017cc0218907e639639322991b14bbacc567f027bee22bf3e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf500d606b49946f8035bba23b3f439901facf958a644834a00aee837dc21476a9e33c34d75bc3830ccb23424603c620a6eaa67f8d418e47a92a53c988;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a52376a0b8231b4addd1ebb9e85f3134de0fee0c2aaa94494088a867969a9311de644703f393a8e76bfabd36ed6ab22b2b8cb408c597c208687836a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd853a4038f746a04058b0a55b7451aba98f982f4946ff9e4cc544216e443304b16d441a7ac64bcc60877bcfc567c99a60214a4ad4dd872707027b0dff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6207586812139eee185f5f1d095ded55e2a8b346efdc63ca7be085919b6751948c125a69560c9d7d44b6058a78d3f7ff7aeb7bf2738349099abacdd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d26892bf3ee855a7425169e7f78c255a24bbca8007e5a9884c8367dc8be1f82e53ee0f3389f9773ab9d50fde8df0c50f8efc07fd23bd475f249fd319;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e6f7e80875ec8ec25e931a7feda43ea41c2cc84f742bb561cbecb0d01ad11a2e898303ef1ddc1dcbd490f450d61adb8790d9eae851e31cddf5476aea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f8ee2d686e1943fd564803778b51c2f15173b941cd074dce16a5977786830518ef8674ffe9ce777247d3f8e5c09eb6e6f351de04806aa4b0fdf40a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0ad192a6efd20bce33d481adbadd3779d17a498863ea6128ea22e7e5f36b4c5c337301ac60a22b1860980f26277aff7c5d453bcfbb731d287743d63f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c0d5d760e3406f84451399a8c4b1cf552787c3ad527a2e8de9d501c79911565f204f2c6149da7e8dcaab66a924ab6d3e983fea4fa2f308986cf9d9ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fb1bd146ead7fccf7f8e5905b511984706aca7fd3cd397928fec54800e3ec121e96753555ae6e89cd56d225d318a7f9bdb73d26370cc68f2cc1c3c99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd06261bfe32d6f57744d62232a2846108a1d51995e10f04d3f63f3438abc504aa2a34c1dbfc38725833812c0d1a3319ead3c8f1e6b2fc33a2e23b768c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h584c37a4bde269eea70339d459fa38f6736dedf38252d6146173695f01ad20793a406429b1b2a7ce8374a9807cf4e372ddaca629372c4402e140a3af9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h743db50722673755c808fd3f37db3ca688df45581512855627a2a6edaaf94195d405a0663f7734eb711669a587ed1b43bf4b4875325287a7f88fb532f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc0e4f94cd82430b2d8f32994f8a7071493ba19b519337b2948cb4dbf99e3a22e3336f7cf1b5e79804c79a068b8446d6ceabd7af3e944ef60c1f1fdc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e646722ee113127acda573467635a4a3f4d5af617ce056b5a86e6d53a080610dde554f9d77b577af207eefc1c04546cb26254c181f3157eb6e309a1a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf271f383157a16c8849e582ff082f4b951853fe0442d05be78c3c01fa0ef1c18338d58e05a3315577d9d685b217c14acda337037e0df29a4cdd8c6232;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcc469fc5ccbf9429b3ff37b9c04f3f89131974c9ef103871d897d63971ca6e849d3abb1b598b53d92e6babbdf8e29646ee4112a34c0e348bbd025e58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c300aae0f1c1254a5128ec8ef9491955858bee2bdcf68127a15222a1060c2d3d41337676ecf995184bc897d5d9bca5d0149b768c0114bb45b5d787af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a49bbd8fb891b44e35a2c752be57d9b01b55125873d79cdaa0ee42aae6fe3a3be5c91ebc2f4bd27401c819d7883a873c492e67b05222f65205223859;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3002079176d0080c7c5e64be97c60d2cb58caa096bbaaab7b145f72bc83345b031911de56b2d6608a19b935ea8960f8452de25f419488cc284a0d29b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62c23d8d093a44e463e3bd80dad4defb0c01d79f000c11ce26a5027e92cbfa865b219defee4c33fecc9ee58e29671e8dbe2a25573c0530325bc56af2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb3992951459592e207e831a2df3aa028f8e40a35331660255be201203ab93633f7fe8c3172ebb4225d02d16d71633c667b42d73943db090e06c172d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5e0848622660267c38018f72f8c7e3e2309bf6010896fa5b9339db8d7ca1c18d444908b4106133664c54b5ad0be9744f45d4f7a01a5ddfd449e66df8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h401b159b8249303169bd4181dea3952cf72a02e1a63d13b5c633712ea842d9d90e34daa26f6a4ad4e404e0ae554527a78f78cb86794a3517da22b8537;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6a9322dbbf5132a4528514999a28cdc8c4813a663442bc6ea062afbe247ca1d3c0998a5982f1234f6c95bff44a3ab162eb90fbab87fad0ec41771469;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde31d9580f91faad8fb8845bf9e3ae70fed7d4045372a2d2245efa4ed30a6551c687be8a88ae29d8e1b7a00cb907d2aa3292d8b53555943ce0c51ceff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f20820c7212c6c1593b27416cfde5e02ec056b232f7bcffb95ac1038f04e4c637bb3c45a7406b9fd23641f14d757317e74e30ddda1990daa5b765a9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c2cda5eb6a19c40286ef65439e064abb5abeb7456f6bfec46c5544f0e057de099d1a62bbaf3bb667eccc4c851c3ebec8e7ef1961acb4c6b4d9fe78f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habc6f48a629755a70576f47438e14c88651a536a252a3b8b1db8b71ca90da177986881e49457d97f57113771d9bd3ec8a41313e25f2c9993327e0035b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc815ebaab01cb005b0ba5f1bae025681d9c3f96a6ab4b66f81cb415dc77cd690f6e023e8e76e0a8ef2a800910c86f0b9881550665c02748f6dbf42c70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71153feee6dff9c15d4ad0d8604e37458a8ec332c2398b3ced22c1aacb53a8ab35c1cc5f5b6e8b13b5c2351787cc4d6df04d7a7f362db7b86b98b8dfa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac7027f2dc51855e5df150935b2db62e38935f7e43a3ac82986fc5bf1b2254dacfe3185bbbc15f986315f042438afe6be310b833339102d393668f09d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf56dea30f9313048cd66362e53a20e64d26043c29e8f451965075d630b82d8025017635e2d243da763cc5feaa0ab1c8dd90b5ee801db03fc50ad23521;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha46e32a15ff4d40fd3ec303292ed9db8d592b4fb15d52582c037f2aaf6ccbad306fcd7c1cd0c0e465f9818820c7ee36f38db74e8632727fd741bf83cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfab194a0b89f7675009e55eb8cf9d19f7a2814e490b3d2f7cc56648b2b6bae9bf2804cf5d7b577cd0e1634713b5e73c05017c5d0d680cb855a8c56637;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a8339dbdd7717f08d072d5d3d58f2ed5383c7d1edf58015e8b3ec1e3b52be0fe3d9088cce109aa2fa7defc9ec7123d08f362c36df2eb4f6a8f57a9cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb30537427e7d5214f80af2d0cafe22a09814d62f4ad703f449e9c0a4481fea941f488f137e22d1e98f9db6c67f762a20d052248a32b85610c982a76bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9b2645c2cc0c199fc8ec96e2b23fd5cac7a83e8caaf2741f7a08745839c3df0f84c3f8f47ad87e99db10ebff7515623347b0f695298b057bedd39c27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa9a0e2832956d9505ffe4d8cd87833714d78798fc705bac69178e9a4b6ef4bc3df50da145e24707dbaf7db413a922442e285e8e254a0223bb1ab4845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h674cd93ca28154e783077ae4bbdab2106514f323f609071099fac57e127d3fc72eb4c0cfe00b49c2109e3d29e8001f831d1914b55b96427b5db522763;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8be8b12a9ff60754bea801d40024b7d66423735d6cc088a2da9df0813ac253261ff65fa15dedc20714378963b115d1dc62705fa4838c7aa6a88ddef6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd68adaced3942dc2bb5dd417d6438cde4dc84f68147fb1e4fb4221815d2890e5ddc96be1b8a76440eaf3aef24525a81c1a7fad2ab70f035e14ee6442d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha44b561a68563340fa3e4875aaef89a64c1430347b32e340d0f0e9126c525ec3976beb1217aea674bea6f42003614226c5f6cadb127530d068caa20d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73c9ed5df974bdd7b8fbe14a49b9af329e468d140b1049a5ee6cff932d4aa14d5129295ce6c38dfade304e86eba071fb391b483a4421b9e3ec39e727e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41f7e2fc9d2d565733bcbd658065227eb97d1fcb6b0c15e73ecc36dd1a95d364399510316e32f64a69b581c565f00c3936a8af2431e955a241c06a9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7057dad61d3c6f294dc9b53ab92c11993192ebe14fdd66a6bc8e331dcce5b85af40fe80a5633506fa604e1081ac463eff944241569c4edcc5e3bf90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23c989632fd6f6ae883c68c596dda1738a7bf242dbc0262510d38afe8edea75a63db6d4fa1c9317bc40a19d0cf0a7d7e9a9d48966d1c4105b7b405beb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33c0b48c9b4a0deca96eb59e71fcd4de6f2bf1fb44b03f7fbdfcc2131f24ccc4ab7de31e123a4ac98711ef83bd6ca3dc88ace31b6490ef61fad97f131;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf9d410d36ed0c15fc5f804cb03709acaf4e8afd8991f9a8737fe8aaa2b90bdebf974278302c752e4acb39975392e191794d155790fa562e99049650c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd050862fc790a1db5eecb8cdf2e6343cd790a48249fb0af1ee7517538bbfe486259143aa1762c1082ebc22380fed9d5e9892f39d5e39f4e2e9837a632;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8267bebaf34ea701e18f4554c6f7c34e23a5ad24b7eed6d76ea6b5bd11073bcc26a4e7718ef55c42796e165795942f1fc4bdfa4fdd7138187ac341e11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5022c9ca3d2cf4bfee263b4e3aa34ec256a577bcd27864dcb1c623ae71a5226de537eda0084260a5c718ac6c756c8c5572448902ea6eb1a9a9c22097;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1287aceb157bdc538f9ed8d97b4efb9a7db06b3d1b061e8fea49865a1301b538c56edd57ba6444ef5d765316b3ca91e6a9fdfbf56080f12d9fb4b9eb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc640241e3e115b62ce5e496dfd1ceee684dce9148c8e368245aab3f713040a700a1f391a689dcd000e1341be14041e2f709100413890729c8c759890b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ddec4eed7130b5b818a0a0c4811d54c9812eb75a2f17995ac485d0a9b005ab3066f609454168145c58be7077e56515f08cd84f36f1e5ead02f231809;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd0d121f1f37d55d04033cd7273bf3c942138ebcf3f8358e1b321a98ce50cc17ca95577daf70518094cd8a583328f3229a906ebea4ddda66d89f0cf39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17e2761e2695f636185f34118a39234694d14c2f9fe600539dfc46d4e33f389b39c32e47b830c865a9155c50a031246d414e5fa14b5b51c847df4cae6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbb0144bb25359e2c620b6e5cb8370f32e852fb31d7e7dd6ffb7963bdbfebdd39d0aa4b679465a6b53181e2f71667d44196bc22f2320212b0c58d38d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he734cf4d12e44e64a5fd1c9e24d6a3d6767d7a21ac53887fd60edbd50083db3b33d8791ae310f33b97d143cc447356ac36d521e8c9a98dbcb39588d9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h451035acd328b4e367ff4f7cadfb6289cb14e2acebe7dd219bd6b61afe351415673500404df25f3f9950dc1abb5f90ecf8457bc5ae7722810438a7609;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2ce72b7fa0b5060a72aa95bf98c0818afbcc44351be35a75e033a0e09c006d79af72c9e709d385957b9353e28d3328c976ad270cfeea0f4c373ccec7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7e554d4bb4a05243d5040f51eb298664cc26160a809bb4a8619097bcf4d6143c1bbc2f490e4e28ed8dbebaeb48aff3ab7ee0de3364b722b3304a71eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h814ac37cb61f57f22d2bdd29e13444d87c339735df67681b04982e241e0c57872a19e7ce48db4f151f127e23d1db88069d006f2452c4427ae49318c70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd04bbca2a99af146b176839744c1410410e9da4673bb651a4f29ff41f5717c0b347c2794ddb9c3a31987b831f6fb77d60e8b59d6bef969c2d3d0f35d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc618374216687577b5bc931f126b6512657f56f4e58af68f40c35fffd6142b72c9570da926725e8b61db8e98e8c407cd1c6eebac7837bdb3fd3e5361f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f91d4de4d52924f616385003f2f72c6ae3b334ade4c75b90e48aa18d4b13d00410475051422a27a0d547f268dd92e040ef804f32d449794a87f0f6f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdd2cd93a53ec656ef8056465f5655ee2e7178f8a6635cdfd44faf689e98cd822fc5175d5c224da6a65a42bb22784384fa146f139e835528444d532a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d890dd4afeab44e5f3714d9ea961599f001ca8d02d0ccf8b39f6c0501a22ce2a0d53a57eec7c0154a5575b9956fd0b5a0f0c6eeda4e6f87b6e4b6c00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h578a32644e263fef09e695690b6308586c114cd6d4fbe932614893f2b8c477583476ffb1a57faed934bc5d41f3bd395f7b3616e68a94d991c8ffc02c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26417ac3972ec698e8424e7cd88c44c94ad2670acdeaf592ac1465520a2ab0c20538bd59a606d0c50df5799e51c0e03e877a21db2d3cb4eacdd97ee6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h140e96214963b83f8b5ad4db398e27961f8ca52a2fc5ef1749c9a717db7ea63882bcdbb848ce53bf94509fe5bc706a70546dec7fff59afde72c22e341;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2ca5e261b924d30f44d79ef1b2caac399cbf521ceb681583d53fd120252dc734ec48d7b44e8d51ed9ef98b537d2a98c370e6a115a9e7f9ef8ca74403;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha12b7b162cad1a3febf43cdf672013428295fe03b1263abcc32debfeecf97bce8f18f2a52e72ebedf3531906747247a2cdf36fc347710fcd4a6915334;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e188e045137a1544779983cec32a225277a5747b604ee70dccb9c02a628feb77ae1c7265d7904d53c7e4decc0e9666d6c3edd7cc887b53bd9e11d39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc18071432d3b9ba8968c9cbf8d98b80f94902372a61fa21f84a10a0e3cecf4f674f8681eabd6880cb93eb79adbbed10f936046d20e6937054dd8ff4ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3bc06e7836a8703546e2828be4837a1234b189b6035ad007ba45cf0917e1d8b5ac399636ae8d3a6d3b789f90b1bccaafe4ff5f88b12382832d969f84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f12f51f010030b0f80aef07959a452d203971b32809138f63f2fb486b3dd77b10e081e156df746fa4735256a6f1af083572a4331a7d635a47c94f60f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97138cba5d30b1cf8e4f8fed6db573200ef272e3ba253e463261f91cb75865adb0dd8e8b20e3c1a682b414656ebbcaa9fe6870d52c94818b39a352922;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f2e917eef3bbad0a57d6e2abfe8d1b33816ce9ed02f826e24ca459a8ebaa2b0b5213a8f099ec2d2e8a3841f7a2860e3c8a58c7c1448a0ccd32b16a6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h734bfda52ed89653f8b3f0e6c91541d8d0afb5b4cef9f4ab65a51bd1818a82c0528ef5de8de4e788bd25e110b14a1c36b60d630b85c120b00b68828ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fdce85df27363b5ee39f86f0fa65c96e0d79d4a165f7801ca862ef042e2035bc1712ac0591f8f0907141626d417105582d50fe664784260db3154b22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5657edab488ad5f08d8cdc9d13ed1561598905c32a2bf22480751feeb47f626744e1e024dc65e64715837c1afdc4f82fc28ffaad4728e46925e768fe4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3f5b1d112fe03387320bec5a318acc1a753b51ba10ae231d439062af79b58ad8228ab28255f317b57f769da20c3beb9ac8ff18865c7dba1dd689615f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16d550ecdaf58adc438293d44f64a34b2933865f719cee2e27143fbc36cefb4dfd5314f7b0acb0a4ff4da89cb83320d3600cc916a968f50b3dbcb0316;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bdc0ddfa8a7a2639e650067026b7b5a739f3a9156afd706c4eb704174ec9aa09ff11a07fc187f573166dff9922a36783ae4619c329f77f782624a336;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8b5aa72dd1869bf185af9634d289fe56b17e45e9ac8b8d756c040e8a2c48be0547d3bcf2bc33175c05353cf93e8af05f24e8c3f1917bf6e672e4c164;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3756d5bdc1ad52cdca2a90c305ba2c49b2e1bbdc32d39f959fb013b021a696c7c8b8818c41dda42bd2547c35fa5d56bfba5ea0ed974522ae083e9ba0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcb591d36fa771c6c81ada03ca906d0da83944d254f46d0afbf119acf32cab8119c75c59fc8c3864c555c474ade020b45c61c57ee8069723bd8ce4bd9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3b555b425fae576328182783f2e0c79187eb24358982550a0bbb05a7a3701387b32a4fa1a2a693188081dc643aa9a88f2a8c09cc60a591007048c27c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8489bd0804d3f62055d811542f494b46c8fc36ca5c5f38be34bcfe98129971930ee8fa691e8c9f2f179dc3df51213ab8df3619a826a4102494c9cf3be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90a741c5ce00cee87be8bbf1b7ad86aa7eef317cb3215902e7aba6d191284e01d6f52ae003fb6b72514e0c09aad534eddeb3851eb5e2a80b5e51a93d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88d96173bfe83f7d8aeaaac9164f82636e8688544e6a47759d04c030131ba624dbe1e5c05e4ac7c5889ac5d6de576cb8c23a2d1b0bbe97595ef40942f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc12dc1725e12f722308ac1c362b387ef7c44f15560be623c489adef839a11f401a308f93da17663e62b9d8626d393196fd5270d20d0192ffee2245de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60faa468a2c69b988b961e0eede05e7360f3537b26ee3453a93d4f6283686855a127fc9351814cb65de1bd253ae56c4b79399ae3b33c865fc10329f14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644cdbad48b5b180647835f8d50e8e43e1c1533836cca4cfab4ec75df17a06e64492f0f972227c3859cf2c7d2d27d449009b5431bfec9ec54bc582bfa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7641d2032d111636a61c87750cb6ea6fdce27a3cab9092c6cb2b9f112a386110383a328ae96ea01f8a7b555692afec434c8c9b571766a4ddef35f067b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f665eb59475c6c5304f26c04aa94baf7b05775afafe6faff2d6d1646f67afb4fc54e473986b1001015c17b7f468ca0273e7f0dbd267824cba8111281;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ce7cc0f9943131fde0fff43bc90487d1f58b2309bef39c742e799322a6ce0292e37438eacd468d1bc5e54c378350139b658284d3f5ed68a96ba0c11c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf7ac2f8ad7d86138e076d99c61d41623488da27c5350ddc6d70ab0cc9bcf2ffc596404acd8e6d50cc1b6d9728c42d687c8405e3ebe20675e962207f0;
        #1
        $finish();
    end
endmodule
