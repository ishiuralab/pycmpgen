module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e24319d44adeb5f07f8d936e9987924ae4879a67a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38faa69b2af8f1e17653a2980a876dd6b2c3302209;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16bb88fafd84cbe8d0652e24f0702bb9b221e35d58c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee032aedd8310c8d993d71a066c6d41ca8c8b4d127;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5ccea2ac13f72d1fabd95c29caf493dfa1365030e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162145fce5d92566975c99d8ba7b7a53d067e07e8de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1971e48e669304bf30d4521d94f3e4b389fbc59df9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19716ffb058402090055a69dfc2848a44640b717b4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157a7f1fecce3b4d188d7709b6d1c2a3db32c9d377b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b6077570f2ceccf40218044d4af6cc01a62bbe2d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f2f6ba5a0deafea0c1609143786770e7423f97d24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83a01e35200714e21c563793beab98fe76e24032fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7741cf3bcb7de74a56c3186c4521c19548fb8e538a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha548e3b16c09108131c6dc3671eb2f5a463ce28673;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b39a47f7a22355149d0fb7e111fdcc410b9f0bdd7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a83fc96189e40fbc08e13927ac6aaeb24d2169baa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13678ff480404fd218d09b3e0fb3f62a58ff5f8b95d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114d543325df6b8656a19bcfdc1af2e95543a29907c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec52327d2141c5929a2fdf1b56bb35fb01b41fc534;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4762d619869f086ac2c0bf0c3cc7b4947feacfa3e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha74e942cb9eee86d4e8022e539720311c2b95e5f9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1390aede7c1facd786f374a184b50266c368f0d501b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9df4563bcbddd01fa5497cd7fcf8a4504130c6d469;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h559a6ae01c6ddd29beac1e18333dc5be4414a71c81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86806f22b101a9276f7ce01a918a701f52afe080d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he60117199101e6e9d82e51c529460e34a3f1508909;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5439210142e079031cd54d22c879a0da6ba1db967d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccc9394d162a149862113d3fe1ea911b8a0054d0b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h696ed89733ee1e5692f469ed1d79e9b0b0600c37f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c98e55245c2dc5548b55fea96df75d713a840d0b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f7a84f98c47faf4358fe70d21d3cda340c9f65962;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf28aa90669f432077210051617423eeaa72e2885b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195e890d9c5b92c470a6bef41479341364d12f4b09b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f72b2de109d4e288cbf766a6404bb78b694db580d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bef26f88ac48a6dbe1d81c1c4e9c584a5870d2694e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa346f77e9fa91b7efa1900a5c32b57649f0728e7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2309e3e777e8fde90fce0332fe482d7b1d34ea598c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6b5b26ab97197a0860bbf05ebc3be994a92fa3026;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f93a62da6f8807c92257ad4570c6f88c090a3e45b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bb80189d95788df50ed40f31950a94626875bde3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1040d0d01ab370da84de4841aa0812373ab1f6f69f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c4e1e2c734e828765f5a975aacd0f300611d1e653;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75b99032eb04753dd619b71f017a75463c17c5d427;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h268519f5be0b1a6dc75ac08297b0c29bd67731515a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3276c079ff6651c89279ddecca20ce5f8fa53eaff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170e51bcb91acb1834b9d4d1fc30187be818f6077a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9bbf9b69bb39a58b301fe866183822d5db6a011b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h43cc8ea0a690da6b43d4e7361888c016d3750cd448;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5c52e6266ae7f310af1791a199c14b97af5fdd524;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190639d3dfdf5348c024d82e871deb1d00ed62480d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d884b064c3aaa9147cc1fefb79d4fc2036dce12efd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8e693c96859f1004a67bd4cbfc3a0458f7c900787;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146042a2ccd740cdef3779354a75c7afd3e45de12c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4bba723756ca0d5f12fabc96a32a6e6dd93be634a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7bd1274a0703a99f03c95d130d7d376f326a19b82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137dcf80050e57c6652e6d7d1898f28d69d2c528717;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e45a91961750ba21397ac0682511758396c122d96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193b66ecf0e652bdf4c766d1c56d54952c50039c0f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1765177dd27e5cf4a4c735c0572e12193be2dfbca8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f271849ad390dee06ebcaebf8dad5781a4308d95b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd24bcbfe732721fa0db4d3c864df64d3d3d023df6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f219cfb9cdec88d757114beedcc282fcba60553f09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81ab44cc9ba6966005cf3caf1b420b3ab29808b54a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc59055e8cb1a16598b2eca55e8c2cba515fe3014f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5afd39a12ddb3a9dfa4ebebc7dfbde57b9fcebc634;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d243492e108493842048069deb320b034951cab8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f86a22ac6a62f07046ab70123b44cd9be9fdd6cd09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52b7d183704036e2a89c91b66eeb0cbea4fac6b03d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7010da2324b148879eabddef4800ae7d4609751121;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16beb370667fc8c832650c8167442c131a81a734905;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf41971e222d6ed11cc845929c9ef0f1173426ad72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a1549146d42aaab00f6909c0112a618df5762e796;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7566f7e299afe730440a83f02ae325410829208f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14eb0a272dff65cca1987670daeb2bcf18278f7777e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d97f0bdcdea1b0059e137d6010b7ee1dd15ca64aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17cd2e18c6565ea05b6b10ab31836d53be325bbca7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9fa9342e49869c138df88f06cb2377aa8e149b6e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h495013a3f053fa7279d21b94160bff6a73003e74c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b7e272476b08277aca6d922eed90507c67f4b5e6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heccce13abe77cfd102ffc790e74d416d496bfff825;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec0b6e51dd11067e92cb6fea83dadf17a891d0f835;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb54682e5ab1d870a167a248e8208a29fad7c35f238;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fc541041076ae7198bf96ab6b5bed8c4cb9819045;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ab618765b13e4b85555f75d7d09b9054d77ff8540;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha96d1f2503f1abe8e3e8366eef1382a49237f87f45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3406ac4ad6694185230b5e89030c7a8280db700a9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dce6ad39d0329a64b6a7e18ce97a1a64e5fe7822db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ff965f3493b6abeab6fd78a25bd4815e35368d843;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db4f4b2a0489e304f5c77fc13caee7f91e7170cbe0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hebe544ec01f0cd506ddc02ba61838f6bd4aee69c97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he42f4365c08b9d0fd8a3743faf7203e9bfe4f75400;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1719602566be719938bbe1d348b00e7de7f4db00b51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac4e1b7065321aacc416f3d0e5d2296bdafd1e1ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39745bf1447546b4c41b1795f8e0dae70f3e8a4335;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd621d181c1a515f4cac541c4e59f69adde21465737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1900c598dd4b2e8487bce67a8db8105663cd741740f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc0f9c986a2b8bc29f5bcee5c917a311e4551a774e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7271879d0a5284a3ff0adaad3c0f8592b03cc4754;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ddab96e4173170063526cf2105282dc2539b833d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5016331a5b7c833e7daf935c6cf19c82ae21a2204a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1123eeb8b15923eeca42c3f4f3958905ba277a55787;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9dc4eeeb69f46e51a1d90e2030b4a5161d73b7e20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44d26e7cdaf5711c077fd94564c40f7af4b197495;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1257da6f5a6e04235309ac189150150f9482d68aa83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf33e5aad02f17d8ab871dda23149ed0337bf8a9cba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8201d9958f5ccfe35d095260859e113d224189631;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3dedf2a77d7b760a034575b38f3b500364c29a56f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d47390acf73d76f0c892bf17fb2efa066e4f8e1b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea32962f6d75a8d55c6b619b78a02a87ca4f3e42c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5732cf1800f9792a167254a508eebcbbf705196749;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de5ad27d04b32f57c103a01394272567ddf2c94a23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15451b8ea57508d3471193c44dd27b76311cbc999a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc1c5f8d2cdce1a271baa77889f5ecb21139fba199;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h586db23d5ae41c9d1f620702f33b4e68a55d819ccd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd9eb292340a1b40bf22b614e6934fd2ecbbd66845;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eaa8fe8472ad5e8e1a302df2e35665752c06273565;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15170292ea4b75b6179c2dc1a3c0a93cdaeac002a77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1569a09fae4003b5f0db921963ea3c7c2e141dced40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h713bf6e2b6b80f1d0bbc2c82e1b26f8bb247f0aeaf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb56d6986e3a006cbc9f6f8f32c4c59289762f1586f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ec66b956645924bcef8eebd9ff01780d38f0b161;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae8eca26a5560e1461f0eaf77249dd143d7032c652;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b271ef3984b24aca27937506939e1625a13e2c3cee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e92e5560ea68988a0eaaa9b0d5e899f3d88de09a29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h745794fefe1e59d6b178e64f14fad3a1f3692e4b08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd790670250d05edc9dcd154e8066fd9435c7976756;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9dbef523f6905c00a0bdc768e2741f54f2fd3a18c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fbb43d197a82e3693ccfe0ca50ec5deb3efc6c2baf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1841bdcd9ea6363d4ca3f3e4f05ef5836ddb948d265;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he35f97bbdab5b190e0eafe27df2d47529b547e708a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c3003b68548b57475067c35796ef0d73884d73571;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ebb652b6a5d6cfd032ed2f379feb4f9df35b89628;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e713a68c3516a51aa3a9dc9d2698dc4c5fb097524e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h829f746dd20c56290890454553ab5374f94c12b24c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39bef9c56ac922f4b6a0e547e797dc8b9047d437fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f55db549ca0c4c87533f414b177d99078dff2e836;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a1bda752e4ef447bd6ee3db4a50eaf8a676ccef6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bd406db65e7c966b11696cdf22c45248b0e1ce6b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1131a25ca89ecbbb548425c4e079995a32ef0173d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f08583006d6cbe9bba0b8a6fc77a365063a83f636;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195be020b7d7cf70f67645790da5708c17c96d90cf3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19494f524fae7abdf6d217e17a25894588d881df60b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148be8bcef1cdc8d136a321cc04e1686e5f5dffaaf1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10fbd53f779a13051e39d19979b3c95bb87c21db8c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1997430aa2d5dfb1898cabc9efb9d5de08364446a25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af5fe5748f120de6157d654af821e36a87dcb4bea5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h251bfdf5d0d7b73464cf58a9afa6dbb05726fd49b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40b60969aaea0ff6a42feb5c132c5e122e0dae6ef3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffbfcad036d16a2fcead7cf679625da5ee79f8d3f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa69a0e5eb41781ecb9a01e2c0f95ddd6e90060e0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he203a9712a13d0b4cc5dc0cc1b4144df20a0c076c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62059b0ac990a726b2190e87db6ddf51dd136d139a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b45330145802ecd043ce9b32ab064ec95e8af1711;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12a02d9ee599444d515a767870dd19fb2b99b4692d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5ed88ab2dcc6a3488cb9c711d426e1eca7682fdd3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194999301a0d0eab27888c9981b045abc5ee7c5fc3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ec481d346cedeec67670bf53e2e1fd4c62753a214;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb47218eae55b9ab8e82ddf3d8a91426f889d80fae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44cd53631b3fee9a509d825845980ac473fe2de1bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb243934a3f02f2e4b7f50a720dc14a5e2fd8ce2f96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c857698221ada8cdcb3dd9bf51e1cb289fd546ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174948eab00adbaea2c24612e5241acd508d9373b65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1615a9a0d95248f90a051c56faed12630a5fb99dfc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164486b5cf10bb57e7ca22299338819a8b904f94fb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4de006120d89784a696e38891f304c1835a1a14af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b77a758f97f76c2823b26e57b872e09fa35847a06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h864b6b9cd35a33391e943e5ee2f068205328a243e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66156a32a87ca340cac74d69a1f1aecadae6774457;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26c02491d87449e3e76710b03b960eb250cf1a947;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10830ef80cde5e1d4cc2d955ce04a02cc094236729e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113439484ceba538139061195b6b16a45566914d5a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123f80487d3c106fc4fd7121cf3613b05c5a0b4b63e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40939c3c430b11b651d683bf7476020e20dcb35053;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78af6ee528dd4c5b3b61edda6b0238f3dd87d22759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c88649dcb7d28c20e30b27dd7611030d7a293cf56c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1a7d52e429926687c1915855b9c32c4a3bba5476;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de6b55f33a722b706e38c7a192cbc986ce2de6073f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb82b58ca74777e05ed6b2b0ca1f66fdb62f8632983;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58594886c565be13103d09491e9f85ce1f38eec6a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15bcd980f88a23d151a72899daba4c70b80f9c1c46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f381a7a627d2c9e49a527af88976627f5fe6b5ae1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2d5c5b612c138b4ee9d9820a876e79d7beae1f4fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he36093dec5f6a3ad88d79c9ac498d276fa9a0e4c7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b0a2e9a5138482c08145b8d686c1cdae18994beabe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6138a7e842d0dc8f7dae95536e31d8005cd3619c9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d039ba0fdc2fca4fd2c619c9f9eb29c45dadf7f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83f7898f21f6ba4852cd794ddaeb944b1f5672d9d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ed25cc59436c30eb12de9e4ac0cc30e39a3c8b035;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c608a660e538359276a65e000e0946371e3ca3781;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0a7dc29065c495ae2f71fee681311c4cb9522a7b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7220ca1eef808e560beb9854b39b6f1b6607a538b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bac34a3456009fa17ba7288cdec33ecd6bf3f79b50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5353558deb3fcc66cad5c2fca54ae56ee308e0a8dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h984cea4ea450b63ec3e7d072be5a4c80793c615337;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cb2ebe886fc67f13dffc0dfd51993647f19d962a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac5f436779cb83e631287ae3f4ab194f10a00e4544;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea9767e0a6c3972e285ceac14f3b89e7cadb3f3f39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f5b88e81925fcc6e32b5e5b0134cb8e7ee2314ce3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8f8e385fc3572b6f183f94681ea9817aa77a17d2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda6a9eafcf908ce0eb3048132e8efc3d3380fdec16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he078a2b2cc47f1abec7863d0236c2779d5e7a2281f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e835a8e4ecdc3ac17a96a03ebc371cb822085529a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdced115b19f88e56bbe5beef11cd2888518a48a3c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31be49c2d8aaab3a97f15bb291d53a4aa93f8acf37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a26afe043b3a8ecc3f3b2befae03d15b26b3a3fad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ff87e807753b3cbc3b50a319dd7e5b7fe39b9847f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6fd3a1387dc32868e73f368319a370ef7b3734a93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha54e9fc731178945d53ceda4801bc58d87285f524c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144df8182893e5ad2f426d0421dbd443ef140012a87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4a3b506b5bcb2cdc29c8c3de39988c3498732fd78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3edb7982dcb88d14d69f20b7c1240cb43d74916d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159e794516f2b2f3918324d3f32037d7942502baf8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f37219f85b8828b015ed6da602eb183d772c765766;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h620719a82a2be0c842655e6ffa2f65dbac98319878;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d684fe08791f613f513550575e495de6825af04ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13017b476486205ccb08c9ebea7e9d5cd66c649c121;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9d8421ea99aee81127809dcfbc85c42c2b7efe302;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3ef50d778e9273aba462e5fcba3bd66390cfd415b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f7f93b4291a9ed13f320222885bd5481d45f08cc93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62f53c7f36e97d360d00a32fef5c4b3e1571e0edd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1984366d1b4fcfb9a671d3c4de17303584d4e99ba44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11aee8917bef8622fea38e0741fee8f1dd66fd69764;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h667543be2d711fd996bc07de1a7a5f3209da026ca7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd03422f82afa245babc7484bfaf2028538cef1615;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecdad492cb0aa02fca4a567f518f3e4b31afe65522;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d04900ac47b78547b30dc4da0648d3cc766f310bee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ce204dd4ef3c38a6a81bafa7fdb1d9a29f3055095;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e26d3dbc373d60eeeba656a31046722e0e3bbba5b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea6b605803232b88b8967ec63162e1da9831e51ef5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h468d98a00564ff0a7770eba722aa697ed4ef178d79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc0016c4dc600d589ccf3d1c4312efd691084fb912;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c1b7b9e7031aad720831b9c176160fb3b6b99387b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68617ad685fc0a6e2bbfcd7123529131c44b7f9b8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa43faea0dc23dcaee912cbb7183c2c44563be11cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8876d7d427e83f74a30bdbbaa7f9b3027db26d1ab1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc2215b0f5873837a411e5a125dc48f8802d1c5fdb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f63b4f0f4f1293dd0441784c2ee52a474430c7d6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4027cd52b8d7f25e180dfc368e15b2cfce25b9cdf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8fb2c8c1ec905179cc2ba3fecdf78d98901cb5a2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6eb86a8715d95d5fe372700bfb9b39a77de16a7fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d84b4e1f99e277814890f9e659f9310e3b24095c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he462e2738eec4325d77d08fa8aa10f6c68e70a3948;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a0a4a1ef8cebf1f99aa30aa90555dd0b1a3c6f8cb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149d5c12258f46e7fc20565179dc25b10b60cd070fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h995d49c066a739d2f4447b5a5528fd19c31e9903af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1422700b628d4d8fcb94937c6955a8852c0861bbfea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71b28f3d770824cbc115023dd2963e875361815d65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h487834f497348dcf17f9e8ac7e23307d6059e8f034;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2461f4acc15572d13fdac0019332332227c282a009;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbff55b1e475252d5b7a3fdfbb5103eb0f7c0404acc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1d66670046cd26f890e0a4a1cfb1c4c2d3c2a3994;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd732bd1d7a4ac0b5fc1d875450a43c2d650b10bfa1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1147e7a7a54da053e722aebb76fa786adfd9388bf4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4498f95e1fb1a667698b4684d42c3ceb3201c4eb9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h139231ae84abf0b07fddcbaff288c2f477d95ed05d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1644fbcbb89f34fcbcade290e209d55af1331c09d24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1934074bba3efd4905edadbaf214d75224598c6a53c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c779ada436f265d3293c95937e41e412802f45ecd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hebd5f8e995f342ff5c33e4f2ba32a2cb5c615e2448;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ce1384847d0c91ac32ad6aa7e0a2349348d364b62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165f97268c31896b9b8dda8dacaaa64dbad5ab7163c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26f48e5deaed4f73c0939f7db0ac47b37bdc555278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb6abf4e8f3887f8bd54c1361103a74834a36035357;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16df24090820fdc0e5d53700e97745d92ceb3de94ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcba22c41f2a7b965e04863ee522f53d0fe529ab62e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6b6cd5d23ab4f41e93c10f527c50e3e8e154e43d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146e8738645049ed5a145add755f9527e9dc96cffb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha91c15413f53267551b0d627e8028ee86596beb29e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd37937482673e48f112b4a4ee10b1cfa28582404ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1deab8f3339eb66ef0e31120a999dcf662970a3296f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14550e42f628d5894fc7db139eb2f9b8c0330d9873b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6db0d876764bf9e0ba366bb818876a578b3e0ef3e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199cc3492a202702c30e19aecb83ec22750c3581e88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17cda41a56950d874e7411f7057e54f0d0a00ab8f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf9143fbe898c948e154135cb40f3591ab47936e267;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1040323b46e58b248f94ba393185eb2af7b312fb4c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h771e53f1e189916e49a7fdbc212aa38e13c2edc46a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55cb644dbbb7bb8698fe3a0ec69f6db7153dbd1b29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h490945559c1e2cdb49ced27d0f0cea18ed0d2bdde0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102f45da5e5ec6463e154f2278ea704c97eba04aaa9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c283588438a27cdf05fd9aed069172f0f5a15f606;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1541396c8b88cc7b0c80ad8211dfeb4ee502a33315;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11981557fa1bbc161dc735051bf8fab640a477a3fac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4173d2aeee8f6886d1543dae818bd1544f9b4e08f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e5c1302be3076398a2434fd084f89561e0dce2105;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1904f6bebd558bd5af55ada4d379dde1c8bac80d032;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h37bb33574fba1045937a2f9825e47b84ba0bb767b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe1d953433cebf17c72bad6fa600ff7a7ca33bc496;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13422f5068c30df2e99d633d781069f5882d6c725eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h974cdd71e2afd52e10d7ef37919a72d06e86a4e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d29aa529e99874613c51c04556373edb0a863018e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fd5d764e925ae1add7932498b548fe56b061b1d31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192bd6034a53259ae4b513d3822c40371cd5d3be0c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4adcbfef5509acf5d352e8245d76c32b784ca23f69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fa77701a78dcc14ee88d6e4390b8833be481b107d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h446b66fa686907bdf940eab00df5bf35fa2c8d0907;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4edb5fd4814a4e4d77e0f900a81c01aeb7f341132f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d9889d6483215b1e01abd6440ab1a1d495259fd98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe4d1701fb0a7c052a403d000c49cb6c228ac2b508;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d9769885b6af9f4927695be3bdfaeb1e2f8a45c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h310cd5dbf3bf639af535778b5e2755628275e08f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h465ab05b5ac0b988a9e2b9a29aa66394e166ddb6e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b898a2ddafc0e967c32ef3ce7a153e4630e5114b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6494f1eef0e4ecb0381e4cbd6a8735181c467ab89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36ab0ee4bfe8d04569719d098f002837d8ed269a9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8fb7d848ef52b836b5f36b0ceada0f5aeca5f5cf74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b3a9297cc95b1e22d0d7bc4fb89fe23d04fb3f257;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a22129d6baf30ed6553e2baea1861f9f862af6cf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4f459300e652a2464da63c51b96a1e68875f78141;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78b7994748587241aa9433c1799f58384db9ec424;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123786fa2bb79487c55e865f37bb1284e43109f5ad3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c6ed47d40056761dfb2d469e6ee1d132e78d38a7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b3a7ef119eb5ccfe1e09d3c333a67300de5c06945;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ec064f06a8fe19a1f732c9f1b8164233cad968ffb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4ea071cd7915cd6fa01fd10eec801afbb926b8081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5fe5332c2ceee5e8cefed34c327b5adc4f8451fba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e8f71ffb0255537e726fc8dc3ffbc29e9557c1e55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dec888b9276327df46eacfba71e1b6638276ed9c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3051b37a10a7e0fefbaaa81bc8e7d2702c9aff4644;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1600fefbeb995f3b3c5de6644ff5b59d6a8286b3375;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2c799f5342aef94e8e4269284e9b9367cc4579262;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122c26405042076666c62ebdfb51cdf16f84cd3eaf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17eeae48a9aa5f7e92bc040648ecfac8897e0b9e540;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce77065be6d1e4dc9fba8b51e8f026f4d11bae774d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187225a40b7871c23891150343c73ed351c62ea676b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4d586070c7c26ba40e5dcdb35fc15567752e42916;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h700dc100dffe5c9cf40073ad510ac08def1a9aa454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8bc842b8083f72f1859714bff613ee8bfa8a11dacc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a90eb4a46a2169285ec6ca353a07dad9031fbabb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha051e836f7a24b2563fea34832c87f7f7a16ebd28f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ebbc663edeb5279d5e43f45aadab0f8ae98c1ef35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ebce7cc966c5e7881d3f6bbb8651e3e19ccacc7047;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1807bc17e06cd2c20c088cf021aae3aa7d931c7c832;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169d007f3861c66691025e157bf946b0068bc636c77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c6ee9be52e4bdb7375f46ccdf980eff46bd649219;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74f2a74d01a146adbcf0e25d18eea7e22005c233e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174da9e7be3593b74b851f3a3ccbd9b15362978097e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0a380b9a2e7e0065bd0a915acf19ce92259f53124;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he05ccf33d8f60cfea8594487eeccfbe565d5d82654;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h886a91ba96104516229d79f6a40125f4b71e741d76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa8be12aa2438de5c7071a6f3fb1ad9789dc8d43be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3802fb3c4bcaa9dfa3415169f3d063f46c71f43864;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e93a60ac785c80e7c317fc46097713eedb03424269;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16fc9b32cf5f314083490f6b1b2bf0a4c1527e889ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cde40b64a4566c635e3a9316492d377f9b0b1b586b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1040b6683ca188fd42970e969f5958d7c3459c66f4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7f5a8e412b6c670e9559e58d80dac4a4cb34b04e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16006d821a19113e0b1c889c6cb484f3b074fcc44fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ea33ecd065c1e0b9075602b262a30869a7a6875b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heaeea15f6cd70d31c1aabc54a668c3dba0777f5aff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107bf641ccf5ad5e754069354711440c8653db0e03d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192cd39292ff070649847f341876b0d736ab88b56dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcd7fa091e78461e2fb9c2304e6b330664cdd441d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e9a8277bb0b2cf9aaaf2b7d84c743033c5549807b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149825820efa7a08811e2856ee70f4283be6a16f019;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175a80df38c92cb8855a86652f0c5cb302a242ddb9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ab1f67187d5442ab7f9a269e83f42a71361e87fd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fb4ee0f1a96693dc7ac7c2e42407433f42df6a03a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134fd061a43c3022c8ef05f67bd405e273955ec77b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e9b421acb65cbe1524517bba3d305156dc9c4d73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16945249b40ba4181d111a2807e4ea90b1803ea2eb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199db78f1884791cdf195d593da7d80e6a74662dbdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16251c6bf0c691a9b09154258db77d8f21223e90e56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e275e5c47ba67128c42d292678107babc7ac46dea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1162e1b9c732130fb2ea2da847bf125dec89a4c3d40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1959699a339cda286d532f55803bbde22637c998507;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141b6677bc4f302ec7f5cfab2be3726f3f34b10307a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef10dbe4edcddffa3d0357d64307039a27c87874aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf886bc69737ee36219a9ee7b4b44831b0edcade407;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8259292253f698847f627e1b5f645efa53b1c3cae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he93ac91649f53e9f9d65d310a278eeea8ca7bc16fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h270fef0ee4a014672a6b4d24e680279180125f8c8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1328c832429738fa4579c4cc5124f65f51104fbd4f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b902fcd556c79dc979d6b1eba5f867a7d8dd5d7791;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha68ff194e50266e84cf796047b631cdf14290b4c73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e46b8eb50dc6323395bd1a29ebbdff93d44babe196;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c97c109f387a050c1efc4988ff39310b2f8f9e87f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17568c2f205af1af548b64699594f85e2c749de0830;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172c13b74781c76ae98a30394ff03c7cc4a4a1c9452;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b5c787484c2a37ee4ee97101783dc6db114515c86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12990d2e484297f548221dc203e812ab5fa5a32751b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1313a521f313532f228b38006b08a8a8c76b1abab75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0ff9a814130b6c7cccbdab85c8aa255a29604ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdae741cfcc875014cab1df86a7a0b73338d6f98b5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2858b551374b83cc0723ccb056e6d7e6d10514fe72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14aeb61a78167c79e6c2a4a25f3ee51694f4f9acc78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a47706c331be5469b6bfa8b009ed1906268ec887f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87f49f4fcbc4704698aeb465d507bf3cf4ded857fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he566d24082ac0fd44bbc24524a8905fa4ae8892d42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb84834fb554a67225bbc3b5257753301098f8cd62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13878d77f10bab2dc9d5179f37282bca0e88ab6b99f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45ef5fe79ee57ccb924129e846c9ef2ce89fb7f083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h925b96053a42c082af5f9dd5003ea49ffe26592411;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132ae34beffe7f69e3912e9c192f00b2e3955db417c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3c5ba7f7f7d5a0bc773b728d23c95dc7584fe157a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f50e7046ddc81ba6ac045ecca2e70dec795170f2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb52bd927b88c6853f44f8ef23fa44506a8ca63fcd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a365ea5320212cb655c3d46cfaba128508896057b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b993bf018c018dadea44612a4c56be5425e449464;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f753a442ef74c44b205dd29fdae306da9e419b707;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d21ad0011b6277c0ed3494a8f06edeaaefda12c4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4a784c7141a4214df52f1742a7887d7126c3dcb49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf9ba695d6ec74352d42063a0c333aa750c4722770d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fac86caa62991db29c7c5f0cc20c0814472f1f3d16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h967110954d11b625edfeba616d96e1c50c992a5d13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f76461e4b24f42133de1d634294f964d8c9f0a1e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59e135175d2281f5e416c32d66e995fc40179c7244;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184fa612e8cdc7dbbe912412d8db5f792e79537a86d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6b7b55b56d916ae2bf839a540313673dda2207fb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c57bf5e8c035cc8c5f7a6232393375a86696abbd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7592b5145ef4bbb688ed6f54f36f434af42437c0a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee34243cfd8ceeb70b967beb30fc6476b3f5f4d219;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16796b947e509f76ab80215436f6eb2b0818473e89c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc90c7cede713f3fea9a2b23ab068a7421c06486e40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b051b61a6786c6c73617012123506ddd9d5f6cf2a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9cf7b35b1106424934f183d0a5460acad9a404565e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123adcb2a29433200155944eb176b59a6bc26a42bb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75ebc3884d9b493b867049ddf728954238093cff81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24ec07f46e725c2b4af75305dd9f959d68a578c20b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdce4c6f6aab83e0b2b478f116644b4f71e8c01fb86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7a52ce34a689f927ff804a29e2021732cdd983948;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9915e0a3bdec75ff53e9aa86c575fcb0a9707ecd8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h932ebaae7c78730781c7d93de857c56c67de2f32ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fdd5e9ad63b98f90ff0f469042b3bec97674e3ae9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc11fead7b2bdb6d29316410f53b4f8166575f9c29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90189f1057ff615358854e9b3901f21297fe1dc023;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a603b64fb68355b63167de1ef1d77428b1f45e27e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180161465f450b5c5a3700cef21a630877fb257fa20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133e506e84840780b540bc58fedd56506f978c7a2ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc4fd6ce608784fb2aeed6be67c4cf9a10438872e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb50b1f877349c05d6cff10bb6cf8d73fe3ec94a872;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1474f70323fc1ec4c3cffc4b6ff994f265c9b92ed46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd8391bf1f6304d19512e48af81a5cb7f6b805e587;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1736583ebf2a935b5d7a18a01fb2314f9adfd3b096f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51b150237d2e7691cd6e45768e4780c79c37944d25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h654d7b44e0d31ea00ace9a05071c686f3750f8eae1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130fb614415f5b772503da273316e8d29be33789f76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1022aca965dff96e2cb54e73c27567787897dcf7d58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ebab0aa6e7b6ce3e6091f52c344316e3859091fbaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127ea2459f6e788cd40be807cf26ec68076d5a50d52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd185068dcdd8bb4e83085fe3114b7d176dd0d88b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cedbb610bee686449adb02f53a6eeeaaafb5e0288f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heefc75c97622a5a2e5e94586cfb8f5500718393413;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cf148125fa809a700a7267c0732063ce79aeb797a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11aafb345d91de250b1ab666fd4561a8aea41b80729;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f2d7eaa6bcef7db66df631a34b9c2c4809e640e37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3491c00d7122eca2a529f0b738de5745be51051046;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd820659db7ee2b1e8a3aeca95f77ffe71c172cc90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a5ac1747963f423143b4e25d3e312159b9700dd28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cc65ec36bc8445c6bd280170d78d006e31dc0bc89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea5b64875b1e77cb6ca865d668f7bd5ced810bb490;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0c4fdc64d8d92345b3dd495d71f03d4b716d46744;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10cb8d0dcb004063bcfb1c63b88b9f9a9dccade2c7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df6801f9f5dfae2dd90fadb6f5671a0cbf158e3ed1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bbfadf9c12e141efa0a9d1caef4401b15a1b26ad7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d704f928d47f6c34a9206955ca3a076ef1624ad14e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c0cee48cf3f1ce3628d0c7c4d219c52508f3ebfdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166347a4f46826ecaead2051b588107d8cc7d18ffc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85db4bd5431092139084f4ed91bed9d9f3bf65fe6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h778043f618a160aa66f16022c23c0fd634bfcd39c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148aadc4bc735ba79a60f513db4ad8cdb7d39febfea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19996a7f17891744e2b00b5981b1dc31ebc4df79430;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b08d7e5191c5202b197b4604f41ee96f142c016f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102192c27e6c24f65caf6cac945d1ba36a19e0c0bc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3e932fae53bb78c3fba90d1af13f1e7d4333f41df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86ff46e5aec2a05cc8d21321fbc154770b9d2dc2a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c630890bc660735b4c94f1cbec8a2133c90ccea5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d88b2b9eec04182228eec31e1aa0e2ee70897f089;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1734baa8b2abedcddda1252361381cd784144a73f82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193ff86679e8bcdee84bd6cdc03e46928d43d23e523;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c4e70297edc6f43855b7a2a025b242109c724d292;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1709b99cf186bd0086d06f3b3d3b165bf971674712f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h437cc4c9e1b7b1ef5653ff028cbb45f08792561c91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72da8fa28b14efc1cf561f14bdf5371a1e8aac6850;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd37e58c95076ad21c3e1e3206c87778e12452ffba1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d96c462550aedc5c8c9e445f303406b16a3a46dc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4431228b6cbd6ce5b8854756e50c67ed2967704b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cd0d0285a24aa7a7c363228de6a5132797156e1e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5a352728e0b405e891f177a70876994962ff240ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99bcee092478dffee1bf202aae6a1f244b3b7bb9d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44e42fc8d267fed63b3a507ced0e0135e281fd3457;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78c0e9e352ff45651b665108dd74178cc6836401e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0827b5e09788664574699a0a71ec69caa6380bb9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1408d2ceb600815df8f5750974c7d69af1d9e1f8c6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e0c978eb4fcba16eeea226809adf8a8448e2745a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148dbae2cfdfcb8bbebce52406c18f199399739cc5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198448bbeef60d01f688e33eb8d3c6c8efb38a9d7d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb904ca49665f38de2aa66ac8bb587e1e8723019609;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f83b915f42088b267aa95bccbd831804474f665bca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a42f50c6417069bc3a7c49cdd75dd6472b76d5c8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94fa9560c6dc8cc3b34e5529c761936b13bc3502c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc9768a05209bd8564d53b0a3e39bae19445f5aed4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1647320a0f5b90c15904c5a7583478d5e841d4d9f39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9308129b169f0e32ca9c903d08c8f8f86616617b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h302d4919ad5c191fbaa1e871c95572a44790fd154e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e25d7793b049be498e3c69fa3243021bbf56939e85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102daf41ba4aecb650031c94fc0e01fa249f8a4d97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc5997560a0857c34e1f59536ca719b9c149d6eacf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1329eb0012434d79fbc3fe5b30dac826c2af0911559;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1612d996830a7d75e53b45f33b977248b338456b19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39568ae95ef74f94823713ef7dd1ef454bc61de7f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba4fa5a1baa09dbbceb995c63f8bbcac1c942888af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17287b925dcedcc8d21c62a9398f1cf03c6c52c9044;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb3dba1880a2d6c04884f524d216af59ebf902f71f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130805c9f310d429217ef7ee82d6e8cc55410b73f5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d8594cdb2d7e1355ee81a890cb28145185f69bbf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fa4dfbbb6b418306e639ab5d527b6a056cdb5d25c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a6a3269885a164add0002a7e2a8e15a48b2024ba8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be0736707a5a12301f12462b764e5cec21f55e0dff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ba871796b39c248c065e0d366cee9998dea3a7193;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66e9f736db2ee2ad0887a084569e44d3faf2cd4cbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h313fafb76b03f7105f88bbf394a5f8c3dbc1bf5e78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85d13627ceee35a64bc559afbb5edfee697b81bc95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6acac6436e7ac4227a457b8fd82e88ddfda8cea93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h67eef9d99c6a07659fbf7463b8aeca25b49bb67140;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1872956a37b61d53d47c24ee3e763447d52dc10cd96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2f5e6a0937b337aa5700307afd9c425c58457d68c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c28fac7b30fb446c80d1219c01fea9b2ce0b850fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc995b67d35f196558ce7937dd4e12444170df09d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1516e6865de2d0d94155a3cdc95d1e6c74e6c7ebfbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haca3405295f7f8a3ac36e20bfde69042b58d383ddc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187bf58407551202047b4784fd85276f6d4dcd80af8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8d1241ef0c9d0dbf81ca771b1bf8871d3d43909a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e9e43c87f2dc57c8cce1e0fddfb92ae7e68b7713;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h572a7e8e1409cd2eb698cc51123ba1b3aa5291dcfe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12dd088105029f87a1f5a62c3d912e0b26775429593;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0b09e679bef5fb6155e4d8424ef31a6cdd3690eff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1148047346614c89f2c34c89c38690bd3c30d4397c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f007e46b6db31473bc37de863ec0963fc6df33f2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10426362efca265af1a8f3e0b5d1ad9f45f060642de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bfd4ccb92b7023faaeeebcac39ccae731393c617a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14284e02d9d708f6dcab907337562a875f13a55974c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2f8f10ad74634f5e51afb03204b601e1df99cc5db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42560505c917752580cadb8c8b27c4ea33e1fabd58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4bb38de7ca7413a05e09b74f94627eb2b177f53e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd62eb3e7899919831f319656f937ce59610a233639;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haae6dac78b17864115c99abc607f06bdb32f1fc807;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7830062c30b74c9933c3d5b58ca51ed19ea7450ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27dbf95642baeda0bdb97f40f7ed4b2379ec591d52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hffeac7544290ac8fdcfb2b5978039adb5f12f6858a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d79d887bc89d9e25eb60d6f96cc1db57a850d0da2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a9ce77614e8ecc7950c3ca9f72c2961cd12a98539;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b87804ba18539364d7c4924e41dbe5817049ecf14;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h360d0602d58483bc9aaf0f6fa607503b69c36bfb4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c94c85bd25fc90df50f70640b6934b7aeb4bc1df33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2403a08bff459482614a810a2c711bdb0690ee350e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h188de5e659ce75f167e336b435313c3e8e005994afc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h910982e0c8b9129c6fc12e684c2fa20a8f6a04fb64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168bb76a5eefe023de42c90a8593eb38bdf68857452;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92fb9ea3ddfa74ced6f2b8e48a5a90d71d1967867b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10578c0f5ea71c3a71cf2194989980bdd4efe783d7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b4b9621e1c2f2747be68e610624fca288933a705;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e06175a33b9d004d561bd39c6753a7015cd6378e41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6860951703e15307a965e6ae6e8fc9011aec891b70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c410eb3b3494a8bde1ee5e1c7afc9d7f89a1eb2f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c501828f29f77cc09332a04d8de720f3cd86c6bc3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e051717cbb681b6cac1fdd3298f2f9e522e2d78fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13758be111a39a9b9569acfdd24e535617d5939e81a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc30c0b66890c84d6bd6a6776b9463351da5041394;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c60b3bc919fc789cbcd07ed4d7f326fd15c4c238f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4725beb00c58f4287a39d8840cd26b508f1df4086;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ce4f89a05d06e4eed9957b9400478525547caf355;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10929601b169df75a5e0835edb5077338957c16fc24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f637d96496e0a972d4effb23e467bfc7fe954b57c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16fd1dd3eb4b17b3b6d66a4959bbc38d18267e8e789;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5eabbc0640bfade3617f6ce292c3d1dc3768bc0f13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1c577b5abe4c410c87de13186f761439be901e7bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d965dba7f31d15408144d625dcf21c124a93ef869;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad8d1854425f2c4e98ea112912b548777c7ef7f77a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9eb01c755fb2b52fd11c937b9a5bf41d7d9087b95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ea97469ff8ec97462c203f9fccd1962f235c1063;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fe08d6a80eb0ad2bbd3d33abce066d669b4cb0eba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h25b009bf49ce39da2b513995148edc13219ba62772;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he98b47911a077e2a07cf240126eef9112c1f5274da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118293ccdf49721917395bc1ccd9829e87dbf7f9967;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f5848513f2805cef1d9bfffdda5c65ef093599d4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h136dcd15e0e40fe396300147594f788293688feb19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb00ce07f874add2204b039dae30609e19992cae4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha48aaf4be71b0717f93b82d23de1ffe54d19420513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66136449e53efaf9cd0578f19fb7e997e4c7f2d514;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c4c455937c378dfcdd612ad9cc613ca2bbd1087f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6802b9fe21b151e7740a8832c7577dc1f309fe75bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82edd857e4ac3b505dce87951f17ec1ffd6f42e031;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a75b998b1375f0a1b2876f70f970065996d8be8ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf40736cdab096f25e8156596f123a863163ad191e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101fbc58195c1d8cddc79f6bee36e0549f0a700590a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1001236115adef8ff4e14bcf0e03f49b6ebdc141821;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b44d0b245b8fb6227d916ac4548559b0106df3fe8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1579852699b59dbdeaa55d0b5b9f55ff3671c52175a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac5d1f16a91449b3ce4d55cd23ba27b727e77077b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec91f2519429acabdcccedd818bcd2308984319db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a93ac9edbb721f8612ffb03664f089f9512e80e83d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3da1e3ce7af806cfa2512bdcc506a14206a920bc67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h319d3c51d47fdd577cbdd6d49a8e9a19b84cecc646;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb309126fc6da503d4307b8be1687f6c807a957a7c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2984295eca71c37107bb19d037720b4105b1dc25c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf02fad58cee8c94dc972427c6a2d525b4ec13f94a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1467c53a1d3863f30486ad34408c0bc2fe52fe47059;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51706d3dc16afb87cc7822b9fe06ea29f90a47d5a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2dc0280aec3832057939f614d07dc55d06c13c457;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108793ec6e15a25ae0f761139beabb88a890f122455;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c307feab160add463e98db3e7011bc28c42b84ee7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19090dc922db7d5b9fd6a3ca4ed48e89fb0956d2579;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17eed0638dc7665a4fdd54a5a89ba819be7766e9a09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1029d89bc84d92fa8cee159fd24a378eb8755dcfc5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f392794dfdaa93ed5dc7c4a62906dd925e8b4b98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8a28ee85e69ff9e080a372479f4ce7fff0da47f53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1146a1d71b84f5411129cb8cfa25ded834dfbb8dc29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c9837c9107d7ffbac42ea3abc0d9ac3122c499c3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a57ad0966ed0bc8b56aa0333301a070fb2da25f40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6d94a9d424963d4bee8e46c9d274cbf1b5e1538ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f344d7f4c4f458c485a3a05780360fda36fcaf0ba2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h355ad501cfe20340c943fff4e71dac1677d715d042;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h829764131e5874f7f146f61972aaa40e8d0c4ad345;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ee1b95191198f9f98f45d8c29d2498fc51de0b1c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4674eefcd3cce9584beb38b16bb009c4bc27690bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a21dabbf28636c4984f1ea838213c7cb6c8b2f557e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf48ac9be6b6b4bae2989fb6a66d5fd845cb40334a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ec0f7f3d1bebf20d0de33903a97de7e79feca46a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hddc6495af0ad635da211442f6198b92e0703db17f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12989886e7a49f209a73900ca4da24b447f351e8b81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13365943760cf4a457afe0946e5bbd179655aaa956f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13032437e78e872b4732bc1b49a0f93c1e5379402df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8de03144576f2c3e112eed7811cc0af1257562758;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11c4119aadc77af964cc4a13224ea573ec4b93e11f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1e50aaf16a729fafc98a56c1c582ff863e217588c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e72321b7c437159791aa390d62d7c6a07bdbe17382;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197e1beedeef90a66634eadcd4a136478b05049ebb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b995dcf4ec6071194a82f5ccb270ab8949e060a915;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h750cfa936d9579608d51ca450d22f319bd937e05b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f20ae112253c862262999ea221b8e773d31a6c608;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc95c0d3c4153b08ef8e8a03d2abcf7c6f8ddb2278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e9d2a659685c86318d8d72f45de7f29a5c8e6cd40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5045318f876254e9b8d5e2f67c9407ff1cf4f93f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h630522b0773a449e1210683c2e927c8b8dd1126a4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184835f31357e99200f647483b55b22fe6154522990;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132d1cca4a54bff8745c5083718a1540fe4c5ca7f65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d758ff05502fe483a768bebee1c5517df16cf6be2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haeb1be4894a534b91370213d3d7ce9c024a6e152f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160fb803283fe79d6bfab12dad44d82f22651fafcbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10578dfe3d2db3078a99ba18b02e2bbd71ba30ce484;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169f55f4d9a8580f0875383ee9672539ce864ea8fcb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185abd475193953a4e958d38540dba85a195b9dbc2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h657221d970869b7c1802da7327ab0add0302e2ddc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda95be578bdb81f043e0e3f47b732f123bc33c035b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7782290edfd5758855cbcba2afc9ccba68e9f2c237;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4a1e235a61dfbdd02479b384ae31d3466e2e2dcf7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4290975b083edd0cff61d9c51c5606fd9d671e06b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e13c8f8137f6344b9bb86268c9c62fbc679fe7a5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b42992a72de2dbf6f18b2fce1aa9ac60122241f35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15749647216d5f750b38151ecee78cb589b6d67da47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c39c624e069a7c639f4f59013f1e5ad33f30e4b9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h789272e459e2254f069a4cbb164ff7c6df01f4e8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3610507d414260a2f55ac0e1a9f4623c214167be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150878a07a41fef2ed0c101630fd552872d3508c983;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15546eb457dec0583c6141bb2a39b093b1a49a57887;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed776a9fdc5a7d2db29bbf4d748d520a74d8d11518;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf9a0a3cd084eaefba615c31604046d910e4c8a3c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3ee1ba635ffe7e6b3941b7fe3e512d8f4099dd914;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a7385e91ffff9882cbdbe9d2dedfa7772d8f1c483;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf9e535ac9c6eb65586fda64a33f0725a843036fd1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54da49d440a17da1d54e9be177c42c7721c78cc9ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb05f34a2014111fd42d5959c4eba8100bb00049443;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3a6e816aec71b9ee11bbbdefff91bd197e808a16c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b8f42446f93a55e3788f95fe94467c53bbd80dd50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8fc73a47568844f5d3f8411f45e5e660c86ba5723b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a4eb54857a74e6190e836978373c2fddb7fa96dcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2438c84e27543ffb77d605174c8b6479b08a0e596e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1514d98996909aa70abc41f53bcea9a6658ee5f2897;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfda17645e9a50c98e4fc9c8c9d302c4ee928d71d04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc034a7f97ddb10daeaaa2ad84f79bf7246cf547;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h104eb18cecce79e7ef479bba37e37937b4b2034cd05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd6787cfcd074d9b25eb6a8a61db914806737de054;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae94753ed449dce00a711da503d8db7fec9ea8a3f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10070ae1b0bb7d1f6a739fa4a21b012203da765d71a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15336879c3c9ea08a01c771fb03114913ae61268e24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ca3bbf9fde43552d6b7bbb1d2c3f2a2edd849ee4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b38ac7f5f5d6d2c99dd6becaf32a58b27696f91bde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6666638289183b0230ce9f991919c1816b5709f358;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2fff2b505b9081f29609aed2130a056cda7379759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14834ff73e32cbda73e850918051ff85b7d718b4528;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8dbdaa144718ade20ef58d4b64bae46b76b5a7d587;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb6e1d86eda9c8146b9d80ad636995ab27d27b8e9ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134795f9737d9d8fdda2693416de24b603d121efac0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161b68db40b2ec681485e0e2c66e197772c5d26a9c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1627191c9acb04782f8671ca5e170991b90ed750d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1684056455baccd4b99da7135edc224185c18f633c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56490052e83eb522c6d81d57866836d4bf59b5e439;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5013106bf6cabbd73bcbc658b991ce582967057e42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64934cb7529a6b4c832d57e45c552c66ea9fc26807;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62121a33b0ba1c6e0aefd8b46032d6cdf5fcb798b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110d008356aee69041fe900262fd8d91d92a6afcffd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b982b2c54ec6765b272f3d217ff89a635a51053e97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192e0605b2e89acc6bcee9abf9ebac62ec7bb84bca9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc11590289da6e70c812155b3b13c28ca46caeb5a43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba364dd815e206d5737031809687d8dedb0f5a1c5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95cad22de90ec4769f4742737d2ce6090ba5572431;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e3371b8a351d3c86db6af5be928815899e59a47ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f128d9a3a64fa2c095e79e39e55e14210c2faecfc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69fe349fdb11c68ef431bf70725523a1ea51acc026;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bccabef5d58fd9b0b12ba813bd45d8de1e58edf92e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ae9890402012b57010693a35ab273d33c0a10e8f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb696baf7aa71ff93b08c04e2efcbb97e6c3cb5d4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b733afc804e6f866143c95c298b973b9066684514;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f19ee2962a521c79160601cd09ea985dc068d30312;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a92456d910be3ac18fd9456aeb923177ea7826efb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h834c2c901990e18f646fd2e78d0d978eb95a92dda7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f0e8e11ded834026b99a57e9b15b3e02f9a54ef72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40645894eefdcd62088c7bb8045128c5620705257c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bebf38cf9654a4b27b9db8d4f4c6bd66a8470e6b1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73f74e8cd43b1c855132eb5bbdff8dd70dfd2434c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158c997216ca102925342b08d022b70a44d1ce6850e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b3ed4f39865d7670faab9edd638929d8ca8cc1812;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1628ca7668295726c42c430a665e3bee606322857f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c54cde5796bf3c11711b21cd654677df8d0a062a0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a14bee1422a4f0540d268c43a4f281fc08f4333bc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b74e9ab72f5b13bea038f2907aebbd4272c730a0a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b97911387ea91cfd0922b72837f5cd3dd437a3b1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4b91f8e3041340093409bed87771573558e9fa248;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fb8a7219ac46a2c5857fd75bc6a090394fbb735bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e80ea8ab156d1324b831f75d689104eef7962c2928;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9d6943fe5fbb94dee3c6bfee664ee396e4706e3b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15cd74103dad35b749ba3d5bd2611c7e140d57e358;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119784e952adf55e90a4016b0a67a83b0c2f2b61e29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccbe90e02ddf1f7a71a331f015465be2b1f579c734;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d1627b7c0ff059fbfe112dec6309c35de5f72b92a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17060127fd0834447d541b0f88e237c36cb4cb83984;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3dcda3a3dd7287eb737c70df33c4041b524fe8134;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd135374ec7207f1bde499dbea80194ea3229e1993b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13056d4063c00e43b3afe6a3fc5bc6b274670b86609;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6bc8f08c6e99166e12218d02575ba337fa68e4e7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d62184454e2039a9c45e9584b24bd63b3f1aadbd1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf5d8f94e901e6c9b561159aeb7983c2e6a182827b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1878ed40d4ffad15e2903afa70e0fd5a5e09b4c10ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a784a0d4132f037df84d3ed86055cabd508e49b61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2939b84184e1b0f7713f1431e043baf0bb23976757;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf862dd99970ffabd1eb2765c05190b7099279f41f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h583ce381ea25ff648e470d5fc8327a766f2387c064;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha32fed4d76b9ab796d5e7dd45f6b264d7d11c134fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c410906014e92000434e60884094eefaad39cee966;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha242a678e41e8e49d6314ceca468df004b5285a392;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b338d9aed136326c2deb032d2f62af406b62a14c9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2f7912f226b325df9362f096ef36ab696056dce12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c38723c28c6bba68a16162a65f7145314ec62d6a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18752d5b10e9256c8b871dba9e90b12435438bc3ca8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb32c1573a30afe94855986c4b4e32e89c76361a710;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b58eb0a18380f84270e1f120fba5406abdf96c37d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21f0f1aea1034ec501e09db21cd984e16cdd74f768;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163bec3f1cb5c2163942a49432db6a9ddf7bba0037a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9b645df0f2e578c9cbd3aa92ce2bad1937d68fd5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f19491e9bccb1d3abc419399b8fece1ceb257abb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153d73caa59c12374623a0001c814b5fcdb87e824ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h931d64ff39b9e87dc94139fc10b2b6c95180366577;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a4c65e322ed3503c726e665fbdb1749271b78d6f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125f7ad6fc633c8869d85a00a26a5b050f60242afb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb6a8f539f069f26e852f7eb093449065e06cdc1dbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9e3e868d5d55e8ebf993586ecf88eba714824fac1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b499881324db9c1394250d49eca31a1644257931d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cff645911ba8d8d975975b38e5de8894b86fe8369;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aca9049ac0cd63cd88e4ea196e3f194b85224c52dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9409f08e3ea1b52bca8962964904eda29a192c9f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b80c4bec2c8ce474a8d3a7061bd79ab25595776e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he129b4b58200d9a26389de36bf6a52f2a7000835cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h729b2b47bcb33f264e350daa19ba53e5f69124d487;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a887395cae0652a5d4029f3aaec1d9e5dc72ff14bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ea4e6dc3e2067e4d735a0d440558c13e00e66f6e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba5c26dd4c85ec370b003212d3994eac9e4821aa32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153779c0236614b8aa8908eeb9349e814636ed1c23f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf174b987da14f8e5ca28b8739fa75a3326e877d77a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8730f81ca597415d7a1429cd3c352d77dc2c0d7ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc0bfa4a06a29970b74e66a0f4a99e35db2ace84f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e8d9b18e001c0e35384c5c2272989ff0bb5958725;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fea9ebc2e303573dc93c1661c93986878528cb78cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18661494bf9d751f0dc3f179a14e25afc561b42aff6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha821f2aeb4a828f12b22eaaddbd9f549331ea8077e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1654c1b7c5b198952d42e26013117b1c62b1ccfeb47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cbe590c7f447a80639b7b0fe8de6be598fb39dac4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73314d14ce85d76494d7989ccf7bf372d3e80952e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he52f24910f118f4a5615a19bff94bc8fc9e3ce8afa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1973b0f7c9ef0fdf093b16a6743bc96e5bdf111594e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb08a5d340fa1dfdadb236ebcd8cad6c48f2001756;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14bbe1d5ead3875bcba0bc51ba22a65853136190ab4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb111cf8ca5bea64a2ed2fd3f73ff5c24590bf0c386;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1878a92ea4eb9a4ce786ed1ce04cc94dd7cf83e55f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e8d3fe4081bcddf08882a71b640d556d384f2054e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccd1e1ade97e3e4c58e7a9e8d10c17e0f75a699f44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haffbbc64391d6155ee308a9ac3332a8efdbee1aea5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac73d27a403086e817325b664c587f15064eda8bf5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1275eed85c66469fe306baaacd2d0fcbc2d7c5496;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5daf4c08dcaec1c71b07b41b4ae09164071d46fae9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103351d4c2f77c8d33216d5a393a5af14388a9b1856;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152a1bb8084794d51178d81d39a44aac738d522264e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfbb1dcb6f029d2f83197fc97bb83335a86023967f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f89a25547c15b3b086d7f7c643b7399fc64df7d88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1623f6bf6e73c68a188136e6bb3e71f296f7364cf9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d40ee6a688806809c8defec691d608e7913499e27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dd8fee916c7b7929a8dda4add465e74cd879cbdb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8274788e8e20c720616cb92719d91227da075d7ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb63658cd625967e1088fe574e7ab3224ecdb64703a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d45e45212fb1836e93a4dd796ef367211c45916d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f63cc891bbf720d6b3be304f0125067652624f057c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0aa58804ba0a2e9d395f4dc3eb487e727b44a5f78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf7898a2ceade20cf7468d401246e78c4018ae3d06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a9308993725a638db71d61bdd923397c93225924a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119eb7f0521bdea266d5fe36f9552aa966d53840de6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d4f1a9de040dddd18c804417638cdea1d17d48eaf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142dfb01f94f8245f8429e2d4bcf44e80636e1b56fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d8fd54317b2c57741778e5d0c3cb8180e4a722914;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b57541581c9814f552bc632b0f8ec9c0247c680b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hade0ce1a2f79883c074d37c621dfbab932f0b61006;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93e5937b8f956b21a390f0371865f771302f9cda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcdc1855d093139eefe295dd8934c17fce8a72775e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a48b7f7d39ae9ec9c0fb91bc533a5fbc34f2ee119;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c514d506feae2b4637b636e8622d2d8ecc886be75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h548946356c1858b66d0c908cd81c9156465c756295;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecf2167d37539446fa84ab0c977fd79c9e9f8ba786;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1454ce2ce32898f9104c734e26ce5ede6188d665777;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169c649982a1c2cb11c07d69c4b9a8533beac18ee5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a5ea7461c24aa287ce13f81dd03ece5807ad1e210;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffed97ed814752252904e17592b2942ab7cbb573c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18138793a6229a1f785901ecaac5bfd5c822aa79b9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfecf2620da8294176d909bf2ee894fe7ca7f311442;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa994da075e0aeb5d7e65128245ef2f590baf53eb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd45b007c1b75d13ea7236ee6d91202c11739228ed0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f85e39675c2541d3adde7bc4f4582d0a42a391abe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22683e9bd93e251a8a91c537e39c4259373b592759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177bdf6d6cda0c7a025c1465280081f1563706ac919;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc9da3690e2d9a71253494ad27bf48641fe8be6799;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d64ab91d9188fea1c40c786ae58a7afdcd7b68b7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1713668ac747aeec6d6d3c850a52ac1f95478f9d9d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ba6b671f0757a591e806708eacb54539598fa8810;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6226ab84f55cdf4b9674e0e10c6ea2a5310980e335;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd24733f52c759c0406d25d1b48a04c74438e03f90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ba699337e2c15c62c8c41d02c05eb1db436b93df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dabeec77715f175c11eca203ea6edf3ed8614b2e82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da367886236d99e9cfd87fc41d852377e806cbf962;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7d894b3049fc804cdfd53012ceae29e0d894eb57b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e963c2148fbf513c6dd1d8e62a78dfae6782ceb5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd04718b39c62fd88fc53eee2374940be0cde170eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h67d70ba35c1c4e65e3a832f4062147c86d33a7648c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfac5921145f6253f7f0a896ad985fe449b3db75b90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd99f2697d8b090c92dd2b819e2a7d71efc29ddcdc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cdf486cf0548eaf7d8c398034aa91dce0944975425;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1234ff3166e0b21fd2e9029e5602b88cd9efde69569;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b0d6cfc607b818ed99a08c1108dc74a0270990cdb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e56165c838b86839fdb2de18297faa2baf95634de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf08d8a8eee1781ed4d3b85dbd7c421807712f5119a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d1c98a240e1358840d5bf7b4fe455a0568026b7ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h603553b5bbf473803b893a0cda6963173dd7bf5796;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd48c382eb5fa98ba5b2ffc1bb1a666a26308499acb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a224760e019b2768009f9e3be3732ff286af74dc42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8265072a9a54558d5f80528aa5db32c5b58bd62be9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1dca966ac82e89bc24b38dcd89cb8da1c7e3f98d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b583022a65fbfe93aaabf4dfb2b80fc4a53bf0a19e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a00c5c6a9e218002325c0eba5565aca99d5de9eac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea2b924005a2c0896b08b395ffcd607468e26cbc68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1330c3a188ab62f356bb3a05b01319d5bed7cc6ad57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149f357e7467ab6f5bae9700e425129ba1b3ee59c6d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h690bcf5c68f8652646f3f5c9c20a8727841128255b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cbc47934f2bcc4ca6f7aab852c8f3bedf0d03f418;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf1a315ac3b9f4e865916833392279001fda0650c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc321e609c6634d59d36c75e4bebfea057f6df6d9a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c44f615a818271a2f438c81cdb27fbfca1f8f62a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135a29280f95a51d386995f77b7927d470c1e81b34d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131bac41cb7838e0e222c33b915d169865ad2fda13d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b81f486aac694f052d255915a2c1be5f82baece3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86795bad0e43b27d034c4e2864c26b1c85e66bf5b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef45458ce34c3550b18426ec21041c4f31b6d60bb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1006ffa5bd75d783ee4d3aab5218109046db52d468;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h221e13dd78a221be6107abbba8411121036b5a8bde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1760ad59ef1322b0b4ed19e6608cbe91cac7725c558;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f810c00addb23562600ba639ff67ea89aacf44502;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10caaec0b49374cc1407d46679fe988e63e8ff7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1849d23a1da3c84991d7bb92aaf2eb7621624335582;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6fba74fa24fecfcc4c966da2725bd44699b9dc23c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135684450404110d1e7788bf4f0fed04fb44c54cb93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156e7f34372ff947616787374034ceace0fe9fb20c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182d8f770d21407c148f17eecb67864cedf0b7601d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c3801d99d3c23acce867c91fc44009747fe52c384;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d83b925dd851a3b21ca867b0a97208c9068bd31fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a42d8d1236ab972e0444aa54bdae8a959c59ba12c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175cd93b58106f1018b7f67d4267d09572f93238692;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1065412aaec587d8e407bacb9cb9ea2e360646892;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178a83bff62db77f7a8de1eb4b506904a2d4abc52fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d50dfe0642e238b64f8ec50e5f2c3d606a7681a741;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcfb8d0427e9247723c12d204b25081d100baf024a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147bac75e5f4b0359c802ff36220a7615b942a7897a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c699883df89d99b9effb389f3d6ccca60c194c8347;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91b766e6927332d7fb9e56abb0082408999152d3a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1faf0bcedd8f0e9e34daf923755289deaaa351d1211;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d3a014a2d9b0871c4150691cbdcb0d6f1b0f5f969;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56d6f9fd7d6d4287be1d0fb238f8f5c245571419a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9b294de8bb9cc5a39d434b64bce67318fcf3c0fa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa3430ca74bba8f632fb0da9017a14cf740ff09244;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e026aeec6fa3bc6abf8088a0f15f7ac5a7736c89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103e86fa53cc91ad626111ca2636fd34cb14cbc88c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141d189411eae2848a7aa0866e64a224faaad8e79a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ec67b469d5b061e836341bbcec3c9df947fb9541a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138e617983ea9550e6c5b92146d964c27bbe6c525db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8d330c1dcb031a4649f076d1f570f1866dc623338;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70de0b17cbc210050c047ea00e3b00b43ff3b7075b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbbac420b242970ca5ad69cbddf906d43192f2e5fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4b4302e3d186278631b6a2b0e503cbafeca88cca3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19853847c868b99eaf6d37066b8076a752cc89f89f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3142e19f85150ee65336cd220036d7f002f27e97ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7fe5ac43e6ad2a5bf71e42fa189d300e5116eb2692;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e76da99fa88733517fffad05189cc8688b1068c49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefb335349e9c012fac47363819580101d67c592348;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d8fe7c222082ce30af14cd18e33c0c20b4e8f3e6d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57ff177e14409ccc991f6acbaaf268c9c5555a1d32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd887ac0d7741b698a4255058dfb4c731adc58a6efc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3116c0c37584ab25cacb73391b90fb66c98ae580f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h808bb40f778c134513a229b2b7a4d0917ad73ab75f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d87b7851ed9a1cd1c0335f3659ee55ea834fc940a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1045bdd6e49d63d24318eb76534dc6b6b4593a9211f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15abda7295044c8fa893fe6a6f3439ad1e48671f757;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161e4185f1cbe56da367ef19a7cc64fb5a4461b9ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de37c155901d06024625b493d48c7cd23165959508;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176139292a8265762a3e867c26a9baa2f3ede9d1662;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5719569c98f7894f56910d8ce338adce088c4a2591;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b4152a61e9bf58af3dbcd754d55871bc9e36a026d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d22161c3c56b630c3f829655667a74bdf6f412a5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f2f5e379c0b459f83e118c33557b7785e4d3aecaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11077bcf7136b79c6cdc159698693f3cc96a08f0479;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a5c75acbe88f792aa089ade60380f576ebf2662e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14395a3cdfc66a0cd7f3d7213b81a0510dfce8ecd24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18684ca014079b16ade1e024b7b7da44b69e20d20a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b48904d18346286c06d317f3020ffdd11aa2c5442;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197f16fa736afff72fdab055ddd971c96ff26202864;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7c8370896d00082cc901475107ca98fac49f69bd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c01b9dfb746b114d3ee07fc3b227248f7861b041a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18455fb28958380a4f74b31f2fed72d5f46286bb726;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab1a176a99197961ccb0768f7eb40f90c21a74c751;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1971dbc4aede6f26fc200b30ec4c652573fbd422e88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1536d4fe3356dff51df896a541c21efe20efb3fd78b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4ec81e44ffc287c00099adf5f3b9c5008a2714231;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1deeb190785cd77c4ec4ea4fb1643e9d3436f8529;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4357f60f06b6af08b03ec743118547caef06d78372;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9abe46ef458e97f2aa466663bd9b72d65f3247640e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3551c7c60bc360af7a649df5ea08cdd49c24f898a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12cf102164590d4b7c7cbf1c06e25e2e50b393f8e16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1564462bf7e8bed0a066d1029aeb393fd1886c66d79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecba2f9f0376c5baba9126ecdf569053850458c9b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d4941608be6d48409a0c185af1055b4219d92dd0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17aa01e295506c00437d4aa9ae66ddbefb53e681c30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5aefb03f2bb7a040ea30ffc8b6656fa5ec5d7f857;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77ad4f855fc97ebcc7677bee7b726a178de65891fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9425326529991caab6755e696ef659d689fb26743;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea91f0c2f00d9faecd235d60002772468d74ab4d09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19baebc9ae4171750a2aff954a9067aa74cb39cddbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b606d66042d3a9566f51e6b24eedd6d790357b9bc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd23a1809a65abec82f392c04afa5f59ce523cb57db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb81fd2faf6aa6f43a899118d52f2f7cfb5f4ee24b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111e3204a21b02e33bb936414af7f5b129eef19daa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d94fe8638503fad7c7cf38bd838b5bd51cf499d5a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51a098aea0f0341933ec287704538e41e8fc56f39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7ab975a134e27eecc662db10f0c4fa5c8ef1b6320;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92dadf07d5d822d24fcffef71c0f60cd33e602e4b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1728a4361b2356c76ffe50600d1f209da2e8959039;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e991297874eb4d1100eafea5706141bd60bf0953a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94163993787eda40a303e88df4fc7d317375b2084f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h96529b5b60466caad3289b40a46292e378686998bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e3218cda1660fa5a164aa5a65a09a4cbd98119b6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcccd9c335d1fffa60c1f6a2fea0263b867324e9f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h46fe8852eb3578855a14c388f56cd55eaa3d38addc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h570c39ec9fb58f23141fe43e5279334a94419fe097;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ec2cbad01c9eb75d81c302e4a6ae4c654aedbf6ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce3fd9fbf181c732552c9ee552a35e3a38f9237e76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h745913a76d305d8e1214d1d13e74bedf346731c119;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf60e3aeeba4107b9bfdc29313cf4e7d39f90edda1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d82896fb9ab0d8be11a8330d931307024ad1c459a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142afc44f9d3a52d3daeb1369419b1450c423b3aadc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6f8d19a98652d6c8e7294cb2baf880556781a4937;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a4f57a59024334097e7a421f408dd5d617c222a1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h859124b85f8f4e745a87bfd441ef88e4aa33092c1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45d9055a60da655a6d27070c575a3b5e6374d40286;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89076d2f15e8b716fd87599d8072b14878fbee85b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb25f713ce222f39a4e98ad74371ccc8a14c63c4b35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1793b4afc74d8136230183716183485c0ebda44bee4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb68280a9221d53dabc6b9d07f5914fff1aeec17e4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a2044eed935046d38f1a9a5335bbb2700c229abd9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140c8907f198e545f9b4a4dec7bbd5b2d61b707dd07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1846286e60458260ede2e24f43b59cabac94d585dcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94c55f9251240de0e3f40637137462f2a60c42bf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h750265df98b5aaa34486aac3dcb27bebbb9e9166e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1626f08c9bf48937816b1263d45cf036ad6f0bbeafb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197e45dfcb0c378cd6432762fdc1e44d4768e322f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8c7f8f11bcedc6831b0c1d910a1dcfda8b4de9095;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106e12535c432a084a627b3a2647d31c25680187c86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e16def363e7e66171e19c5f796e6d2c0681c28f49f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85499c6d9d7e94690ffcab7103a56e26d903c0526e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17c4a166d9866fb50f32a8fa434e4b462b17d64eabf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29db25a096ee4c07c66ff1d1243bbbe774a8118a31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99e1d2662b5de31d9386c1b5e0d07ddda832d472c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d9bbd9a008b0db6a776ac3ca264bddfb392227a3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcaa2f2944ca753e113aed9f80292e53b24610e7ec2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0823aa4ee3c532d422e9c90765074b612a2c3e10f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a9a2a01e54817403219873aab46a8693926903c01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f65e017662f3f084694f33bd12008e8929e23ecda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haec8f5469f13874ef754f0c8137816b26325b097a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c6696fc01b31f130532ab3792b6dfbd36202ca9dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134175cfe914d9f8b894df1c3b9a5fa8cc043e3e513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147749150bed8cb860c6db37caa5b1ea9ae5a960aa5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b7d8148d6610c1f3481f59873ad3df8cc3136bd75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126574f51e86020e65b5307f05df1ff63cadd344fca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175f8ddf75120d15b145ed80a1208fac7ff5746034f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha55bc8c22149210418810d2c1040c750271acc7190;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h362afc4dba6e9556055b57fee3badd2bcee70ec34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14546d388cb39e8f431f26644d329786b5b5b80fddd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1882e8b41143b75a7d3e87e63d36860546c3f268496;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172352eb7098daecccccb657ce5207be9e0dd6ec645;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab45ced9491d662e1fa5480d1c06d979a4d945bf79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1515f784bf4aa8de516cdea8cb769c1425498e9f41e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ed025356458868ee09e17dee6f0db7836e601d220b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8bb7dd566d96d749f34091d57e0a16a700e42fb30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f2be027de069907df2c46e2163f58046dfc1dea3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168758a471e49a7eec5a7ea2e96d96740e96771a4b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb86a54cbd04453d94ade103c8d820c9104c2701f8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd39a0e1c2f3e6387004f23aea689a2049c510acf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc43bb99ed4c09fc4b7290991bd2b6146a5372f084;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9fc9fd8b654a49af4ffadf5a14acf62a7e5ae3c86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e411c73683c81e5f15b054ee222a5bb4826922282;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b25f2a266103be7471c8704c53e0e0752afc40511;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8554c3fb5a540b3ec6090c928ac226b421c5f6f5eb;
        #1
        $finish();
    end
endmodule
