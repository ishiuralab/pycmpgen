module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [12:0] src14;
    reg [11:0] src15;
    reg [10:0] src16;
    reg [9:0] src17;
    reg [8:0] src18;
    reg [7:0] src19;
    reg [6:0] src20;
    reg [5:0] src21;
    reg [4:0] src22;
    reg [3:0] src23;
    reg [2:0] src24;
    reg [1:0] src25;
    reg [0:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3])<<23) + ((src24[0] + src24[1] + src24[2])<<24) + ((src25[0] + src25[1])<<25) + ((src26[0])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24edfee5deb4668d9bd1188f662633e3a8367caae2539bb11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c342446f015767c47e8ac1ce0f29b7f09d368f641a2d72a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80a59e5650e7756230a8b6d5e552ba26a67bd3db748680ff6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h511cfb4a6a66a1114f8b0f4d71f89371b00e047babef4c8dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f11cb0af14bd18875b6b0cba0d87026a295ccdea0b1b2eeb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4b96f6d418a2eb12c8d248c2070aac45744f3245c29d3ef3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33d15e30d6fa5fed20b8c92b9fa3378849455d81d5e4e2b1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82caab604a6286086c51dedd0f5cfe9d352e1a651cd48bd82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8e1d97a4aee4248257759bdfc9eb59176d4b5ce65934fdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha60f913d52cd9ac4fdddf4b3251682b847c212dd0f684c857;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb07ba8aaa91f3f99b981e9a51b1ac7c003e930d635b9303ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h912eb45fa98bcd017e3a7c73e5f3e42067ea2f32c57d38fb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2199078d9c4c4bd51d881dd2e43798a0316a23b36657a356d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc99b07e9fdcf2944be5bcd560d6d88e202d06cd7281ab9e5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h620253164e48523930af90685f352993fce1410e21b7ff2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca93af95aa02631888c1972b81c2b87f4ab5ffb48d335dc65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd146fb16c66a81a5f4568e25b1c3583ffa201fb853e593e45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h198d672bf5a5cfe43296ddaa9d85b8a80e870e1b22fa9ef77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h934f5236b70569ee278a86b977bcf04ad8038bb7989521c31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a86854d6b64f1cddd17f1820a03875cfe3439460f89ec780;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99eed77183f7fcc2b41b04f1fafe54912a089fdc978c99b76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67fde513e1b44f3da96423c9dc8a2edc62be003c068069228;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf6ae3b9a0f3862029027ff14f0a53da812a18bb5a9a914ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8841ec17717f1fa5b589d4e66eabdfe605c966ed3088eb38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafaa5830f3e80b9dbd561f1cd4b288816f7f79ac7d903e780;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9552c543e276cbefd96417498d02dc8220056acd0d1a01a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc58e22939d750a25bdb3fc1affb21708bf9616511fd18f55f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a3417f841e3d29ee2bd5b55d6b4689f465f2a8d97b484635;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f08585ca6f6e43b04df920dcc771a198e92f8a69076a8ae1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe703cddd5653cd589fdd07245031487518b55d66cc8ca95d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefb31b235ef5702c66f14ed7824ce77d81807da2f96246abe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c334ac5499c2229d0a83f66181e6dfe57d84bd4f28a6141f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfac10dfc5c67406660e20f79483bd356520953819b86cb1eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8604a77b0b119c7215cf3446d5ea0800250ea7f9e238b7b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h202562c4ebcddf512a71221abcf7d10d6f1f93a53b3b6447d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec8ef7b90a9c5b7129cbbaf6f9559a2f94a86f725fd7621f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5b4784beda9179bc5b50d51efc9e9fff3235819c82fedb5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a93a3378d5caf07fa16b3b81c5c0e231a2be199702ec8083;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4830c87df0c834a503e1408b54db0647137c236e655cb23af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c8058610bb6785a43c6071c0d4fd76281455c469ff59d25a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4096795c3abec13990b451f182c8441ec190a942cb49ca2ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d72f65739c2b7f34ab496f078ca17608dda02a278b964d20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2970ed292b0acaf9f5fe05d95a33719ee72ecfe938ef1e2ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24a0840773bc61a6f19e49d9d3a1327b66aa38ec4fd3ab14c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93fd7677cbaa779aa62748de914843e2f2ee36462a0681ace;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5480997ee085267654b4cc61b32a81e01cceb39ef1fcf9c5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcecf8399888e837846e255e843885175ec2095e78d789777b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69204259a35a0fe993625bce697edd68789a836f988ec08e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h254c56f2cef4c01ff8c21e7d1c7ce08c0d6e47c980312169b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf91aab8c8b16639a78f44cc71251c78ef5880c8d603894dfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h526ceb0383fcb97fd941437fb7555598ac525b2dc454e258e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd7212762179483ee7693037e45ee7b560d61fc0da386de38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h872e909e68b8d9c64d28941f5c64c43fcdbe8788e9a07caa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f68750fe58d3ca6306f5caa710ead336eb6c0ea6eaf5a31c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9b350aaa3feea7951518bcd3e19d5fb44d8ae43d6968055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d1bd9b524786aff4dd29ef475a4dcce0a227fc35c58359d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde85479dde200dab66f07a4bf1e356eea390539bd4e6c2922;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83c734a60a863766d02b19bf22114c9ef74c8863741602803;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66d7118ca5406530663fc6a9361e193859ddc44c5038f8318;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d9ce2a2640373da65579030db52b461ea7634b561463e2bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11e466bcc10c9ebf541b99e59b11e06bb7b6f778e0acffc82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65a1c7a20263bfb8e481703e51344efd2b71d1a1eb0800fba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb74ee747d219733fe0784d3ec731ea21172eee7aef25097df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca307f707d85621c00390581c3a6939bab08b95f14f226436;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h963f7c5f881a57d3470dd2cf0e438f7dfe55e2485b24bc032;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdef234af813f16b3a48f8d02381bb7f1dd805e236b117003;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf45cce9b278638c087742743025e36e5ac22fdfe89f07a2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bf690dd1699bc4fe9032e346214f7bd81c55476615a8a2dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bd506dd474f74ecb736ff16fea632a942f76491c863a8897;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5967e7c9ad2b508647ec1bd3c258ec6d0d5cad4a8129d77f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71d67befd09d37a128e027d14beec97322c9cd8a2110a9ce0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h654ead4da75bc9d3a27111bbb6d18e7ee64206143432c7d10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e067849b146e45731d39e58a5310b70fe08e69f5b1516af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd16b7b746ceab4f98107d766f729ab3646358f3e96fcd4a95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a0fa9ebb491d7e22806f4e4d3889be7ad68eb958b36035ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f5b4fd8af42f9d1831c15906eb6589604e63835cc3afa768;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf4f4083b4c83f7d4b1e1ffea1b063677ec35d24029825865;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c9f5919294400ea9d403b8fbc8217d3ffbd80582abbc4a44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4106713f833bbb11a1f354730549be84cdacea2de1ff5e44e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3663980b10f9e9120e770bf2f004ac5a7dd9664c1642b1893;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3f758e859857e45e5b22f43fd7f6fc7ab0dfa0dcf869bcd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f82219ab82c83306e840a23d351e26d9d084c44d9f5ed3a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50e36b8feb25a2233452678e607365ba8d54298853d9e445b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b3b28aef82ed43e24c1b48c2a89803136769e913514351e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17d388a61423f10933c066806e503d4dcb5be1a9dfd437555;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdb203f948f48a377833685feee1b65c06b223b86bd5b11fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15d66c16f4c398e736cacd9ed45451c3d9e6b4151d63f083c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb06ad1f97a8dd15741b45436c2ee7556ff239634875c92015;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd1a31bb768f3939d89e8eb3124b6bb65edd6e980f850c05a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ccc026f92f5e5249ed3826d69dd439c0de85631f0989bff0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbcc3400bd6a5f8a2d219c2c00b92eb4b7dd64f32856d31a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60cda0668269d2ca753791c760f8f326226a255d5ee242249;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd731f0f5d6d34eb80f3c411489f2a1e11316d3e541388b2e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h263e822ab8f2fc14c4c1c5b201b83873a135ffe0add49bc99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65c839af77e3de351fb5148263e2d67ad18cee8fd1de87828;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd65a160e118f0d292975b4de983faa0e71e5515f6d58da6b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc82a66fc1a0682a482849ac46ff8d618ec952e3c3caa0da6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40e057313b46bc6fcea363cd7d5f19ea4c9eaec520cb1ed3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef1b3a58342e2bc13aee4b35533a4411ecd9076b243cba1b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5de17542e3e0cde0f505cdc2293485712dffe33517f82871;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26f671ba973177971fb759c6ee84f9f1c1f4d84cc61d60cb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cde0c29f490fcae0ccc53a87fae814a26cfe314f96390eeb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdc78c12095333ca6d02b821877c46fa0bc8732def816b8b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac05238ba85424006c05f3ba9d6ef16604e8f09debae5bdb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d05f16cda9a433cbf7740465f82e9d2f26a4fae01ebfc188;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h815733d4e810607b0b208117f36b50ffc6feac845df18f8a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha84ea86a4965bd192f2bbb2d32eaa15cebc7e4e9aef703bb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h480c2cf4b440339cbf7feb564731eed0ab0d3049b50741a35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfee35282c93dbfeecd920f78bc160810e6f0c57b97cadb3d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56ac7e7adcbfe5d12c3cc11756c0f9aa83c778e6351ed4c38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63a1fd06d316da0d648bc726dbdc6646f6d39bec0ae18ad72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha47daa19478739a6b061f75d3444de8386086be89bfbed373;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6570a463ed5ba42d2f10177bcb8f14883bb44fe1cfc50dbad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37497e55cff35a2053a5c4dbf7075571fd18b230a33144617;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ec07e0a08b50ebc410aed898175bb48bc4a7efa79ed6b088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ffb296d5173dbfb9d7d45b46e829a205d509eca57fc591de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8b6952610b41ef237648adb85cc9a007f070ca96ff3dd6be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h254ed1faa1ce266fc53a5f03c79c8fc72c04c570b007c4f40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5d5a1215870ed34478f341f3c54cc89de16a7e177780c72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h378029e0e689c663e264521b78e7a6ea8cd71323c6688e041;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce7bd5b7e26b09d35ad0a9d146eed4a0531569318d788dac1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ed06e309acfb6a6958b0589daa525efb1bf6ec06ff8fd170;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10cc1921f8cfbcdc96f98b92618a118491b6db13d557e86bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha576fcd054f424ca1f7f727aff856278ef90d2c33853a74ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h883d3fca8cfd158338416304caf3b54d9c59dd74282d8eec2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h197d143fef4fb1e324df6f02f179b0ae23a23c3fb5a4f6a69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f303bb92143d278b164ae0ef64b687e4f9e3d34dd8d557e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h286819e57dbcb3b6ad28b8974264dd34a9b324e4b4c47b870;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96cff82f8705880677757e4a970ec64ca0ca8fc8282cd46c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99146183e3c2e62f0ba74e0ec9a81e88cef48075ebb4034d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42b2c37a944c0a154c3e9b17786bd0190bc9bac802ab34284;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c3cad892c37bed3ca7b12565ea4e29e316552585ee75e4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e6ee714f688fba14cbedc3b52f1268ac4b5cad6eed695667;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcae7dc11f8ba2634cdf94a611f665683ac8b53ac7158e647a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb415552a028e180f14849b43e3f90c73eae927eeddb5ab5cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8968ac93385d41cb6b8533879f13a2056b3b90e35a87b3b5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had72991a359b66b0ec2e0eec04eeb562474e7f2e1fc51156c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45f1d906e809de18e34584fd5575721f639ecb4363d28f31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1bc9f5d2548bf60481b86e85ea4dfbcd8c55b031aebba0d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8ffa569b4c916d497d980cd26419a37549c6a59d9451b385;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0fd6eddba54a4f96dd493d907ae19789ead31a7f229ef078;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc668e0abd198b82d87034f73d7b692dc244423b0ce56eb8b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb38824746c6723700318bf761b936e4d5e6e0764a627b1870;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h686c396b4a0da86d4a320058a196cf34901a3d7939bbf6c40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b75e307bfe23ef3136c9003549939dba2649f1bb6b5acc08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c149b2fc93d74092b05ea3e823ed27892fb314e95b34fecd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63f9d76ddb2352100b68dc9e95a4d7443f7170231373dd2e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda4299c439ad62621ba11c7482f7e9b8b99169905ab5ac7da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf957f8b73551043723c36cfe4d82fef54dd317d6fc9a8d0b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd03929a05882b2ea7c9cedff333ca2262f12314c1a95e983c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9beca12e4f5831aa10e4b93060eb421fc86af0f98c3f5936;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he54ca154cca68763fe11886bf96e5abfc8151c53f3510a45c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf10abbdbbe93609352483d590fa9f5721ab098f48cc8b661;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21bf1a438c824faf362b08366b47be47e7db95b6f09004107;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h390fbbf943c93b11086684b6fdcf4a32a840050067aec2c6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h774a4ecc37987983dc5c33e1b2a257b2aa3beaa44fec48188;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38380edc36257d0e34975ae331130bb468475cfd2fc7e6f2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a12d16f49c8b048d691a982ad46fbd7481206e66ec5cc596;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd95f683747e344d67f46a840385a6d6d12f50b8ec47bbe8d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfab329715d66c4b21259c1860db287b403541396771999d1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda8ebef055825c17a279116bfc214ff968c1e5ed1e825d12e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6852454f42079570742c080f5636af72b53118177b492bf60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde2efb21037792ea590c254b848c0bcbf297f4be8be1fdf40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4722cde168d27af585fd8c4b197ef731aa588d37dc6f20563;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3599ab9fe8bf34b97479944a7b0ad9ad7e3d2341dc6f6e0ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefc660d3073ac33088a3ad7491e3ca8d390f16afe3ebe2ca2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9880655084491408fca40d2138d66f317bca079b66426e9e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72dbd54af723acbf9243ac7aee916824e03fb35a9c00b971e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ab05e5032e11f4a33c713b979a7e6e747156967c1d514019;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e3d558f8470980a81ef9baa83a9d924aa92fc46ff71d5430;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93c0369b59aaff202996f56813c4d644193d69013d8567c0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbad34cf476491a5ce116dd6a5a97542b8322705f1e68cb10b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8f3e83051c9483981d21551407c62ea54638f0b93384ad02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb05fabd18f294f97bf597787073fce176719193606d6eba6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0f0f7d54f34b036fbe0263e840704044a5b459db34a485c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbb6188586ac81d70d580b598784e25e2380a4dc54299f12c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dcab5c3f21f3cb3b5225fb6d45500fb27715ec5d52bc6aa6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d609be2600f6c6f9136d9ffa71f2078a7cebe7ee386f756;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5ba3fa0e9726dd8a7191498b168f92608d8445408655701b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc272317647c6b3cd38658ca0631efdeccc49cdb7dbffaa6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fcf1510d55ca1d7e7e3eed1ebb1648d43ccd6f9546b7acb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha94e71aabbdf2004701683bdaf9f6f9b1b0b1292a2b600c6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ad40678e4a33fcfdf96cb58f475d1e6f2469d2fd09ed5dc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h109ef18972eb06806244abe247a8269e109f73ec4b4622fad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fede8dc0563b2c783e20f771b9cec02765170a3c82a2034e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb3451ebc8755a71483aa9dfb428675ba27a74b1277ba96c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h407aa2b1ac19f326a4968c3cd0448fd9e48d90a7a00320c9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfddbc752389712b06c27208b6e0f836665b03a795203fd6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he71a16476e0a0676edb97c2e321ab9201d59ac162febebbb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc44e674a721ccc2e78989574fdcb4c32e4345494f0cf03103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71c24ad33afc54e583e6cd519f0002ef5abaf8bc04bbcdce9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he379bcf17bc1969fb275bcbeec8627a8124f6b7d7de7ad4cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2eb52df3344d77469d61aac38c0908a8a9fbda04838f7810e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b973e4006df05586ae590facf630f6769ed1e059fa626c83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4af4398c0328cb870730ce9533563a3574a99db21714af6a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha707584d74af90befcd6da3829f6b2b50071426a8e4d4667f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bcb2fed59f143139218546a7b86165d8294b9b47cc5fe853;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h130765749bb93e00a2b0cd3de85dc98e142c9033e259394d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0294a904cd84c5e9133a2062d7b8ae805471070889bbf345;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h841ffd06be4a8f59cbe80e3198523951cb2aaa036a2e7a506;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51942774b080cc534f8ad489d5786f7d862f3d75e925c51c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe2ac385a49393018ddae23e00c6aec45928cb79d55fc0169;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h372c775cdb2b2ea6dbbffc72602ba89a2a135a3888a278b7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h514f063fae6dc66d2da3c1273887fa81844b1989352f6427e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbf0a87946a8a692af543bce563b5cf2918fa34582d02920c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a359002ed0739435d13d4d66dd2e078029d81dac9e450cc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12f83e4b6375144d71b9c169899245c4385a26c362dcc80a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f993e0c49f90420b7f7a888e95646f7d6ba698a56229b7cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1b897c433869f0eb09cc6bede21d5a1b5011efd7b88fb2be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcd490ca6de8cf6357c624cc44050995e60d562ca02a5e113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h540608e544c804d5bb512e114e62bd8a2d1d77739f97a473f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7069d9587d62c67ac9fc8b3e60d722e49edd92205415103f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7f6bdb00f1524e43b03cae0a5c1a6193e93453a9f8bdfa35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee470d82a33e293768d14dea8e0821985a2da94733d89e710;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c3350d6004ed86a81fe8d503cd05cbf1fe7c693e5dc7b5cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h291d59375f58ac00d6e3473a60d52aba2e2a3d060c11b39f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf3db259ef7d542cdd7a019a0eda3115c056aee6309b48e53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebb8dae7ec78670412af8f5d53b6bbdfbef1505b15b799367;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h698a900796602f27302c6c01fe8a9338f668cbbdec2123cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8912af6c738aa0656abf2c5d135a2d5b5da66e8733f0a65e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf097e667bb716019df1383b86cc948eda179a29b35c1b85d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c64de48c81d8d9575521004c7bba2c50e2f861ea24be1c7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc14b9ecbfa1471fd46ac4adebbd4ce9f7e6c44e7f6c358355;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51ab67511cf78432355fcccbd6e83fcc14d4796f248104d80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dc608d58793c5caa091f54fd295a29c312e53b90841dd578;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf534ad0e25737566fb321defefc2d76ba35494bfd3f5fcfcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfeec4879109baf2095a16d0022addda1f045b92ece5c20b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b489d520af4d7b634ddfd422c81176aead05ad0c9c84064d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h780f04a9aa5bb250a359834461b7ac3bb36532b68691ee376;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57e20c8c7ab0fb62dafc0e9c90b8255e99f41ba0f90481f71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha255294ba1f87e1a088b856fcdb2eda6dba9b487acfb9d16e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37c7333bc7a52352c19fba4ec52e31d5f37d59651605b3d0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d9970ea6ff26f630810142756517dd70cef979f46540525e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6b18fe9db86a9694403cc34bca9b1ca1cf4c2bc96fd91795;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcab79d846b1e5adcfbf34b8a434fd0a25aa1446434c624da6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa5593cc2d536ba00fbba50532a59eccdaf3c4ad0f1b09954;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1deaa26c8b014679a3a77979eaa99b1606abcb3f73d412bdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27ef2aa281e296c1355d062804dd2bb5e6c16b3f4a4dd22e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb061c12b0da205ebac7e22fd3526ce7209740f384fcf6a3b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h393be5af8d7caa834e202d4cff16633a90f1905844f3f0256;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b6873e7763fe6c0d21dc435d1ce3f74e930f55f07f0de37e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc88d7eb07509c15b3b06b35b0deadf29d7841e2a07f6359cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61da50cfc0ee9f6fc5646bee92cdffadf10aa29d22df89321;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ba8d45ddf64c74a1fdde80c47f0a6a6d0333be8dbb20691;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9e1730608e9dce3769a22f229b8aad4fcbb2622c0f0d363c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddc13c4827a6584d166dc0e57c9b08ec9624af842682aad37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c8770996f2d7d747bbbec270aebb816fce179f091fdcfa79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4ae64b8552126bbff3cac52deb5ed80770e703e5ea005c62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf951c74330098aa820c4768f0e23a5068b7beddd14746b5e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc21a99aad23298f61aa7c3fec9c75df175f715f8b57f14118;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fc337e35833721f8a36725950a43f1817a3a3e9448882763;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f3dd1cce9ded3539e2d2631518eec205601cb889bb6bc781;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19162ca1eb46d06dc720b9d3de0dd07633397a3f6b6e97db4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b01f6d015151aee0cb4f83a65d7c5be8446ad55a49f64f03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe2a193545598ce4a43e96656dca7170ad9aaac9f8b8c6b1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a4ea2cf0e61d5fd416ff64a4ec91dfeed3543de29bd1c1c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc89ab5fc09f0da30f3b930793d0b5beaee8f863781945bb7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd28d85eb192cb526b14809d63007ecb66ce1b3b86acf6268;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd70414511f6a1e529a281be703f3a7351bc6d9369a7c0aaf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcee0f63c83dc338060e7022b6612a308aa80ff5fae38b00a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6bf03f725b4e7bc6534522ddbf13a64a1bf9bf77e5bf0be2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h872839bb131721c4b1591b9e267898ace097c73b3337cea48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d475fd2ce5e8c79fbc8fdc2606db7a037b9404e519fa2dec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h799bde86b4d3021a882f6f898c3fafe9f5173a67ef38c8575;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32e801897d23f4bd07f042c73aed6b2342416d41441b85adc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a913867159df78a4c8ec3503e1f32b4fe10a177b82a293b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45bc55eb18cde1f350b6dc301c2cc042590ebc92302a4b745;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55c1e35456951b54b1bb5a7d830b43cca1164dba7e38c8277;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf51be064d38cc72c29e5fc699d47efdcccbb4e1029ee40bf4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f73a3b8d7a575acf1d92a32f30404692d59756dee29a1389;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a6256124439343b90d0e73faf049f2051beecbc20e95c057;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf4a9002e3806072c9edc87f9876b2c53b4a5fddd41dc7e7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a6872099c72a7f4f716e022a76c98f6d863a68c6b1fdab92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43d1dd954872c33e16b6dae0c63390a4657f8cfd790b82ea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ffdaf7f9a5a01db22cdcc32dae520ac2b1058a57c6b89904;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf201c4adb546f0a32f35fcee9d1f9f8863cfc294e2eee0d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h586f75c80122fdae89998fc82daa416e029cb4baa0053e070;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3ed90aa05828017295b794537dd6029209c4b21e34ee0f6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a06aa12f612bd6fad31660182de481bcfcd7c01eec7d32d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h891948e425d71f5b358282c1011899a67f8b8d2d736ebc460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3f1ec26c12b298d5fdf821ebd2c87be5c4458b7a475c17ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8e8ffec6997d07ffde1340739b08162fd9b96dfeb4db1f5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf892901bbd792ad8b62f47989d80596dd9a9d1ae3bf112bcd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedf4df1d6de7890d9a18f10f7529fe92cf13ea83fc7b5c91f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8551623c6725a2071b0811698120813869ee1e24be986ccf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haac3b4129509e03672ae66141df88117d116b7b56b14da4a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a1bfcb7e5b77eeb0415c52ce5f03b424a96a0086e714d63f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6309372f5c5456be2084ae4b257a7e0d082a52b343d428ca2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74ab9a369fa010caaf70a58dcfb387e6ce4a646a4a1ab70d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff80c7f91175dd3f37ff3204f18a6a9e449cfbceb05257afc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c5456be71bcf1b066cedf2806f5d9fd31e1ee7051a72df7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbac06d9fa468bc2b25342be915099968563ef2dff42a50a64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2aaefec1cbf693c8c3fa34ced407e93f053b9678022c8df8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he472235532fb19152295e76101505eaa73452e3754ebb2868;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h932de1c6a3bc2ee94b00d062c94d8910a69ed98f5d6b9e252;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5bb22d17a2a997aface230fda8d8dc33c1910e4b947a9c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c9ba7f8c0393941871ac77d87048c1ee2238c19c68184aea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99d56c78d7e38cacb29b23acad156350fee89ed3d5261b028;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b1656d8e1c17df9dc766acbb4a93b486d9e1b1071056c95e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6cdfd4ea3a1db2d90555cc035768a55219b73a3e67566382;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h155c88deeba8a52afa88567b018c05ddcc8ea9b7481a9a339;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4574595d47e37cf24f51fe012eb390302bf2eca72fc37f194;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6995dd3f5d3b61a5019766ab3468758b85c5f8dab725d4bb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed1dd1c927a85f31108794c73c0d430414b158aca06d8c80b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3418a6ebdc3f745da72c7c6e84f8a6d4fae33cbc782a2f018;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56746e1fea8d83077f1402b89e1874c298841fb56d13c6936;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ebb04a4410a705e642f436e0cb02aed448f273b610c2c61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cd8cafc2cbe55a1b078f756afa6bfb174f1949e5d51fbe17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23fe944f0deb365d49436c88f44a9ee1ac085dbd6bdc2d934;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6e17753e99c81c968c490b249c19905ee465ade7bae3e273;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b9cb69027796f99daf4a8c06ebaeb24f93a912d494e95947;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e83fdb4b5fc8a8620262ac6c678d83384f3c824b609aac90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8724e7c2676bd56e0f64dfc1e4e87f20d173d24b52c9dc2a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda6519e059a340bb467425e0d35219bee2368e694a8f93177;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd840de8c636aceb6ffe2af876a9277db46b11042cfe78fbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb1007d67f37af84662390f33d9fef9194317df2bd5e1be22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2a2a486a528fcdeb6052faa6838d6874d6d80cc734ea3ec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb4f1b7db4f9eca3c040018f633ce2497c3f5cb29f29f651;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha002d48114a515be78c43b180e43229dd6b76fc11ed56e61d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67e81c6e0f3e62fbd362b3cfd06bc3f04d45c127f47ddb9a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb63ac84a4c6ad6c27a63838b7c3da1e7b52de950840f2b4a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3debba2039520adba47fbd73021e58146341c2c492bb1182a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba9332c01f1579bc76dc998810bf7c70d11e8b576ae78a5ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h985104b5d053d71867f8d0e001193266e47867ff7d631503b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce2cba1ab5843eba22cf08847ea5692206e9c29b843de94fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h347f0ca9cd871c6bbd1b010e911fc98d53338a968a90e01bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79516db4280890cb3e3b6977967bf555f86e8c5e28da1048b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3e7513bf4753dbaa5847cbaec40e29a58c0e1390feb06dfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13c63b6af6f0eda9044e39d75e6a7c3f115bc7225c1bca69a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ca71e12b59075fea1c2c265779f77777745270433fb1e61f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d0b84107d2fb4b5a38e588b6d8d07722fbafae70d7c010cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27aff14ca22a7bd4776b39a50b2a06069d260aaabda9250da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5e9210daac3e25ab527b28efe0ed5b3e1f31f72259da5212;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dfe71877f324b2b4828b404f9f3ddde0afd49e58c245df77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7a96afa237c363878944f25ba19f44ec7534c05d8d192bcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71c75c904b5404730c2fba56df5678db26b811c3b69b7ccf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h184c14ab64e37676b0b36004f341cbca6b9c44a9440b5ecb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h774a23eaaa598ebb36240801124f1ba0c5f8e8f2d25ecb7cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h508e66900f114c8974ef503fe0df7c6e2ba7de30d7ef2627f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc30350120f5b8db296831d7da01dab9373b7963379fb2d00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ec17339534799d2b9457e773b32f8838a500d5aedd4d257;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he250fb58cd70708a2a383ee89e5d3b08cc17cf25f438e293f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47b7bb6445da2d9ef104498e0a1867621b0bd7893ff901e41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h622aa593c093750cb5f9a977fc7d97c168fe328bf8533c9e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a8eebf03ba11ac91fc6dd2d02fbfc708d3ff74da513b3941;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33e5db948af7018e2303ca436de9560981977c23488a60734;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb703333449597f1c4beec172963ac2d11f3a389bca7cea9ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fc4b66ed192088dadd53ce95bb8210a67d61310728263ecb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36b9bcfeb75946f743752d3e60538f84d2ef5b72dbd318e3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef42a0d610ada5c42a8e86802264f82dc0fc582eedeb9263b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b1554425d19c40787f4f96c0347317241d1094d380ab498a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72cdb6348253773b7a38a1dba276c40b8cbbd0086f210f1f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45b38c77d9d95c3c95119724df8f9a758f5328204f58998ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a810c5b8300c5688a7a336850917194bc20c643905b316c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53a6c24bc9d7f6688cc192bc056343de048371aab33ba6c53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h266558bf5de9bac25610e0bcf359d9dad25f2682f8d4c4445;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3f502e370728c406e886cbd46899bab645086eb9b630d103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1b5deb5d024c2cafb0bd268e96aad1827fa635d199e0690f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h608ac44ee257bfa97a28133174e5dcc219dc886ea6e767b82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5364f10c292b1fe2fd6ab2f4a397036f3e25642f82e8b82f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2124493cf0c8674989d0e0a93e4e3e5a5addfd2a3170c647e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a751cfc238802039620b1367d477940ea633ee85bdd32bc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49464640fd2d49d31d903e72d2981dbbf40f6798ee8161a82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfada9caa56a45ddc73c2373f2f6c4efcd38f4e011e75b1e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3b2dd6e0b44ab1bcb50b9b3302682eeb7ba28b2f83c11fcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb176e68c2c6cccb6f390869af2f72909a631fce4665dce1f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eca5437888d6adae7767de63e580654f0f766361cb1d25af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76d2d94a32f76e5a4636ffd979dc7b9646b941cdf399cc320;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fb92ed832aff3a48283f99cd523f005eb5c2fb0c9762e9cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d648a0dcb231f1837deae9834ef8e45ce7318be0e3fa9efe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29cf63ae006c12dcc434b636dad48cc0cf3a1a3ee37128556;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h616588fdafc8db31eac6e18d6fb32f5fb34a54eb4869eb3ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd589b82f3c5e64781fa903b43f626b9720486618e4b96efd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23afb6a289db9f63ec80b4a0e02241a52e491b03ba96ba11f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b3d62d18d0250ed8051712c38fcca9f9b2462d2aa75868d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heef9b61ea028101cb8cf8e19c6545344fce8fcaff8e670b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c073909135105dab060d64aafbb077e9c020403c3c915c4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h357bd4fea2ab2f392ff883b7e68105907476475b30162e830;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h804ec7175f90e85d681f568775e7f28ed077caf20e7115e9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28042b5e0aa5f62c5ef37df39414f73667a510060d9bcf1fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2035f779bc7aeb8d89d99622b72338891e78e2c61e6cfb8cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d47f123637f5c6f273416fc055a9398259e990509b4d868c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7dd5aea022afb16d5542bfa315ba36b54630074b46ddb66a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5689de3e376d142f70692e579447bf4bce4226f494c29b705;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbf7da6dc96b548801b3f0b9ee5845ede0c433beca76ad95c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1e648f6cfc93c597a9b4f02eec7991779a025c8c3bf6234f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87323f1c46c604f45d7049dfc4d937ced668b7e8cf8876738;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66c19ff6457ef9fe3188048b37a61aa5dc15ff714c254d940;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha28625d36a52c78e786fa7aa6d6974823fe2e3c957ac365ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7eac2d18999c0bd4f6828dc4298401b1ec459b2483a37cf13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacd1e48722d8069123e63e23ff48ed598ec8b281260cd36cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab7c6f8c4f102f9fa5097a6d5f73bcca1a822e37d2bac9c92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc414b07d85979ae6be0ce08c3bbbffd5c40720f1592b45bb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1aa31bae509e25f6954f75765fb19e0a24654dfa395230256;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h195b158ad81aa1a9ba93f6d5fddfee16c47ef5576a3588756;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf15f5cff7eb2ca5c22bf583c50160674f19bd021cc7ae648d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7022f00c44f2eb6031d779a4771b7b4377811f0b7be5af5b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7910ae722c396c44e3fd15daad7219352e5fb94df78e4f185;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31d480d57e6622f33885009cbb18becd1796c837a1fafab3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bcf7063edfa3c94ce7e13e4cd012cc8a68702505235e7e0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfec9cf128b015df5a670b5dc6690e2bdc558485428de6cb17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf40ce38b969bcfbdc85e694c82f70a9afeead497c38400de0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6f78797be58cb8705c4242125d69cf75588192b46d715b62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b1d572316c782b4c0cfa71bf3e965e41ee333e3469925f22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77cc7db7d2b93e949ea87197d45a0e16df45e127b0baeaf0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h494aae32f31ab9a1c8304b413cf0a9e511dd3f593fd8d9597;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1df682780aeaf6b93f09db51a4f768b9c99a536038196e6f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9094be0fe68dfd936946a2bfbbcf2b48dcd473413975c320;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee2b1e5f9470a22a682c406ae3d0c98830201131015385b52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99d61e2a3bc1b9aca7d1827a721fe02497ea1b5ce6b285a6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa3abcbed878e6c43731250494c2b9e59d9b54fb322d9f78e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha317c904985108e367e9545bbe5c8c3e04e3f694feda6f347;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb185d5d9a34b0520c8cb52ccd1f4bf9f2da47057d92d440e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab2ff71a1719d65015b4594ce7aef24d1eb2daac4671334eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h891efedb0e826fa56eda760dac86551532d2ef4a6a4dad7de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19d1658a3c7cc512b9d6d5ff4197643118a8a62623949cdee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h158f959da28613224ab7002adb84cd17a84ad44d394d7d52e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h812f76760dfc353a0de79c986f200b0b1e820c1f99461e548;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd255ec0b773c4b21d1537a38d9fe60384a84b79b6c31dc31b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha780ba0d82716174509574de74cd846250fd868a8b5af1984;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8729e12860311fba98c70170dd49dbbce31c90333c2dbacce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9825fc6458da9030c9c6d7c5fa935aac629a8d16a2c0c12d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb69324f7c31c81ba044eeb8a8e661e112040e92f9d4f56bca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cada9e87f7120d9f91f2653d9f14e8434bdf2b0eb7a0d7aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec690c8e57699b073e909daa12e103ec20858cd72bb832364;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h825cba7cb845c81d44d17cfe4bb27b6db71474ed8790fb62b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbce771935cef6e6f3b5f92335cb7b619da7c086a2d9b23e22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h162ca23c3067836852f64ce299ec0881ee88422ade03ef301;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e8944e9668858183d8740988e5a10ca35c05fe43dc361503;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93787368dacfa99c4b8ecd6e0c5de69cd4972c0bf6b6ee4c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h723bc79edc38b16f46b9a6c74f2b65a214fda450929ba51e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24b16c6ac92bd79a16c61b9c1d245f656f46c11afb781373c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d8c01d431cfa52110eadd813c4bbaea7e629cdcfe7751bc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h834ed87b8d05940538bda91189eb5fa79670ed8668c9fe5d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99bfd090eb255fd0cc3f6d04e85fb5b7936b55bf60b68327;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d15f05b4f2a9e1e7fc070982d73deeeba0fe41243ab62214;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5958006dba510cdb2fe0b38f251340b4000111bbbdb96e13f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3705716a353c1c42681c35c93730692e45f26fad727ded9a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14985ac3704c44e7c447c0188110c9debc96241350798f4c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcba4895f0064c0ee24d0fed1d6fcd64cdb947563fc338292a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9c20f1d352e3967ed84f0face5fe28235da9c975af3dd609;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35e089f1c61eb6537dddb17825f113b10fb8dac126a9fc441;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h618bc7891b1f78fcd3d8c0f0bd1e152c791009078311c169e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbcb4fc9e1e8061453ebc6977a075891a6186e9633d150c36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c059501e61fc61aa796bc79dcaf941c73489258b444f6334;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ee887c2669889acfbe7f9aca2f1c33aa053694a4917e6cc0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ed639d88c7bcad19cadd48bb186d19243a0ddfb2c0fb019f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafe2d614a57ef8e224610a294a0d9a793ee8be08c1feb1b7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haef3a166884b6dc83251c45ef9d3f2e6b2cd5631d3a58112f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c84451e7bde9373feccd11859fa909907dde6346378bafc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d9337b034b05870e12d16027d30dffeb4cd6b6a4f4f740af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd26b10330f30503578f3a657440691c345213accd64eea6d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc735f94d1d029f90e79df620d3743972f35f809675a7023ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf64f0b8070a9a9db4dc9fb366120129c010d6ed5584b54cd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47d69589b5ee556bbfcaf46a72965fa2190b2f8fdb5c0d75d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd78cb3c94e6b38b155f733ad052ab1215800dffce5871c516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc804203a57665e771f2b9d438b0b3b1e13797f367b10ac721;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5d264fa5cf4ea9d538a7b6832292eb147786ac575a8554f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba4aefc17243b73cf07c208ff4a00c52d1fd80423b5b8de23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h397c0d1448fdb9085f2c39e28252104e91605f5576172bfd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31bc5dea3c0937cefa58d693c984abeaa8a9aa2d95600fbba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb60574cd89c7f72c553e9179fb29d80781be601fe55b38b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5986e1ed87b3705841f5ae3636801e8f413b4aedde97c80e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8b1bc50539b8c960921fb08ea535b579ed8b4569622ff6ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fdd61fb0c9e7b8a87a2d7d09f7535c5baff7282431d79787;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3906abc60426e64da5335393c2d21636cb9c8dc275b7c5022;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7866b003a600aa781b469a850185ff488d1495cbabb0ff1e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc310627252f4342e92d46c225daad4529347cd0694d209527;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h717959d5be6ba1a36394f0df884301e2c3f823001cd755de0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4e9768350ef496ae464df67e2790386c501feea8a45ff403;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eccf893df86d9e9b32c7c1439d0a9f1bb1cb30123448d50e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4a70e3901d8998fd9fca084e8d39944dc2c64c584698324;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf46fe655b5a42a8691f9bba301a5539b57e94132f0305701;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c3ff89984290a88b57b71e22ec27ff9eb11e5d53fac0da00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e2f9e705f5d4431dd2cacfd9adac9122d491e0c639d93290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5c53bf42629b9480b32703b7f0da052c8e62c907667d1fa0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55f6a79c1977f06e381ef2a9e67b001633b09be5e59479ca8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9627a1493374fbf026a9612d6ff9e75070d892adf233ae89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76d6965373e098ff42e1b48b603ef49c8ca2395bd444ce48d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d80c4f9fb7c56f3e203094b1c102ece719dd7cd27c19f050;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1b1282ed1e77da285fdfbfcfa16fc34e1e1efe5097210961;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10a17651592be9cf6a7dc8d044f8614f449fd24d734b5f93e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h132856083583e40cf8cae4b64870b70f568566858283e0325;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb99817b416f10bddd11a48489378d2640d95349318d459370;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dfd9b3ad94937e01d6dc2d8a399edc70d9d09891014d04b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f2f768490279d8295fc9f0996c881f86d032feb2b464b801;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff5f33408df1835e77caf0f22e58e7641b0fd5338b031ccd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8cb015585f452900cb6e8f1f50f776e24519c4bfd3ac9c26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f2b09cc8ba14e9ad32ef5d394b38ded4fcf629d8773899fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3694835f1a6ecbaba4aa951efd840e768b6b3c350eb1246f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34db1d43ba1d6d66a04c362879570b52967af52336da73d6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h704fbbb3843d2fc439853453560f4442766368a3f7a4d59af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13f1ab0002528eafe63873b742e8954518c90cce2afa88a13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he086cdee95d1aef7679702b78e864950edab78d7b56207303;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5479e93636bef5241016408d524a71599408513de9c3b3f39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc698888ce8b5e0cb77fa838c014e7db3dcb62702b44138055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94f53c6bd87a02967695e97e74d0134a93614f05bac2dc4f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h866b65f1c98b410d50ac72d817ef47030601fec84d1b7a4d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a6f008f481014c543e2a81c6198498d3d31f3ad483799929;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha58dffa97583eabd5f331b20dd1e0b02d997b0847c0cf9e05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eef76fae5307b390dfbf12db6b2901b56b4bd79de88e9a15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde90b390e7515fdce603fe7b56ca9ea3a4d670e0ca24d5826;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h989c55784fd32792c1629d4d96869be6fd3c3e224261fe9e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdce2ff30e06677d6b079c29d339fd13fe7537495c4edbaf31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7540a2bc2cd75f80a91c73d0e5303584b57de59bd34f79c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h722cecee83b794ac3a16ac1e16eea753404333ffcbc3b634;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b1be015dff2ca36d11c4b3d6f90a1220b2d9121f72f9b4d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4c311a6b7749aa2218aeaf27658e74a23f752cfedc4c3d1b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccfaf660a314607210d2cbec2fede5de8d86a0702f95c36f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84127656ed71cdeff07fd8f6807de7f1129b409539ac41421;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heba987c9bfbbe2169f092d2edb3ed618507942dd39bc1a349;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28ad21fa356b0819df3d60969762bf52b43f2221406e6ebdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5736bbc4d203e51c7bec0ad29e2a391fa3eb0493ad9019ab6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab862711c1ea85cd2b6633cf4c9ed280365f19582073c4221;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3eaf4be92114bd35829891f73387a3d3db006e9a2ab1b3c2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h424925ef75b279ec0848acfbf9100b9a30e92ec82ea324ab4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fa3a838b0ca5a724b8cb580ecf12ed5b94a80a77fa68afa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a1e030cb7c439c7f5efed218c15385ef382eb8a5a399cb56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9222e6435734626bb89bf5d5f2951571913fe59179e8dd5f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f2cd2663d534a0fa819023672a1e469b7399d11698f7137;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4460492ed8ba31eacf2d160e5e8e8bb9713464b881a4e5f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc073d3d99dad0e92d0a3ec27305bb12a8a0f587101d018791;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf53bb17a0d76a624f62179e1cf8993f48ae4f9d769e4be7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7584a3846f6f7cd746cf0dfe99b024cc04d3ffa23a495cd86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a66ce0106f85d1567a2e9901df8193405ca183edf88f7a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65965cc160d5c51e62cba4cc4247f480833b1356d4bdf93a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d0bc6e16db38b07ace6c9ebf6581230ecef631dfd48f3f22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab8864aaa9613095895c4545e5f7a39effc700a6d59fa1b13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha519989b4cf79e193109ce1ea5c6c382069cc3b4859911db7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e37527be847712ab99190b7c046fb5354ab33f9894326cfb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1fc9ac52683c83355e6311d4fc3a5e018a037401b19515fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8b6c1c370fd56887d5aa37828f6ce407012f96ac65eafc7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ccb9b8aa9053189cd67b2fb69f2077e275397c5e7a9fafef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4385005746157813b8b286c2e3e2c6497227db6b556ecd0e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f3563cecdca31dc1b48011b582ce6fdf24c32f4f6095ca1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd94676f40daa8d37c423ee2d2f9660db7b9ba2d9b7b4533b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d20d7a97dae4bc1b747876552d963e3805431ac6d937ba84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8998a6e77af1d22808554db787acaa4fa4901aaec67fe19c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50366bd07835287e76ea197723675bf5f1d2131016a065bac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cf66ed94e8109054bf1d6f71194287630893842290f20353;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h448974b075457e9ee92af08fa3d9535889484a1252c34736f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12b5d9663d80a604b1309c2c3b07ca3548c11a3029dfe2c5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3af3f2b975a8c04477fcd7e67154a8d7ff52325e663eeba68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd93b06db2b53ee72378db4aa58836261395c8414a91e2fc7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eae73414949c52d8db5839c676e0d69687ce103332f35f59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc63dbe4c40b417bf287dbc90266616921d9fdda500fb2a13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51268664311385e6e7170e434302333e7be00cf0633ec7bb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9591364d2df12697815d70de9f1054efedd86b174ff15511;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e04ea8a9617b6c71aa74f3f584f2e12d2281a5d3141ca251;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c53f2dba9d471052810d532062af575ea05915f63f9867b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd00288e563af4c448bb31bc487d809b53f14ca96eb6d8ec66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91521cd54124f6cac0a5c0bbe5b21756f15c9c649794e198f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfa33ed391bac8c5787ea70b3ead6b867998e824c1a1105a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h152a59558b526f7abb6099aa886f4008160cc766ffa8d726b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33c7f33d5d5e7f20a6c720a4274666f820f5ef32c3d702832;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda723ddb5b60de3f3d09f360103c83bf2100b9627ef17c63c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64320550cfcad5f6b5879c93be412caa2b55bacb5ae6431ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5170735518f47355ddf93af0bd1fc95622dc337bd91feee5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5213042643b2c27a080c99f40ffe7fd7f530c2fe9d95d288f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c0b5a2ec5ace3e65d044f5198fc39f6c0e0e3426545e6b6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c8d8914e7037f2637fb8c9829959dabdf788e83214d40aae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ed308d3f49f370261a24ba4f14a46f99c4f4bf30a4f4b05d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h546d7ea6eb228bc282f9eef819a6d2faa00772ab221da398;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9db4eed2cf8c6ec1953e0c25d1490013d38cc25f2e477385;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3885e806709aa6acd0414dac2026fd2d4554fc5c1edd64d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h844a91e57e99ce2b5395a334e931c5d4e770eaa0509ff72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dffb454a28087748850983305b1c60cdf191f09fc1cce31b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fe6d8fcc8430264dfcba6d5a8ae4815474c76f83b4038c02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e3f4f00f21c320ed5727110122f6e44e181ffbab5c1fc985;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1e92d2b7700f8baec0e514f4b47981e11129c11e416c3a6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c9b1ed94031fa5eb81cbb7edd18ce700004d5777f016d04f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2891747d36d15b657a8643dc25683289a5df382f831267bf4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c9d11bd3d3ad64c4e710b2550ae75f01a7314016818df979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6874cca75c66aea68f091a1e6981990479ce54259360c8f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0070e0265191846704b42a9ad6f82bdce681d888da99e682;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b64184ac3b56f13d46c3e12664bc87a248eaf4e912fdec82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h953bb164db57d916f689ea4a263bbc25c952e3e67fd15ed7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eb3c82bb1a61ce933f8ceb363793ed183e800d6892b3f966;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3d934988c298e6d6590c4160c7a62ac356aa7d93be166fb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd3dc5c15be4a3d8199dda837f5d36ffe98e586ab6bb696ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h706c894b2a156b52b252d05688bbaef0b8d60dc65ecdc2ddc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h852d47568a93816b0b92dc28c93563cf2ad71420c3eaf3fba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1beb528338d200d5fe9cc69e08400298dc7ddd41a7223e26b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3d64fb37388916486fcbf98ec913ade4d12f74a22fd97fac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9ba26612f1a2e53f98dd29d701233f0f4190e7da0d9d69f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe9feede122b940701bd82505223f18df570245ebc7c13fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8dc48e11761416ad41db3f9a58f2890a3cf626ad234548e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6616d350a57cd407f2645d9426ec1d1494424b734d3349246;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43464d53e98585f053be3308339d5378377e817411b206102;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17ded67a490f73caa5ad41dfd1ab2f3871e53f168bf2203e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc44b57cf079403e754a26f147227262f3762b2c803d4526a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85b511ba617fd29968bc28d564516b0beef867aa6c8f247e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31335046cb3861e67c71c0f63e8ab52dae7920c5fe17ef25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83fdc2c958458b62a5412503856ac0be3a9816e6c54cc6205;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc11e0f3cf5ac16293e12b1a193b9e9f515f9f3a5102a8b4a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf82ed2679cbf26e5b71617b2dd95a3a1987473e90a6c0e630;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf2f4d29221b4dd74131cabb1e6b36aad900dd55f0110cda9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8360a4f985fcb0602eb3e2d277ab06e5c4ff62e81d438df5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he290496a8ca44042e4f42703ff9db3703fc9f59107419a9b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdc28ed614551ba355bafc60ec6c1e441cd292732180b9ea1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd419e255a00e185a189b28a54e6499276e9c12cefcc238447;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e4797df5028f6864fcf6ddc8944f57b6247f45ceeb4efd37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba888dd100ed734c6d5fa8109d3cd814f2b817f01df20996a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d2a9b3f28a89c81b63b42b75e673f189b26db09a1f5687e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf15033e8614e3afbc9a60f3b8d754be7f17977fdf732ecb2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he567ee44d00aa8177b1465259df14051bea2a28cc35352782;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5520b252ee7a136bb523f5b9e0760d483bfd02354507075c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6b7de637168cc1baf1e078b17860029f619f5552c385c771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h574f11503f3c3474f215eb714024e220bd68f8bde3dad37b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ae97428d45ee24c8c8a77086497b4454ae358d3af821197b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h626b9eef76ff4fb720c8110f949b04f28c816434bae84bc3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb406f16f418001df25889a60b2068beac97c2b32a3e1f42e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2850f15bc52f38048c90db957159e1b0fc67f9b64ab693a34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3f547449a462b112346485ec095e4c229621d017b11863da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7777fd3ba21973635cefa24ecc67315c18302cd03ba4b31a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h239e630d90bef55101104db7ee10df36d5c994af030121690;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41805ef59e198b280874be5b41eccc6c1613bd430c087af4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9084197b31752f98d4b8602a976b7ac99d3b27179c81caa71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cef6226ce94c87d255e3580369ca24a5f5f4a6cb631b16ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h796ff4b03a10fdf3401ecf8b620079d9c90d0d77586b8a578;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaa67f113446d8d22bfed25fc7a6b88d51ec12b2a3ca7930e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he433f2f7847ffb938d9b61b78acc63c704a6ffe3637a9ea3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f81b9546fc9cffdcca91c5a0a7587013df3dbee9ac258d9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd07f526a2dee81ba34f8d8cfea30ee3c8ce6d49bd88a4ecce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43e55535f3940d0e8062beb19bd34ab4df73412b86f899039;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf22d8542fced01946ff5f0797241f08e5ee94a693b86796b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfa7b0971f8a1f238760bc6e23bfaa381539a0c23b5177739;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e626a154d34e170af07541c1a11d701d3f40b55e7c960abe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aa38dc6a41d89f7cd8aafaffae3d6b40adb1b68d74ce4f43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde4eb8b50978b59da7151daebf3e0a3aa7e30d305e9cb446;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h123ff45a771cc0e5bc10ce5f21682e42b5717123481a0a9e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6146ce3151823a444f85a689fb0e56366ffdba0d549c96a83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h136cdc6425d0e24f4656f8e11c18d64f68e469b1b104df8d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c569c105c7109b12a0188e1e001289b1d25ae339c7c04728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79ff584877661d78bbdf57e859b46442bd1b1137c3a7bef73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1eb67b494517c22f7d2590abc7d8f678ef1a5ae8d37cbf38f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2044716c9363fbd997b4bf1b6e38af6d777a2a675932bc3e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5b222f2e95dcea73af75a142b1ed3352884d17fc26090e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6789f485eea28826a1b5e11a589091c2497dc8456db254d3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he960afea56e9062fc5651bd716e9e49036a1a4deb26c884a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h847d60ff51a2cb3232b17abcc6867325c31a432be4787ed4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea6db986fbe08882352fde5d8e9f8b292155cd1b77207d46c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc49822fae12c18803c3f8aab34c19937b5f51fa18d40cc608;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b5b555c02f50ac948f8e782ae5626bc5876365a186ab2d7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc544cc142e801cae9ffc9fc166b2c3132efc5809faf7133d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf10c05dcf8a326912fa8bf087caa51c55033d298e2dc44717;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb9b444860872b1e5725b2670fd4c9328efea8a68e0d43437;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h393110684292f562bb06ab598acd09df153a93d5cf4938cf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd24d6711bf5c151fad65a2a8484bf7e6a199d76ece4e21bfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11ce982e6052d3643d4f97ce2476c85adf4d88bd81d6f4003;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd482b56999724883dcf75178cc9443069313f22c4530540a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf70ba7caddccabebec0161de02ab27ef1670413c5b55e1fb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h815ad00c2f274fb5971cea49b8792457b2e47d26f6f95036e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb47d88ddf57f4f0dd5ba90f88ce6b36e3c06a5343a17a913;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80c515393ee14d848a2d0c9563acf66769df91910cb2f5013;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c9bac7f6b6c6bc8e61c7c580d035f8e29a44c6e61d32f3ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haff9d3a22f2f3e7e0ede02f8a477956f4862a05c358a12930;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h896fa76e0f65870a0465f3323ac5410e8d78fb85c66c0ecbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h464ea78d118c07c43f8211f481f8138b5be1e1d0e96f34f7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2235050c3f8a98b0226ae58a3769d7511efb5e6bb96eedf71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57243271fa32a6837f5645cdf2f696e87bd1da6649f360a8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9808e194995fcb9555fbfdf86df28ebbff3069d7b2446353;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2b3413e38aaaa969c7fa4f982367b2781cf1a53c92fc1681;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fe182e16bc55184673b8e9f9e4889295a87c44c5128d0262;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e780f59938aa71fcd4cf0b9bd1a05c7591ac919f546ed66d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d6d3b345b775f38474c4094ea711d303ebcd944ae472cd6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1287b5844c63fd37a6f8e115012ce3788aa66e6ba66364fa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h120a6cfd883a20842544130016995dc7ae611551dec4192e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62ae730228ef665d5d6f50eeab297cd45a6d31a9ead80b7cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9533c15efc2f93257cd86b132f71e42d9f6e5c1c50c45a81c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cbe96f612969f477a7324d9f874f6c837393dabe026a53bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44e34c4d60cdb2f3f769d497b8e56bd253299a8a68494637f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31a806181fcd7193cf22582b7b85a3fb9c40231d5a75a50c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde40a729b0d3bed4ce580543f7c8cb9302beac108fbe3376c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ee10d0c139aafd558e0bccf8c8f3a6af88df5a90fbb8d986;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c74736c358b75976a86a7007a25d7a429d16035570edecd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc536716b30d3f0d63c00cc1516a5ce3d1d9578dbc56ab466;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d714d83dc8cb01c4fce70d22a99521fe8ddef02042a27762;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96032eef1a01995576b84be6a08618aa5322e928234a55a80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d6b48bc514c624aa426b6356bf241d111525813a901dd532;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha06e58ab5d393c49a362a0ae84be9a448468e50e0a6e7b275;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f3f1f73bf744210766773e03f4218832f26f8f0d127592e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e41d7e38568b1a42ef396b34a22ea8b93ed0a4b5f635a658;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e92fee3cface4e15756bcafef6c617442018777235230403;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d8fd04415b211ac02fa320ad29bd83de4b158e7219aa201f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had3f021198075985ac506de9213beae0f2d403d9b1ddf0bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d399331e0c630e7fc51a87515cb2abcd0ed36f0c8808198;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc687cfde4f1757a5677308999bde628205bca1d98ea2792e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82d5c7ef5498696b26eab9a3dc6b55e0b9bc2f58c05942768;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h739564dd817bad4d9d0cf7aa261df3e822adb70a98931241a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd829f9dba954955a1e1a9207f1044bc2d1d2d457f4286bfbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ac5b2a1699a64b358480152199b913d7a7869da83fd96551;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9e6783b4fdd54485b764e08def1b376db0cce6949c4b3bde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h389bed98ba621c2d25c41e6f271be3e77e5082a7d884dd061;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce838d30ded2c66e6166c1db54885a787495e3057be49f6f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h671de69b9c449f3551905cd786dad4cec2dd3f61cac224f10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa1f747721e79f69f55f9b593112f6dc5138f819675bbc064;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67e5581ef6890263b27cbc37ad04555537920bae3f8687d18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c6e14fe48c15a0cdc26bb5426c99c07d48f1561def572a60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0023a854698554df975b163c959dfa1044d0b1ad24bb0814;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75aeae44bcd8ad24fca3aa7e8fe7b356d054a935a339fac31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19fa57510b6f2ae0b9eec8399930f3779fa95db9ce450d16e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8677c2b805bba6f370ed56c4cadbb456e3fbc3b5fa56ec251;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h318bef058b76cc03b12ec657469852fc9912f0d16b6a9bae6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48936e84c1180900d078f89b6fe27ed628b4b2a3c3042e7c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce93c8ed347960c84b3057a84e7cd13e3bbca7ecda0674757;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1cd3575ca1c893be1318d263189bb42433207935bb3b1659;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d44ea56eeaa755cde4e54b080a984583215e7c93a6a91d0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8bb6a06f3535b1e8bfaf914c2317442599d2ac073f8015bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habad90e0ae0f42e9e0a4ac1f2f0f039b66dec2194d11446d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51f30737248234ac3c3b16d72f4bb00c6e72e2ddc3270fba8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eb998c4daadb90c1a91f0aa2fe90ca650c8177bd9807d8e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h523eb0947f65390c97ba87bf68b10b11d3c2c61db5d5ffff6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3686f2e0d57fa7b2f1c1bb19afb99a61de564415bccf61c6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3219c197a1ab3e7a65358eef529213fd8411e31a71810ee16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e955da94920c5291c1a56857ac3abaf3b964de90f2f322d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb623b49f64457d4f023a533ce4fbfd2e038e9f0593e80c113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72568fc4b9f908d9e3196bb145c32e3453568aca450914363;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h211c941da18a80ebddc560c04aa74a20534c9a906c818b333;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h668e04c0e4ca4aa89a18f03a144d689528489e116f88e19cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heccd8cbf90a54484319d27854fad425aa75c97621e6255ad7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a007bbca5e321fd0f8ff8f2a8dbc8343c2184dc2291e57d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31ab0b04cec8f8fc8f05f7af4fafdbacaf7a03ce74b7a240b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30c1093b3279798a64ce60ca1b2b5ec6bc4e24b1d9f3cfd7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf85f058b75492782c065e94d96d1ad6c462fa5dcc4c6db17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4de74dd9ca476b8fd7a5f2b2e653c8fb9149a2277e16451d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he69f7af6e31a5e4cdc6c1f7d37b9c3980d36b6e8587cb6fe5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eb8d49d9bfcc1e8e15265e89495d0146c8e3f1db796eec89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e2062eb9bdadd80deadf7ad0fb4ef4b3dd0e93645df8d8b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb533e8dc4683e14f5c6d239b327cd96c334646c7698f6156a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb484108330fc4e1f7316d80783945a8fd873efe3750a88498;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64815ecc0525ec67de574448a68aaccfe0a5afba2fcaa2c98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d3fabf6857229467f1b7800d6bdd73b770b8795d6c6f62a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa106be05e74fb65a76259fe2927f214decd070b525fd7fdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0ba862a9e76ad88d9dbb99923c98d0eeb2678675d8368513;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddb5065a662f96799aa142cd0710b978223ec6947469c8655;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7b1899305102eca4d3ad1aeff935eedc80d80aa944ff356f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ba02adf1127e3b5bf8e95862f51319a5baa488711a063b85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ad3132e197475f512e19ea0a88460044f76cdc1ebaef637e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h249023abce0eb2b0b800fc5a0788315a3db235a8e7697905a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5f04d1ea6a15bd90521535f5291e767d7429d2d74fd1410c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb8f208fbc0f8af1905740e12c0b5c78a724ef43e39bd3a07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ed3b3b5c0ef600c002d25927f32ead887e756afb31d3a702;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9977af4285a6d23d8ce7cbf3475d1aecc6893d6293542ef7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h624307c0581458a66a3e55142146c78617f8de485e2521ad4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88c38c1f09d62f9fc8a958e8fae521288cf4894fc4260d70e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41ded2dc375a3aa52c2e1733278059e788690bf427429a4e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef6eaae4b9d3f0f1bb1f0a3efd4367635ec824b82a05b0500;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d1d032a84bc4c1b0309766f8495781510f17e2e0a39ad205;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf18dc0a428a78b3bd67c6bae28c2cbe8506d6cd6407bc3a2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4355126cb46f15fb4a11460c05a621f8de9c0e08d20526232;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc8daa22bf18662ee6a7d57a018ce635d0ca3d11f976096e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ac9f8aa310721eaa4e8bd1764edbd18d5730e1c9a4fde111;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h289fdc0e424216b72adafcf79eed0e236c5d6ef87406cbc99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h940ec03adb81cb557875d017c84b0e714a960f0552016deeb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab5349ba330a900ccaced2b3ed2842bc8a5a44d469a12c3ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a577054035f8aec0a2d96f3928c7f99530dbbcd928c9fd43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ae0a0570188ceb6e37493af68fff254d60a039333a8cdc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc909b0a30af441e86a6357c8ac94e010c43660b2289d246b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9376a279e0f275a9a917e4c88f63583481612eaf81372a88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcef06ef91fc356e1cf10fb4c1b6bb4ade2504231075dbf1cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73a1bfeafa30421b246cf1d62813dc0b870e50ec50a8b35cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heda16c3fd152c286f03d032de809b26b6c8edf454c8476f4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40b9dcd059c299d09b79701d4ecc414d6d2291809a2020415;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54ebc19b60ecea1a6f4670fe319b0443dd5e0aec8fe33d69c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1a2cf7e59fd3e2176328bb9de65a9532811bff8353145369;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63e9d93be4772a206fd362d4a4f6ed85599f6b28db2732366;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65f16fdb1ce5f32467a23a6221c33b5e920d277da5767c360;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h593570a0bda4d9a78640995eb0b9403827710d0668ead288d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dad73e06fc028f87217323207e2cb6fda106b0a459fa4efa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39f78c8a9bbadbac9cb066a1fdf54009f20de6f007cd5b937;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26779a2733032f8791ace1367fb76f3b95557a44d104254a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h713ed447cf28663a3c3f251122fd11c042593ba1f3ec2fcf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96b5805288a4e101b6dbcee0d8813aee0a7f9346aaf7297d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4442f883d666e2e163a511ac34f25b7723f777aa91816ad9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2b93696bbe09ae8ab1eed03b1c0965d9384e16cc35d0de26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h256b440638d19d01a5d63940f2d267231414705dc4dea90dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f8abc60f8eae360c56dcb61c3121606e0c2d89e67e5c7c66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf9ae578fa1e7d5b54de0c587b2d92b50cb2a96c9aed3b963;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd919c66edb736c29881951e7fc3f5d4f77d589c8729b3ef1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2200010f16b4f6ead2bdb4c85089d7ca46c3f9cc1f875dd7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h548c5eed17c9bd2c3e43f5fe3eac42eff91a401e5701b7458;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10cce34f2105c16e49e64eae9e08d1a619ded39afa549598a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d7ed755dc2944c81cfc24e9eba944c7e7ad0d9a0f6dd706f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h647650481be0be23ee079481d4f7039730ab8d0b32db24c47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92f3674e677a64e9667d22d9255e2df64b8f7a797f251e444;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e81ebfc4ddc00c973faaeed9ef2c320a5a91069f53c5abde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3cc99f2bdfc136b8534611d70e3cb33ad76ee4c9618d522a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5515ad4f67ee8b8a38d3551f6395e96c6d92403268af9e907;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h621754448577e5c2854ccaa31a20c356757d390eb1b648ad0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd172f65eead354dfa70ea27e4e3e5d4d86ded481e62ce9ac3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0e7a0d1cb020a4e39c7e86a266479f5d9b7add6df0d7852;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb73678cc7a6b9d0f3181ab1399c83bf758a82c5afe47521d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dde19e0f6625ab0027cc7a1fa87b67e2bff92e9665563bba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h946f910d64d82624352b2694b451b7c49bc9f6b7b875212dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f954b1c38107774293198029e567f1bf1a82fd0dbca54d76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a0c16012b022d949b3ecf7428c0793c98c2341540e75823d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf2041499f7ffee1d628b842409ef8b9de7a1cb5004b3d0bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd5dc034dd77521de34f69b7f6c2f074e9c13fa50a56d662a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h669c762741d13ee29454234d253ec01a81539977acab23607;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h810d991ca9cc286176426c8936af4a120bec11dcec06adfda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcd273795cb79c995ea57400323327eb0a9f50942e014ad0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h328e179bd1e843ca91793f144880ee1db260bc525ff6f1a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d68e811acbe8ea9e8dc273d7fc47e6032a790cdaa985cfde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bc9432a10601703b21bd6db0e4f8b3f97ed43cfeed2fd46e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62d6618759688f8e268fe3047d2d88df9038b70a513d19a27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37ed024c5518560cda2e5dba50736266166e9fc2ad1092656;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdc376d824f8044b0b69aef3fa56f817e895769765274d56c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9510c496c76d35173fe6012877b67706b64ce6601b7cac1c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92c33989672acfda03521dc6eec228dda75aedf5143ea1cf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6327a65544444208774e3700949fcce890c593dff748a92a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a5653e46463fada34ccd08aed8cf86ce560ed03cfb9976e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4651e46a9773316af2e6a5721354f5dcff408b97b92e534a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80e9602e9cf169b430aa33af702169a74f2ccce402fdb7da3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47ed0f1eec28841d4de929127e09d3af22eeed0248036aa80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18fb7132ad3d41e9f0c7eba4c46b8cdf2aebffa4a3ff674c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3244f4426778fdefa686fd458a353b973865d7c46a241a30c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h363329554d5e6fb2aa3d27fa1404582401ea2c222bbaa536f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf73a17ad6a0df9b1bbc690566967e9c70204bf2dc750c74e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7811a25876c47ec6463d833267de04a9455afe8dba49dedb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16b5f1c390ad5312aa1a1337d29646a5137dae6cd1ea3dc90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h997f124268591cceef48da355d753d9d7081b99ab0140b82d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b9ddfa497e151399ebbf4cef20d900ff6df19e8b62ca9527;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8f6f0e0273a8fe9e3503ec79e44c74f29fd62cedecf880a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e3266baf17e75a2103115ba74b985e9862cc7bab2f48de70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he82232f9bc4c84355d7dad636c60673db348408d32659d6b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd71d6a05c85cd0534fa39a42e31b59739579c504a7de1367d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb835fbe62dce2c88eab8fa8f290a166a096e0dd2651a2fedd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5612ecabfd2ce0a01a598899a4a358fe915b77878f9b8f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h324cd3f9e1db77406f87f8131fefb6f903dc93b60579ffd0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb91010893663c9b12e18899fd7a51134c4ab73bc9bda471d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha86155d5ee8a136619504ecc49d65840a04d9ec805a019373;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49a301597536670b8a9856f519bf11797dbadb87f074b41e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86bbff6d033028a8ad2f6206f7c191c6a6c178687eb078d23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59aed4669821f3675d077e141eb8095fb2b851341d7cfbd0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf3a763697d219f4df4f2d490465c391730009ed036ae6565;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf84f5fa3a5f3c179b8fcaa6a902c02311dd1657e1e99c2392;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28b252eb22c3cbd7d01e6e96519ba314901cb963a05915fe8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc6f06a03503c51b43cef0c101429ff2143721726ef98169e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77c46243f45683aecadace4feaa6d7271418f5b5e972c9b3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f83ce8bc3b73c052803c2abe1269cef72dfc97b9f3c9559b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf796f401d94368d593133764afc6ac71934a95004408e6c77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6b44f5e203ed2dded49fe29a1c9b5e1060ce9a42957ec0a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59553001af033fc98d316de957817c2ea87725192eb97b471;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb541a4482aac6ca80cb7b63d6ffa87fb0f092ebc11d99d0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b07533d5f3b570106087f785fd3e1c5434bd35630a5881b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b3bd28c1608c4cf767ae79d4b4e311dd393395abc0c27bd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5d34c0024c7be828d9fca25cf5b5d4985bd4c9145094ee33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c98339bbc86636ca23964d341cce0edb416049e35b3d80d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9d149e62e8c458aed59fa8a056161a2fcd02252f310f3043;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h391fe426900e67cfe3e9f6597c992e139934a081484b10fb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h922930c2586370ef7fb9ebb8303691c199223560678d68a50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha879562be3846db88deed502f968da1b67a17e6b88e420da6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haae0654aa6762106ff69467df2ea89b7fba58dfac301e4c42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfe724216b836f6a4bfcc302f3d15adeb9e535c830c41d7d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9945597d79e905c44bc03e3deadff16ab1cddd6839c071ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h282ac80173acce869dc0bbe3cb2429e3a96a4d6b8116d6676;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h244f7c6dd59ad995c964e0ff2e02201ce929b05fe7ba8224b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h459ae189d6f4025df3fa345c2c58b99f0f35220006cabe18e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd0a936e9a6936490fb51d46cc25d8de1f77c67948f5496b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4be039f21132acac7f28d3ddf1081a1f7db6d92344f96f49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fe342af3758ff907065c2290b78447bf927adfa22bc8d4ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ef001abea998dbc3e6335d0433c903bbcfe265afdaef793e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84d655c5a9b3c75074154a7a18ec5e09809352c249989a43a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde06c63040d1cfe07a4b90b1d9bcff7361d6ae3df675c8cd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2eb436d896a54cb59b9a16fc050221fda2e8a1188f28fff5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he28df5dc2c180d704c011b30a60ecc12ec13168429b54a06a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa0062784b7e435f4c7378b8a63312c3be3abb920072a3370;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45da04d966dea3a098ee7f00dfcf4b152d5ad259095725602;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h980661e1608a9f60445b2dbe3e8bd4432cf0366d399803e9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7000a9ac27b7128680ba6ef746c237952b4bae06e4d8dd6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d8d9c93b9f1142fb9b16edccf8e9abd839ec548eeaa3b262;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he28163632f85255b04dbdf0a4b81dbd711ff55b37ddf9beb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb30f51abcaa077e4a30d38025dcd6b2b012d1b78cbe9940cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h772063f03e83b04b98f613354f47ee802d732d40a4d137293;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h753c654ebfc46d9326267442bd0ca4dda3385666733c64996;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he710bce8a3addc89c827dd1b0fddd428d432addd3d9ac82fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96c42d25387cd792cc5ce0a7dc908afd426dc2bd516054f5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3b94f1cca3110bd2c549477a96e4e918fab5b40d693afc01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha470d91c684413808d2d474d19fe0464c31ece9017cd2273b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5fd19f4d48db91e42efe391820930497993cbcdcab2cf032;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h911d42cc8cb870f3d03c92498cc642bba3cf02fc858f2a26f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4eb2a43f55263a8e09f31775d440f35cc16d1b925d488f15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92ab1ccb9bc0ae8f0d6b60c8fc4e8d7c0b2db17734447d3a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h257c553cbe129f2830a770f905ea853180823437ae7fc5224;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebb01ef354eb8e44922f577b41f8b0511674064a23c37771e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc88bc4fa12c9fb516f22877579cd55065c8389b0dd071175;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f85547451ab8dc93043c5e51705682d583fd7b6f04aaa74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadca905c1f6870ffe115d03c87096e476783dd0aa60e0af7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d95d651239ff0a8eed0ee0f6a684075e5b835ddbfeebf4c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2644aef7fc6de368d8e295f8aa4e22d1d8c0b2262dc12599a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h817a6cf01d2075c12d7aa9e449cc7b93d6dad4ebe3732a8cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2276c5b636d1e893ead8b0368d24e1b103f677627d93d6c55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b25ce4522bf543bd974db534a43a69b32027a5478f317d04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h937b9178d96c8927a9232eabf83a6c8cf2e53130309836a3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dbb3fd34379025cd653d49dcd7b7ac23e5755ede305db3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ea0e8e4871884879b325799276ab420d7aa7bf0af8d44eaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd87e5e858f0e993f18d1d35f23d5425587ce39e82c7ac415;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e80a5e0b4e124748da558e5264521c71e2d0880859aae4e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h768a4ae535de1506d308a9986c2e4f95c909e72dd4f54df2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecde8aba105c6c7ceb227a3ee025fafc2944025dd4bc7363f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33d2d32e0f93db1c25de45cc4e3422f5334ad6c605ebb9ea1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d2e5cf4bb8223f15fbed405fcb7ed8ecb5884fda112625e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31cb3c57ddc66569c88ca8a211338d00e8adc4a55074d446b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5613c56a2bbf952d6b63ab3687afd8119025b7f84919993f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fa2cba7f2bbc0e40e2541523aa37f12c2aa98ed5cb6d9a8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha46f6fc087c708e9fd9a59453dc9174314d3e06ec46a7bdbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65c29b9d0dca6a335d6ed47bf80401ccc012b8dc35e00d949;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96b415c65834771ca630def9e42118cb76ca2c33d0a916e86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha88c25118839d9cb89054aced9fb6dedc84336e9f55e9e67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dbe03e8d73c84480b5bd00caff85bea4b34605ac190fb217;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6d5237ef4479e85ca825b710a538a685995de2dfb81a6177;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b702aa6f7061497a2605bdd13e6d703f379d22b033e63268;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72d14324943ed3db64f5e97936f3b5084d57214cc009915e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he61e6642d6c5e90067db5eff56f124c7c41e7440a34018454;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec0ed25a126f1d579e95c4c039891d386eeccc7941afd0525;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3fe52d614867298d360bc661f8cfa7adcfcf1773338dda24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b88fcaf998122cdf77ee3cf164ea520b4fb43b50c75b1e02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78ab63c1df2ee1610231742b83acc6a1a4621cc7966a1c0b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99cc75748f7550697c292eea36f15f3f25068969eb368822a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3646a4514597dbaae41f7f718d7171af86ec3c90ad3dd47e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34d39a19f78fd504d5fe5ec7e787e58d0ef8d2bd4199659b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2500a6a21706ffd18911ec22e647f89f993cdcb8af56c065a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha764342a232f3db90122d65d87a9ad18cac640a24a53b0a76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb274d54c8703b7db451bd244a61f41b3d20907a06e245c869;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac0e5cf16618ec10f0558c23a824cb8ce9f9951afca34ff84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f2312b60f9166a1ecd6c5961136985c9b13dd750bfe2d074;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b17e8c0c5f6d9b3591c1e673fd090edd3b5b775f23d8bae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd818e3c04a3eddd14b8a9786d5ec89c0cf75129a27b605d7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ea05c3f10402084ec98f220ff7d1000e029aba3942c0e90c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc2453c9b8a90fc7837c1207bdff0183693b7cab73942684f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5902de4aab98d5d1e9a19e0797fb360ab1b56d8874d3bd70e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9887fffeb31e8dfa696de32fd4d0c35f9864317eca991623c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had1f8e17fe4150860f99c75c453d72faa22c42f5271bfcca7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6fc0eba2719d66a9d4a2286cf746b699e6f85eeba5b35a76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h214b0a7ab73cd5b5905a949fd49d9da6cdd877413d9f8732f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he171f27100e2ecf52aa38b0c06cbf1982779c66c4889a4e21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3ecb9dec710e58be723503e28af0fa5d09e183f179d118fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfcdcea07ffb3074f554e4a5edb25abb744b5017076ead5c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h330f0c7284d554ed2509d97a83a745025072181ec0dd4ea17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff2aef71da42a099124abfd825ed5b5e41759615664496eec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h894b4efef57ff996551b47e159dc0ac3d7a2d26a1da9f95e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9c2aed82ecb3884647d60e1d01ffd388d806907224e68ff0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h474a676dc6a3fda90c4234bc22dcc994be12b04fb41cd7788;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5acb2158af390d5b4dd0da661fb47285c155f220c149c4ec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb59a028d7ea255391e46c40e60791f9ded6bb19e84ed1b16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h381a5c6639fc7eb85db29481092b932fc7b227b6c901cdcf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2902984dcb7a0d6c2f93ebe49e9f4c88c44548c7b77dd2c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8692263402d9da9d8570f97acbef41dd880c5c43c99334a65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd54478148130e5e1b4479477815f7fa50af7a09448963b634;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf4bfff534eaf3e03c8fd9e79edb21a780f5d1303db7a180b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b97274f60a7f6ee3e58a5ca270c9253781525061a05377e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddc3b22bf28cf28c1b07b620e416ea9054d5612c732108fb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff0d1c11c444d7c08d4b04c153481092fc00a4a721887a3d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hceab1b3d76f578bd4a80054fb31ad5ce35bcf4b1e06ed18df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9759d3c07b87ab17c7ef825542049387cd6bdcf2ad8cb9867;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee0de5c40c77a22150b5372a8dcc2218ce10d2084eb90205;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c062d008c3e36a656d7de8916e387dba4b8dd395778499e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3cdb59b886b9d46d420737c2984b86956b56f06deda4f672;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe3798a2f3fdf2f48e659a679a6af10b83d700921719cba40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h128aa3fff61c222bedc98e4b74eb64739291d063e7e5ca75d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha258b98787d52b360f76bd80fe0c6ce804775e0f1a652ab9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b3908b5e1cdf57eb5efaba54e58a977885e75f6df7f05086;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29ac8c3253b1f6f06e1bdeb9cfa778df442b1f42ea46993fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbb3a6207df68a28559c028d618307d83e18dd1406f14b754;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf41a62f35544e2f84f31e152e710c320fa7d080142bd0cff6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52d85dac3b7c1892831c5b400c9d2332ffbf22dc8b36f977b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d8b6b0feb875d707fad4c86522f81e1061d76d917cdab17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he638cfc575b2b8122799f612824826877c5999e3a9f6d2989;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd9fe44e348615d6d35e98a5dd29a5e52b0eb3e6904e5f838;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2a67b8f9f9954fc486e3b08bd26bde4633107750eca54a1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc4dee526797fe50a4477f3bc4364e8c0f3c9035d0af80e7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ba951d59d9323a42a205c2dc98d5aa7983497791275663f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8393549759dc14cec13403fe50e11cb0d919afcf044d3185;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61de242e746e06b53f28d03c08565d6aacfa43754ceaf673d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79142d9f7ffb39c7c7e9cb861adee9b64f5c9751dc6f4f02b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1afa1faeb2f241c03f7cd656b8b7ed1dd0013952965f9a950;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb64e4d183ec5055b99a5c6276d509943fee8b9b7bca7898df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28cee0c0e513c23dc9d1003b5db96119bd6aa759d13d27b10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27296fcccbc4b7aea79eb0a11ba42a3fe7dbb583aadb66a10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae449207396586012becec9a98bbc7603f0d15e2a6efbce8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f7e31bd9bab79ea0838a97b73a7fde402436b4c20c21d321;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2c6ee8f14f373c1a9d55e971d53a615d44a96aaf600f5923;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h434098dd0ceb16a8708942444752877d65b44a617a0915e26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4c32a521de9433c599a1e980b36e306712c21a39c15ad5b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15dcad7c6f01dfa1ef10f6aa65ce133c9baa3e59518549fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ace63e11cba1bd0fc034aeb7cd7c8e67690cd5877491331e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbad689eba12c49cec8dc20d939ed3a0fe283412bd9359ac3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7924e256ac4f27b80e49802bebcfd7cca84a3160304fbb80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4947b9a2323a644f92ff686bf63e7ad029535160d828fef74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ce2d86cea26032b7642156dd9ff6e993f907369159f9e1b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e31f7d2decac1402ea03bba151cdd7ffa53c98de741a8f4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd20569cd11d25137d258ef3d7ecb959a6e34913cc64e43d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0ec7c291ffcdceaf8341f457e54d188cf9e0ad66447ebad8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h249ab4092a9d77196e18a19ce0ff8df00020e5f1b63244f7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c61fc4ee20d18148bcd4bb499abd9d72016644a39912584;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84c12c8f3f94611ef540547f23c79778309f9718753ffccf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b930ba790ae898db769a56928803d1cfa4cd52f24bd76063;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc678a26b567bdf76f1168ba56af7e56ff854521d0ecfd374f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h688aaa31b1e75d419342d2e1d218ac758c650bfaf113f2261;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he40e26a85e8daedd1d81fbbf6ad4f670d04d5b7bcf51806bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86465d8ae6a0ec80629a38633e1b48c44e4b7f2aed1f3bc7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e7b8cbb0fabf7dd956c7b98c112ae0412864f264344f1722;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0e89327c5dcb08c68307f8f458106c0ba31b2e3d9ad0fb63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4f7e9964a58a58b6085b655f053eeca2cb8a447fcee10133;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5776555ab710699b0b35e2f550e5908865ec4132c815a47f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h843b57e98356d67eb48269446806c440f099de5571539e9a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe8295de35ac5b2cd64f46f8de5e1275d4b6d754a3fe75954;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbc9edda387f03cb822bbbcba1d5faeabda2463f9c6275bd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf643df9bff763d638d69efcf584718f9a2e67e567e1e0b9f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c780df1c6da4f04f2b37a320093c78f11ad96e0272476ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7627001aaa279707551b8472713e3ed9fb59c2503ddf32a5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd376f46f04581fc18a7e6ce47f32d74a344e8ed3ca886846;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7120f6cfb8ec24c06604b45fc147da893427a248c686fa095;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h596f95f9cb15bd87ce1b26699c0b098cb08e74a8325c37541;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cdf078c4f1d6e8409cf53a84fbe6f09471c974199bd4e167;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe56c7f09d5c26c879473e9d9eb10fb570c4c038ae1f56cf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80f5e10c337cfd84b31dbd1c0f3e8e22a0c59350ea01a6887;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf73633cc3765fc5ebad2ae867ad460fcb9acab893081e5aa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29dbc7316bad4050b4d02ab20d572a8800e58f99e466d1d27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h223ac9b3b759105cbba75330fef207eec8c97c7f77c988d0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38d2837a3a6a198f59a649c60eca779afd66daefc49e8b4bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91462dc80a25f64703321eb10bbe181332aaf6f0e6c67c38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda496910fd9e171e49ce21239c58b266f469b3383aa3d02d4;
        #1
        $finish();
    end
endmodule
