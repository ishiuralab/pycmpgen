module testbench();
    reg [24:0] src0;
    reg [24:0] src1;
    reg [24:0] src2;
    reg [24:0] src3;
    reg [24:0] src4;
    reg [24:0] src5;
    reg [24:0] src6;
    reg [24:0] src7;
    reg [24:0] src8;
    reg [24:0] src9;
    reg [24:0] src10;
    reg [24:0] src11;
    reg [24:0] src12;
    reg [24:0] src13;
    reg [24:0] src14;
    reg [24:0] src15;
    reg [24:0] src16;
    reg [24:0] src17;
    reg [24:0] src18;
    reg [24:0] src19;
    reg [24:0] src20;
    reg [24:0] src21;
    reg [24:0] src22;
    reg [24:0] src23;
    reg [24:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c20847e9bb59551b306da080ff9ffc774bfd6081d38a55f459891d2ddb53973fe3609e71063b815fa79ba82a8a28998b430de8c742c27b9f45de41101e8b284eafa46eaf574d7706349000dc843e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbeccfe668bda8905eb2072ddf6f5755b937c6192141a3066a0b012e864d43b17e542d36244c4eb12ebabf16d549b5fe8ed625159d56452fa776d9f3580c6745b5b2a33c100af3f7abc29d51cf944;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f38ef75b8f565015b61b2f7fb3b67195f1b3443003e426dfcede0cc4b40fed14dc5fec92671c5592fd1a84e231354389ceea34ed79e4ebb385f75f4c158332c3fef7e10e52428c1a346eaf8f3b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc20c134bff632abe01bb0a9aaf3626693304f39ec3d83bfbcbd760a1134fba5ff9e8174f3ca4740858d45cb6d51b0c78b21fc41ebf7c7431ef49e8b73d6aef9fce60f0ad0edaa53492f5464ee85f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190a584390170abb73afccace7ffd7b7aa924712e84be959782cc8ced4580bb497f41d8d75da7c75db08492f46773dd1e15e07491a528990d5d71db7424ec620e6e66040ed1054b975bec95219882;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6831fbb0df88773ec490f868a4b9dcf4eb79ab4e5c83c20d3c08fd2ee2bf8e78b1e9038f32d34850e4af17790ef61b1a859004eccca38f31719036751f83fbc066f7f667b3688b9c5c65282e2b9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3e7b7a31a96500046668c7f0d7b92b220a3bca961c6083b4059d04b335462658e5aa18725f6324129767a62ca16108abc6127617bf03596f73b7314aa59756370d7b15b8e5e7e7f3c5e66eb15eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a3f963f5a7bb52b0eed087301b83abf630c05acab3fd0a6875ae5f4755999c1de71f00377d1380eba1f645e45493a3c86ddd2ef28626e386affc53b461c076f11a95298bda673ffe98d4baea89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec51e28aa4774c1754541d48f40109a6ccdfa91420ada64b315d006bccaef4a36002a31842c68b086fd2006604a554fa6ac3993eb8e79e397fc124e4858bfff3fb7843af4b39bba0a97aee3a6005;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30ec47470836e72cda66b3c329a5c8e73b3623ddcd9b7967f79d328e936f9fc30ad1d22803ba3b90fa536b9b87fc54815c76040ebd3e6fbccf8d6f182d7469bc33dce9dc619d0674226aeab59bf6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he750971a8ccf5875c14c96409472dc034969cc50a2a4a16d61da85655e269405b6efaeae8a20edc8c1cad01d04f91eb089c118ecd21bf61caf55fe7da7bd05d5f8fd80872075bd11f3303590a2dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1068b131537011a9cbb8a752bd34c8342d2ee6b44c254a0bbc478c3b8eedbee2f1785f5575524044ae7e3b93bc251a5fa5848f946af749c43ab64a03d28ad5b5a3dc6b9fdfb3684e6c111a873ca58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h959e2a6d8312d7bf3efc3f33bb24d7876d57e369a624ac5abaa000b0e8bdc8e80385a553af3fde64fcb7381361f6ba85931a46d05713df4542142b9e97aa1eccd7c2691a090f7ebba9a1e346af5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1166ef0589347842a9b6ff3da067248acb0745fc7b4309fc09797858247e4b3ed42d82e273c040f49f8810a35e0a628c16885bfd7e57119f2c288dbb0d195cc548e67ece678ef79c07c6372b42d7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e4ffc36aa834e86e250657bcafc3fde89ef3bc5688c31fa11d7f15d4b86ceb3dfb0fc3a3975096b8b6d58e68ea79107de591b676f81431dc062a1d3b3774830be2bb53c03008d633ba580a5e6f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2f996c29acf7bfd4741120da0fc3f0965956f600038241c8eb3c92ef06da0dcc9a8d8ac6c40202e39434535e98f137031083d6b1551cfb0d9d321c4605544b3927acd3f697ab21f10afca1a7b7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9c6be4273ebac374470ba718a3062a7d4a9117feb7846572df2c4eb67d66e7ed2944eb8662330c875365a077a95ace5e28ce92e125320e9c7688b8a9ce1202168d464cefb3cb802ff6a35b6fcec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f43b015571448064fa8607579c04a33fe76e5036f4d2cf4964d17d6fa9eda46af04b9482e098ece00abec5b8f086297e50ff20ce2bf3e6788aeb326dd898aea99ff3c017b3a0b46266777929cb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f28bbbe5437fd53bebb078da6c410325171064a6d46cb99d40d6d48c1152cd6b4c37df3d5beb95f42a6246cc8fb8c1c2c40141ffbe80a8e9fffa97d52e6fbcbeffa6ba644db1c75eff91b066608;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17eadde5fe669eb58938aa626c5f54bb0fcdebdd4edb3c78bc584f1851463c7014ffe02d9cccb986cbf78d99ad481a36151f5ca415be9f121939d71ed92259aad776c6b2e4bf19f757f1c5c03b605;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171f6c12059e1617e6f3ae9770ee6a24e0a8965408275ffc76471c0145d525bc0d886d672cfcd42819321d969449bd4f534f7c0fab30b4e6a5bbd9fe17b4350289ccf483f98b1b0d2684871d44d36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28d0c3e9bf027ab3ba914ff82fa400b0ff2a82f004621107ad36dd13dd8384c906cfd44bc078a016056930d396618a69a0c3ebf779094106eb6c90c6e0ea0dcc138a71001018c870fd1b3ca615d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e21527cab28b0dd5f295ad88bba74ba0c33464a6a776dda789b7dd8ece8c750d3bc8c52d161aaf98b2ed1c0f2fe0ed1e2180ec221bad1af2f982262b0e1574ace37ea8c5679cbef0cc38770386e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2519b4fa926ced5fce4fbc78b25b968189d793ff5511d776cd948cfbd425079b115c3f54bf171aa1f3c256e7fb917e19f5d5aada66ab5fb5eec38ac5a3165edcd8bf76efbc3f693c6cfb06d4eec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h905f04c444fae404e9aa1f9ffd8a8bafe0b48b07f907d16b365e6d78dbb078b1d7e19ca4d7ec16e75ad09dfd389cc4011de4e92acf1cedb5f18ee85bdecfc059f674bac9a793fdfbb59dae0ac6d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122f4c759387e279ad27f281ec93089c9ccad37faf249097188672792f63fbe0551b91a7e2b8da3b91220f5e614c524a3ac9349e458412ad6fb4a40b08e6fa917ac70b1d2b46cf46c604a26a55eef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecc0f0e02cbd5191b4040ef5bad3bc8c49d59e40bdcbecac4cd7ea4d668c42aa0edbfa2e3a884be3661eef956310cd929511255f5b299e248e9672a529aa3b3930b12b2ca8adf575ef2250a1d92d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2546e0ff2dc4a68be02a8584211b15728026ee6e5c4e68c608282f530eafc86f53628fc2fef8dababab93ca4a995cdfd7ffdea76aa73b2a0f52bfd2b258e02c06cc165f9dd531bdf48b3a6ebf3ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130d3899b40e5e84768dd357d575ce4ae9736587517f779de298865384a1942b26434fecf8bbcda7c22c9f0585af1198922c2aea4157fe4f286daf45c8ad9872d1b689fbd5e4fc0289177c89c19fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a9353498565221693e7805018ffbd5a2c0e971523b0463c9729426a31c3c3176b79b899b1e27114cac27955dedaf86de4fdddac7bbadb22e85f6d325df5fb011dec349816475247383bbee38ec2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1934066b5b04cfbaf546e0982e16e00eee70f1b748b999553b2cb5b1da10c3634809ac8d939002383bbc931fb82e53b5a12e5bfcf368bebd36236c0b96b8c92b263f563ab0466f7f549e53ec919;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdeeaf70ec14cf663c6a98725f0b2f4b69d3b6e88492b50485e8260c743f62b8e8c508142d00682918b4260138bb26b2dfd9113e3d2dcdae1271c9eb56097c15462a327cff7e4c7afd075a9e3d70a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca01d990d547c347833e0fdd58b2d9cbf46529d46259c30ebc8b468c3b416fe744c5649d0a2dba89a1c5fe8132dad4b6a80233ef4b11803566fef343a9eb9ab559d5bb3aff57b6a0701687c6b92d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb611480421a45446fc30540b8daaa60ed8899316ece571830ac4803e360dc8a615e2b97a98460bba183ec9aec992fbc7625b4bb6ac12f2ce089492598c11b2bc8f7f6d276e451c5843fc5f192bd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0e5c20401fa320cac2cfb19f5fe0f0b2e7145b037cb08eb7f3188e32f10becff93ff2a90a8d6cc175037e70866e4133b61727ad203fb4738b7aa6b5c34049feb2f2a43c9ed3a21ec6918566f682;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178fb6d917b4723fea52d7e1be285fc9865ca2b8bc72b75040a09f9df578ced7a47ba380bd792be5a7c01a8a704b94d182f241fadfc72bbde831be6d333673a3286bca9f2478aafd65347aeea3474;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1130eaec8a20d22370ee76404436dc6265c041fb845713406af329d799167a09762f669bfed8fb3d823e46f3d9e0c68b01ad8d9cd8d257f4e4c64d49e12de1431c6b62553ce32b4b98692016f7542;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61522839bf96758abb5ca6cc91c5f1a912703bd8628011becf3a43ef687b53392dead6638c02c64780b1d8dcef0d48241049fd4d1d9de2eb9caed6429e699ce42a45678cc8f59ba9c54ea43b4787;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145f5ee3a56770347d768eeed3926f1d69e29b4fbd193e0a9997297feaea465f47364195ca1cdef911909da87c3e901cb5ee4d8312b3d4c7771d1b33f43afefec93e4774740ea77c156a9122bfd1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182ce352561c538a14675199b7849d36f855052f6f920b8d60a3dc579fd14f3e060729e510a6c22aed70fefc929261c030dfe47ac51c0239e7b841bba2da5568596a4b41807cf9bf51ac19e3b4709;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a609001addde70fcfd47a37fffa4aa567e8a63456984ea820e897d194e5362108bacb62d17c85baf6ff55d4761e7f126f9326ae324841bfa779d5e38b89585941964e4b180b1ef5cef0d4592d7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41d57ac89724d060f23fa83c922900d4a93bbcf8e0b1fa5285fd7b34a1a448729b6511d00e5b4a8c91d3b5dc60704bf39fb0dd7299699c0476678ce415a37a093c359fd860edaca5511e8ba287e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1523f9d6af0701de9ad3ee8620160d58df5666befdc4feeee7b4da81d8edc02213d5438cd01cc225490626009deec5e40f32e241b7bc146492f31b2738fbfe7a3820bbd00a584be19fdbea4c34afb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a91d02ee06fb0eca580cdffd1c816b7daef2cf22aadda346215146f5400372f0ba3dfcbe0e69b99b49309a3d8de90a059bfeb10dbf8c5c62cda09b2c11984e33e9b178d891b4453d90847eb90230;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15567862ee5f4906ff7a174ddafe3cc9774ab66b592d8e85c73738c456efd8d9bec31aea752d07232c4b7eb878a10deef18c8c3fa9e51e98fbf7fee5472154c10c51aa77843878de554086d70935e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f5c18f082ce1eba337098c459f5b13623acd6ebd7d748db468887a985186c28d51aad2f5b8bc7d658cc86f26691ee246b39336876252e145f5d45285b0159e49193cd08274fdc91a1c269989ae8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0439741b61598c17a1f42489db405ad4c3d7ab83f718508744c44074bb9be0376f76f5710313a12fcdefb23dd5d104fb276de04b2ec5377a0e0e33f5ee8e0a9567a4081a95651d2ee8d80243d87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ddb2cf171b5e3a014de5584dc5c0699663aa395db0df77eb85a041adddfe47f53404dd1e9025d392218215882af82ef8ccb0f56ab119ddd8935c35454f9de6b3d05d6014afe7a64d042e6bc0df9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6f540077acc1e21e9fce76d9b72668b3b2eb0c4387088c264c3627f1f5f33b69edb201010a119c83eb015ce9dd986ad8d272aea43373701cf1be68e12a1235126fcd5263a84d75b4c6627b9666a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbcf90ea6ec57d40212a5c8a7a077b122366ccd27ce26861310670440f8cf048d782f2f58e0376917ee072777f06d5b9bb9709b62b8e25773cbcc418c683e5bd29d6dc157c8546b5c21bc3aeeb0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha07210283128f1e0a2aec817f730ff48a574f3c414c6eb34ea68673ca6a084f01ea66acc13d2d4ef17cd4256b5e9a3e7c1a704b827a574f2793cf56bb7767f27835f7f0217a5df348f3c3dc5e518;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h676e20be02a068fad0a836b608fc54dd805a93efcb9d4c63b5cd964df9d7d6256f71408804d414ef2be28ff27f548bd7570cd1b50dfc2f009bec41fb06f55705969ab90a1273ed47162ede9f6037;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c38b00e33b0f5e41d264e62f1283ce9a5a6e84f8cad237ce0b6b36bdd3eaa276cb38dbb5c1eb85637848295d81f8b8336d270a259e65c4bbeeb85f8583b3ef41234b8abd853bf728f4bff2700b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5079db7bbb41cb0570aeded44656a61a0de4b9f94cebb5da7c291748e881ae2449fe768aeb284a048d345c69f0a14ecebf0fdf720b856f7aa0db3f666340e1ab64618205c806f42459a7752109a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b9edf1b8b679d2641688d9ccf607a1577a19b97a71f3aa19f17a2236ad868b8d7ac9ef777fa07e3a5e6c180a3239dde37d445d617584e22efa444d12b0f4a0b3a105357f03eb85c7eb15a375bfc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a28762ea68f9ca211b5bee0881ae3aebf41143c1734286d0cb244ddfd61f5691da26767215dfb7c05b5b414042e298389e844f825fe5a73010b87420cf6709566799028a13b9720231c0fd9a6153;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47cf4e53c6c875fe200c39793e6c1d51e757790ed046b72ed9f5f705e8bdc25be1f39070e92169b0ecc4f5577a3e53951a822a4e7bb0068cabc4bd856bd11b91f83dc19fe9fe04c149c35e44fb9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c77b77f6b44730799c0176f3648464aa7f1d0ae5f2b950fd45b3cb3f5e188f05d92093631344c4d2684a6ba0ce20bdb58cd55bbc5519d7f4b8b4a54e44a3a1605588a7a9752fef65d3640a05888c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19355c481fda7c214b0cd6bfc260f842c66d9c6fa4e2eeed648101b1350e456ef5d2db0861b9dbfe4f84fab94c01c960c881305965426e3a1a1a5c094c5c8301eaf14e68aa5284e3f6f36af86a04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88e48dcbe6e04abb9d362b0a4831da886c580603e5631c4e3cd2f1d2f84dbc509bede5dd48b0b5369c37f2d2e8f04ac8b4872d7bca2479d21df7a337be5c48ff1d509a663cdf9cf709647064a417;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h288511b72a84786745d16afa231aed0cfc2f94bdbf510f04924b515d06654dc94d6d7a3649cdee4cc024ef43b2834f76906bfa29643b2993e84e57925b3acd620cc13dafcf0291a85a5d379b1daa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b8c484df8294767060e7c53f4a9beb81a94f1ca5ce7cc1bda9f4f5e895415ac3e88fa0a167754129264d7e9e2b4315336d09b9b6c92f93b0d916141aeb01077b73fb0f8b63f613fa6760317c835;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fa524dfbfbdf26af5ddafc5e4bed8cb34cfdfc9a2949b113cb8636a93e64b200453b71ab21dd97d5e967c3dfc410b7c492678358e1a33274e110798762d02bfd9c39c6c27342169ba48644bda49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f8611315333b604d4c985dd4b6f79ac93e66d5470f0b2ffa75965e39bc035cd8530cac9cb76e4038d099642b34db17a02280ebfb86e26ed9259099aac4f00876398a846b600acb9893f9fcdd9dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7b6a564fd239e4f03af53962326d11adf0b7c34c210db007d5a232cd442950de6bb3a55624b6ca040ef8573bb38a43a6ea8515ce255c03d0eb4ec9912ae51b49d00e1b886c1ae80d401c0a27079;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bca746732e3e7c8922b9407ba361c1d6b11d26bdccba44668d42160131aff81f7626b441559136d91c0c8b5e6988fd28040aa741eeaad109fff42717a6be9269282337680dc62bc4215ceec56773;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf4cc66100cac45478a32132d24343b41083c993d152d781f11894a9c1264ebecf1b82103db1f540587411ae53d9871adb3a2e3eea40a27126bfb28bb9f4c90299512fca3d50ac3d9371cd983a10;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef1ff6a603e93892f8cbb368c10c37b85b889c626aa0bc8f26d7d1a47477b3bfb70c712f10ff2816207ce4542958e6ea9e7572108aa84da1c6aecc28250eadce1a36dc595155fcb0dcb6094fa674;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3655ccd54b9b4be368a90fdaaa5314aae15caeb404cbe347e1669c968b4b4d81661b38e235f193406c39f9ccbcc3234330d21c12b152f185ccbb56dd75c3bf1aa6fe005752ab76b9d54a9ab2ce7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he73a09f840eccae8331c5c64dc5897db45ff6a11dbde0f23d72e765090e8b51e650e2bc8ab80babc8769676212c9b03971ef0390cb6ef823caa948584a3e2146c01645568dbe2138aaa8adbc1009;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8b1142d9ad0ee41da53ec410c1d1bde7bea82263a8b61fb068230974ce2330a233c3253670299478d6fe363ae5e7f2743e4cbe9d4dae661e026b4015ecdd8737801732852cfdc91327904b6fe02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d420d8b189c1b0e9cfb4458dcac67b1d4011453882ae89dec34e869a6fa47a11e5b97ed7bb1b15a972d6271265810b19585fca8978c68f73087a9126bb56384057e7c8e2aeac1f2895cea418876;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf5d2b8cc079fafabebe09ebd22cf8b0a222d4ddbda6015a8caebe6c4a1e19133b88db4c791b36eeb285176cf0b63fc7a4f19f21bcf5ce1165e131ac33ba8ebe2982e03e837c1a9fd272cde160c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae72c7a51f2e27c36d8f1e16e02b1e92a0ee9688343867b3d0c4c5300b1ca553848be349f2a57e41f3ed9f2bd532323128b1ca1401f5efcba77b6cb1b6a1e63e3763613e41b27f5a96d3ccdedd55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heecc3117b3128e67998718ae5f06c123d03dce5622a512c63a66ab58eece050ff8b9de90a5fd8f24913481808e5d3578a1e5b6d9088f289cf89fbde40574f88d5f540c99e5b4d9affb3a2b9ecb02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f44d9a6cf325ca57cb6325d15cda07432fdf6254c90d1db4da80194471b4f5f5d90a159f8fd1173e2302dc44df17f013f91fb6ff1d677389dc2fcaf2489fd5452db1a07baa8d3133c40a6912c139;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1913c1258011f971679abe0d93faeac780e0b8e9a84d445f58e1867ed7a047139071e41c8f8679b0f25b6b647ecaffb10c865ff0e1de8aa1b74a3cdd16810d2efa7ea01d3ffe4a480f94c17316e1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb5e95b0c169bc331322bef3cad356d34b611c6eebf8726c2b98d9224ba3920f8bead453dd25b581937c1d2ed9b11d465726b5837cbd1849a610c35e7a54ddde3a95496e33ac888d76900177a92e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95851f21dff68505e88b5a4cb543d02b547e609e6ff4cfa1d63d283fe97c2132eda26b91c6fdbc61b2459acf74e2ff7e2481c6e739105185d20a1ce09ddebfe7a8e6aa0bb8bd7435d346cb4e4066;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfb992281a89f78abcc573c2fa6e9e2eff511c9cc87fb2e1f6f21a16db067d46c2f72722398f34f62a4cfe0fae96c0a1000f1ef58c6e9e0879b32d927ce7bf3db909c57108a845d85cdc3c912474;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ed022ab6ee7d69d383b05ef54f50c6e62e7acda55699600c3294cde03c8c93f8b24a5aab7972250f335b5bf55567dfb651903e6999ac0bad3d4984d4d062e7fed7c64d49fd4b00fb048f430803c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14455605bd89b80a19b3ea066d25b1a2a709eb637773a5ff1505098679a0c01f4ad3bf89e714a28709619123e2bfe2b4715d30d17e3bd16a0ebf81a16cee7e4538abaa9c2b41de257103203f01dc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154174d639de7d1feb7903ed6a0072fe9a9596394f2d121622a3ae78abb09ef648ba002845fc7ca970d3c49934e4e2faf35191e467f69618da366f21bd312e5c5ef0318ffb3b1d485679a46e2876b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1236fd5ba3742472d8d4df657e7bbbcebba014e75f7819afcd5708ba30f08aaeb88669730b5882794c0dc352cf7cd958e48aa9620482c2bba51ea5cc40b1e7a660d61a3517c23cb09d215d63bae8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e753e01be988e2679403e0b41187c5c39b582ab66e23a1ba1dbb9af9c525d2d84442124e579a33a1fb360961319de661ecf6da5b475cdabba7af1214baf511123a588736c756cb18755e0e2f5b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1745aadeb5fecfd4ef32de30a6cc7c9792cf9917ed26806f424de7ea2180f8ab2cc9fcb7e4cd5a09fc4b27bc40ae1024516dc60fcef5d2206e6c5c94befe3e0559523d4e81d947ecd731f59d48668;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb83f2156b70a19d0ebfeea4790b0e3df04f23410df6639bec4b20539df97a17fffb41769b347d27b4c649bb6cd3ceaf48b0e7c70e3929d9633f01e5c226886157af774125bddc8e6b64a8b5c3c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d2f40e859a8605a6df2b992d0c8e888b59d0a0de90c1cf512f885f0c7b7bb74b342ff4ae507bfca4d84bdeb4daf567f511a0f8c3127b2766ea920dceb3d71b47ad4f49679699f98b5bf2fb4faf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd826d954f4a8f718e9d1af0416df6101adcf045c0d21b3cc81afc53ae32a61e4bd43ee3814a16726c90f60462912d51c50092dc7caa52c7a51afa35726e28984eb646c941c708b46aa7445e4f2d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c15eb091affc8f0d9773b5837f58e9c6433eea2113e4751b05c0a809cc608a3593dec7cce94fd7d8f94a00488aa20d4baf2b3cade0f0b3a94f6fefb3912ee6450a10ae6f4c5b7a937c381113bc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134afb22415f69d3eee9b2e9433ac18afab9ecadd02c50a9bd757edb17293ec5713f07947e920f69eb98dbe88463b62c0f63dc9594b7feae0aad988fc87dceb96b020fa50b82db8999811c8a50921;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e3ff4b4c460eb46206970a3bd0ce7bcf4172deef01dbf2cb026384623664912aa45189b290c5739d37f3e53d3c695c32d926c82b7929d7c5149ed3765db5f5c7a60f126be9b985883cb14d0afa8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h147c8f192bea642ca542e13f579674ec20c3f746bc99f491a0e4bd38f026e295d211cffcda2b7cfd3555396856c3d994c63099eefb71bdc7b702b1e6001aae48a6b7e352d35889b358980b94f0271;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1743f119e26748a5d8803dba2ef74b4cab2695c62d3b1f7a452c667a24878d744a7b7e28339dbc689a97a9b770daa3d0888e1ffd349e2b8c8bbe798f68cf7c3d13b2f7c3f4114e2cd71a4abf71a7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103e3b4e3bf55b503ab0a1a50f0c060842207c574c20981e6ea711d6e3ad2b8deebace53c542ead4eb8d401b64d6fb51e920d773edfa5078f40b2834e486cefd81a95b9fc8ed4043b7c7b6d0898e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e36a6f7db5de1999742de300bfcb65af56e25ffdb6476efb48ce8813c5014c19cacdd7f0e8832824a5fc2906e6e4185e36272755643d9411318aa4e1596ffc8112e27cd1103c09d21c346c912ec9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5c68d2f62794274784e6b6c5275ffbe0ff4dbba23ac4224dd5a336f71c35d2f0f0104876a468e0913e03cbc7d63fda5bc4dfee2d66631e1ae5a3b83b8894ee87a6556be3db5baba16d9ebd2ae48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186e3db5681aef17710efd7dac4d221fa9a11fb48e16705efa3a096cccf8a3c363907307d5232fefcd5db5257ec4aeb32083cc2e687936c8d283dbe1084fc5428a9a4f26886768a0c42aaf170cf2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcd6ecc30001ece04232269cf3f06da3961c6f913087efb979092dd7cd051757a4c293786f5aa531e07143fd4160c18e41b83c97dd0b9ff8d12076b1d1476b8b5581c1cc3ac9ef4b549d9f39daa0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21054b4eb2c6f0d9bc05178ddd65916010d888dde50e0d3ceb5679ac5eb7fb33a0e9307d91797e640bfc8e415bc1c840dca822a6e4ce76c107fe42cba6cf5171b465c408ccce2cf7c39d84e97a27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b23bbf82224e36ccc80501903c6b1b2330499b1e0b6f0dd6ca3a1a20149896aa588b8eea51fbd2884504c360fb688bbcb302aa0dbc355119985a38b6ab5ef1768a0ab87cd4b2db37c6b8201ad8da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ff965cabf3a9ba28f0171841eccf47a92a5739319d0d37bd6d8f3127ce820f58dec33361391b11bbc5ed177c987f39ddeed46ced7bcc293273353969dc3fe36fcc86701626a2d7722523b8ade1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11766ec95b6b4c801638b9acf70058b0a9be8dd998d80e91340caca567b0899971bb776b8d82e1f035689118a5df905d81aa4fde7e623f1e1792263b00b7d756d3ac49364b1d2f5adfbeb6bf9c8e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h262ed394ae2d2fecd2f44d41e53619530f9d3c82c05037003184d02400cfd77f4e9d66cef8ed1133d6bf9c6ea71cac82063c11832dd416074d675b81ab077da35ff64ae0e0ba8faf32f5a5842f7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc83ec295b13242248804c718416dd252de54a93760bf254b98a344d388726919ded998c44866c2d837059ef7878baef854e4ffcda2b4d4bc2b13089a0fb79318b5da7b769b9a55365832bced256;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4656577d28b670538d6110dbb1de4115ed86ef6c99b810b79ef011c780a3ffb4716e05b58376fe68003a5cfcea6da613cb6f1b936e190dc177cc5aad7fbc0c5b7d290d48b81ebb5a8c46bf2b17e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc210793d212b58657bc9b9a29f8fc68ff008984bc495bede69508b3bf1a644337b3dfa91b641ac7f878795312371cc76584a878bb1748133f81301cb1ec2fc7b11c92c3340d2d1daadbe3bbdda6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3025307330101f38cb95dc20d82bc64ab1eb82a7145f5787104ffa06ebc209f1478327e2cd9afe538c60eb99f741b424c3ec66dfac846bc11e23b9b9c972284a20f010f35b9a61573e35ab54920;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ee34a2d94e3a3b963422933f576d6549737baa21d9615356b20fce530b0d9cb7a7ad3d9ceba7d93d1c87e2a623b9408e9b671c0846bc5193964f34557b4b39dea20b1408f37b5f151c5ed08882f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118256c2fae93d38a205cf4ccf62d4e91959bd97ccae2f497a22eab3fe5f17a61a217589317d6033028fe49503c06f60c6c5daf72d7773f2acf6542c765de8bb6e041d056d589b7c6411c26064db0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5365d1fa988c1f27f3fa5176af2fcc15c1164ff4a45f7855b1042a181ade309680951217589e5df3121945554f9857a75c78dd0b4d3a12c7c93df63fe9b7ee1967fb6e6876d378631d5c758ea9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5b14778cb64091e8dd31388242afc277b7b4ab90c108bf47aa2effc63c2dd95a3faff02c6fced0d9b807dea1d42a45bda4f4e77e2b843e2df9e2ba63a763c21ba68c3fdbc8a606b23b87bd0602a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7b634de15e1b30be8f04e90be9cbfddcf4976f4a7308dd0d2df35cae139cd4581aad1799f5dd087e0e09e8a211bb3bd5c687a34dcd26d877b7751ad28ddd5539f41ded44d550647cf555cbcc982;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15997d7587ab284859d9bd42dd127640a4078d57d58c73f7d476f9081a7d36ed74c40574fbc49ef1fe46d8299800a72fb6bf8ae41704139c079720d3c08c7369ed139cf2717daf3175a02d0b9f8ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1837533bb22d9d2bb9bb9d439cca9c298fa7a8ba3b91887de53a4d572063221ec5ca4bc3c69a2bc77311a92b0d1f822454359369e80138f3754de57bd8f46498599559ae04dfe34c9b4c21039ecb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1d81ed87e92d3acf15deee7394b8aadfc7eff1915cba836cd7fbede5997e01da483610bd6de89d9cb4c00964fd7d07e66789523dcca88cc87f73639b06edf5daeb1e7f20c0ed4c7d1b20acdde36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e77115015ba1d11629ad1e390f36ddbb51e7330d6919b8c5a34682637c9582a393f75e5e19c7576ef685e5b831f90cf6a6be176129fe7f5f10203ad700f613e94c97cf739b57891db466c359d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47dcd6ebcd9a24e1e35f0deb93e97fa0ed0a5ba99d680fc5efd98cb25588c444caa9b9f6202a27be62c71c7e9d80e67a51ded58dcafa1bd8d7b4149d2975e767cff14234f41695a66af4ee7f22d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14abfce7fdc5198dbf6fb7bd2e22a2c0ff42546894125fe818dd17753aaa98073df998990ff2c7d22a11f07c1d92680dfac80923699e2d5af5bdd1c0a6909dbeb31e637d72be9caddbdea6491b882;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1231e8ed4a0e48a2f65e089032781036d5edd3d969502c34c9b64bb85ac5a50fa7e7570cf466afe51e25d76f7e689f2ada212ba46f7ab2541bd4e52111db91a1fad30917fee26914217b48c3f2951;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a352973d76d200ab684b4503be492371e9453b7ac16d4a198dcdb9c1e7be89b321742cd6ee1232d19874cd018dfbc4b162a19cda8c496767992690dc6ce144931ae72750d05b29bbad886b35eea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36d567fe65e39782d4df3ed2f1d9a44ad1ddf3afd35251fd6bd6430751e15ca4a60f610dffb604031a87516c01c720a69eb5708c8159afffd972eaa430e94ba2e0a870c6afb6767dd693b659effa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dffec5c2ca5d474fb6ec7ef136b045e9347212492f912887c3dfe243274bd3b3c6c94c1197d3b1d2bc99f25eb68f1be35426d77fa1c2b935f198b6427bb176b33a01c1f3218f5351e14e22bc566f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb36d8f30bf8a2d46887e8bc0ae0a4004b57d5f4f208ba25f4112f408b7eb450885a4f236f22f421072b8190d6d31cb7fb348ebb12cb82aad49163aa293595c728e3f5ee689a2e662f1141f76c224;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5796d950091522b84f4cca12a22efb371e18b968c79e0bc001db57f53ef718caa4ea96c7565b524818c4530576b141154001843810d924aece96581574d414f80c5f6daa0f6460257e2773f379af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c8044a7fd4227e57396b72b1dd8210ebeb3a508228443af75fa4e211148f6700bf9952d1fc631555ad886b30064f82086c7e32cd92ff185c8e2adeed644fbe521fc8f0d0818724971b3e6015316;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125323f84b7fa964d76947d0643afe47fe73278724f648b7a5697985dd894952ed515aba08878466caffcccd04e175314aa42c1efb1ac8f6e913ae12558a54334be277a076b57566cb68e230d271f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e504ab4813c247a2358737a6adff95c73b5506842202e876e6097ebbc2a64bbb7f0cd52395870e3e7ecf744eda6fd76dd7f87e82c180150b11e2789c8aed23a11b159867138d7221f7b64885d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1876b288e0d8fbfc85b9d214f59142309f78bb3545f6278d64ae6b4e36dd0fedf7179f7c30bfb87b4cc4b280ac264465f1100345315169de8d8bc553434c1d2519b86637ac135b140f7aa6d2e9c57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h424f4e8e302027a68e6e9a7b841edfbfd392411fdbf7c473bf24eb5f7613e1bcb7b430de32e15e62eaef50458b5b1362938a6f9ffbeeb57b763ce3550a86cc007bf640ab5d103fd7988392d4d543;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d612744a5dfc36f6c1a3f72150e8a293de792761c55671ca1622aee02320a3e9f56d157ad4f0cdd0ece9f9a9c6bdf298192394ed8bbb1e9bb42ebb10879c9fb33555f859eb3b76c53fc367fd4658;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1096b091910eb849010a6a1a1a6a994a3812c0119e17808a9c39af6909d5dd8f5ca754d3615dc26a7f2290935c5963d74dbcfa6f4e21783139758baed347f5afcc43112399bc120c0fc3f61618c5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5e34ae8819d84bb8e2bcdd097aaa6e5d86e57f6bde94c2a303f5909dbc67bafa3520bc55f09627d2dcd447c9d7e2c6871ee02f36223821ec04b70f17f96f96dfeb4569315d4bc65d97ed9d8eda7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1877af9c5675d2c6bc3dc021d34ad32dd4f0f82b0d4405285cdaddcbf2f64d76eaffe4af2520c7d9e7c42edf07ffe30cec8b1623e9e3d4291e8aa0a293a71d2f8db90578269674ad9e413b8b362d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc53a02955164ec53f21f7de915252ff0c7395713ede59de4ae70ed8b88d5eaaa0998b5596254dc4862fc89ee0b0c190a0d80c497d1acfce622c6cbc0f77da2d82135dd212790f0a459d7f96450a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebf0a7644d02d5f8f124d29f40c08d58eacf054b8c8fb3dd29de270c63edf31ac8ab7910dc61fef83008c0aac8d6e8f75fd513824913d780faaf330e5dfb10669df3e722eaa94ba155f1ee048e49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fecc896837133786d9a9e65f41ff03870eef4d4070b70012916e87fb1df9afbf39779afb6f91f688e24e658eecce9ddfd0a6fc0b176e3aad757a1a0addf07a5dd3d3aec6c8cce1cac1b76002554a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c92f0d3fcd6ba313286cc94d3091a89abefb59a850e533e44a6666a2dafbcdd31c29ba154cbbf249f91aed949c736ddc6b0353383cba424f6eed895a3214d23b0f6f77b732977bf47cc068d4f66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79e85cc4ad4543246d391ff1abd19dbb7022278f760c7ebeaa9b2de96fc9187824b86d79475e6f99f4d8767f841b4271c81d9c3d5b422fb666ea3cbfdce220a359f7e1074b2fda522fd750fb47ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be5ad749a049694e4006960ab3253561c1a7b6844f99d9efff183a8ccab3ce663712a8159569ea5fd83a79ba0455a4f3a232182c09754ef23e1fdd96086f80686f31329564dce72b504115789834;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121fd0173ade6a58aec784a5e42b6c7db42f85006f22780965d85dbe5a10eb98cd9160920b94022c5b721993fd99bc17b4d52cfcee665fbc517808aeb002b508185c8dc7c207523ce163d950320d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e15fd0031c1066398092f1b9dc7b7bf5160c63de70edb50e96433049dabbdf0ac7767ba63642f03e5a0d904772e63e688ee9401dd4b4c6d2baae158d03fafc4a3d09346b6655b1557021e216dc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bcb7e17f2fa335fa545e89afab3c6c944badac76f1914377561d0dc706704e3b7e751590166f4fb7a88e04b998df6bef602970d133245d2fb7fcd0855aa231dba31d6691309ba0868fd9c26d8f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfe901cc4701c63a49172bdb53960d769fe03b5210219519ea23940bdc28db1fd5a9d5e27f38c6b0ab22be73e4ef8478f01117f7fcf25690e30d03db5a9bb0a919683fdab602bb51b59efdf654b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d59a0531503d667e8df2312ba6b446085b32d23a77854c16aac6a748642ab149f6f9c57593dc2e75e94b35fca8535aeb436e39d82a809c2e86a5b537b32c44308125a817dc2d065fab737d5d3666;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcf036f524681fd84f109dcb37fb62316d1f87fb2c59eb1c98aaaded1e48806b9d93726659246fc12070f23f5e6b1cce920793872c0b55d5d89cf3fc505f761d14308f8a47b72d2b6ed48a6f1d65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81cb231a1e920c85e8a3e6d29a72f65303c3855445618f983b2d37a15bdd1886c3c02ad21c20af69954fd16075ef17ebefc7ec1c373d6b4332765b6446a8eadaba0f8cc9f19f52460b5ba2406c90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97903feb8b6ceca25d749d3d930349d21a203465808f3b6c074ef4321dd9828b9b5d954232983918309008dc4b5553100417bfca3091515a26769994b1b35a26939ec918a4a2525c4b4af0d427ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7f1b6d1b0b1dc4ce100423fc1db067d8aa58875211687b9b41f73496e299726081730c6cf72d52afe6fbe885c5be37463bf850c9ee193739ce5bc4d1b1b1f3c05520275db3e54ebefbeefd84111;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb16d7527d48c4515987b9d41ae4f543a39a452adb3b3c36fe71d62f893d6f3c7cc76a0ba8b63123723a2a5318673ba4433e12c4da28a672a9400e2440d7168b9342ea3eaefd078a2e06bb6032c09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e425973219cd682603269c205d73f0c304e564cecd52842147d0839e14cc035f271729afb0733032b1dd933de96ab86989a08cddd374abc42f3c0d75b630d0f533a7a10ba13e3e6b15abec4a127;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31e597aa3199d39651df222dbff11907ef6813d4b661f054c4d8ee3504c1a89105deabfbe36934e1fa4e1da2e45904c46311f76f6ba390d43e9f49f3d45c5096148fedfe73234b27f15f2a4baff7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb2c8dc4c684ab59c51bd5b7336f463740b8333bb37168de7dff19aa5a5c2cb1d60df5a289ee1774cc4bd3fade6b1609617c8a2b6818510216aa0a218f7ae4184bc6b95e457f108af1e70ce7a53e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h700ac1a8600e12388947bd3a2e8c885e23705c20bc8085d8e43af82636c23cd85f8e99355c7874bbed09cb2a0666072539a68a863eb26cdd5cde1d25459bfdb9102d30bdf6a53c56b38662139688;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1966f2c86a39350941884973ad4822cd1f3dbc40ea23d37f2cf3d30186623ec83dc48a90117f2667271ee8df63ac674d50a9e1714f204bb11835b05e67964f9d4c703e767800e06c6381042cf09fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ad77356ff5b24f88d6b280951913054ebc5d584b64aab84db7b8aa8cf8dd2a422b2ba4c641ec1edb29265264021a9ad9508763713bf2154573206a3dbc7f1a1689bb796fce8648a632e4da2e14e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdbe4c15854252aac3520dd6de3c1d3907440705f3ba8c07d05f172aed7807552df62c01bac602695ec8b9cdf93db0b4e3292b328670eb176ac2017b73fae7235e05b9723c007895486bb5ac1d7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8fc021b15ab4075322609142c83ba713ef5267185c6bbd26eea8d056a6b49ed27cba559b3a2a6959979f61a7bab39237244c691d5e3b7ed20143bd31d50daabdcd11f5c1ef1daaba913bb6c8435c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbd042591c82238938b06ef7f83228473442622825e55b381b81cdd01f9e56075efcc071a890a42e88b04d6cacc6b80436b0095108970041c2cb400c68ff07475bea63242fb0384fdfd97087bf7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe78e8b915346c1d8b6115823cabbc6048a764f61be2df5a058ff066a1fa3f77f55d867403c97b6a3b847c93cb2dc4adab5fa2b5a91ca226f823931761247a10efcfcff3998a990287147f329816;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a27b7abcfa3df5e19969af9475ab81234003655d154afe8dd1518dc6882b6417998fe3329fde8b431872504f29210aad9c7d9f5242a24845a8bac054dc7665d7d75648b0f69e5dbd84e7155dbca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26290d7fa357c8d7917c95e176f769532c72a4b835976ea54a04b5000eaa57e076f437650b944ed4d28e308c377985a817f7b7e16f276cc1bc77561c2b1baaa144f16e6f7687e86f85a588b6bb37;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de526f15bc5e537f96e9c7bc7683a7a30ff5118285f0416f7280f0dbbb1203b48d3ecf65bbdb7537e369fc85083817dbfff1a4ab325961d60adbfb697da23ca94650d090a44c75da20f570afef6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dafc9f8dfae98347eaf51cda343813f92367fe92c8cdb5bf0bc4458a5f8f43807cde171d642cd9f5def106fb765017e30c32f41119543c5d627428904cbdb02ffa4a6f9c599dc662816a7ac24fc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e7672402e359616d8de70dccafaa7d191345f1c033735944cad30815d97c1ccf1b017a2427e2fb6ebf29da9da838dab92278e6962c209d493e9e281162cfac08178272c95ba2eecc7f269a27fd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76543c333205aaf3ed787bf00124d179e63abfa1b59a4e2be4d2e0ec42d76d4f14c652c76fd5a3da9892342f9f1c7ea4c49dd2c4103cb75c6962f2e9c2414b8bf47768c14b2e944d016fbe8e5cc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4dcae657fbf5f41b44cf9bf611fe5b2bd9a380685bc4fcda24941b7fc8d6be7c32dfdaaf19a1dbf036d491dfd0a80c36ef1a38431113d4d9c2ff8a3a0831b1d5e4ad10be01697cf1794c6eccf0b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95b3274d789ccd293c3d0947c4300af777953882686a7368a6fbcc0225047d409a5cd3b07513eba63e1de649a5e87d867890f395569e3a1ff241d3e24cb0cec72de3c3b2bfa13b5bc2f983b56a90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149bd317e3b6fbf0bc660cadbd864c219f378b2512f66c43a6a79e3c7245803b7e7f75c3ffd87ffdfaee6bb15d87acd54544bee4ae383ae6698ca126b13bec5449a6a56f64291a64bf97d64a23398;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0e4d1f56bb1c45aa467087d1658342f91664a0dedaa19a3786a33f8ef3683cfa27afc156ed32d6ce4e3acc6e5d43ae6d0ecf8a3d5a5796997c2edd823b575287c97f810deb442bfad7727c81a84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183dc56a2f0880411c2789d1b888d4f7efb9721a44e557c2f93cee7a21925c6e4459209cdf081f1ccf99c6e611416b36cb8bf7becf44235508b3b42cadaae0393f5fa9ddacebcc0ec9c141486762;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140a48e2c716e70f97c8eeb736dd5f5ad287ba20f8b06b344547bb71ebfbd0656985a7d2f3b7d057388240449c6c5cbde7ab8f48ee10ecb26c56d656c459911a1b06d47892e5a1129d853cc45e5b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1180866a131d497b9ea90e8835791818e56e4df23ee167b0256727917131c7e7ee2bdad79ba617051da221809e38a4c0bf3dd3ef2d6c6e34023c026d085801b8a816de491e9f18ccf30b967b9c9c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcadf06147c91fda5bf33d2beeb8d111e8708f780efd3c6a99ac76f820944706d0665780c71a3195a3dcd704457d51b506f10fa489b4598131ecf46d3517235ff5a662d2a3c820df8f6bb59100338;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h615c78255d38ca539e708b2e4ebcab9079d4376f896aad6a5ec4af2e1ef0a89ce02f31451ea952b0ac50c304b81d1a59fc20d154fbdeff279f7d3f4693b6f4ff1157d7829acb2363e22691a67b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe486793848c5d87c550c8e7ea6982413c4a84c5000547b1287396ff656a130e67a2187f1bb457841a791fdc3d88f275113f1bddc1f37d943c1dc92b4c11b45013c8f8254f7d3aa54445755bc519;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d898bf734f67915a61b61250a409634e98fb7877d258586b8e384cf8c74176f725e8ee5a3398eb209e25660393e9365e8bed615b066e2e1870d1e7c201bf45528a42ef5d8bdba66adc9722b14766;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb76925d6e0ff7209f516114c0e7bd0ec90c8d2917ad69649bde0444219748d1365dafbcd07a6e3a0868d1b1a7d32f6de4905ad9b7aa626ba3520e552dec5fabd6f000d8eb7bb617331633976d9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e31a8906288da1c42e112cfbf0431dd2acd0ce8a61700629ea07ad33355519cc1faef27461e84d099e68de0e1fae474cde51f03f9848390ac712c1801065709198ae5b714e6a06591fbf4322ac6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e5cb7487978d6b11e9f5c05165b7ed9201df8af15e9fda3e9c5b1342056c5ba1032569db587e897e2690a787b66daf2957b9a958a51c200b3c3141b7938765d7943c179a1530d38d683f7ca9243;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193010f821aaa16563117778538b600129f0a68b939f9ee409b97c54c7d5eaf6c1877875f66190687554749f492eeb6592be6102fbbb87ec1c885a65aaf06584a916503f430feb77065f859838dc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6afd8a07465feb4b32059e956b592e41bbe889dc934de2fca56770c038e60b6a5892814ca21b64e8bb53ec13ee25f8312a0efcf06dd98fb8b92737565ace722cf4171cf2c83438489fe9d416816d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12119975342223115a08ca91a28a518c1588c2e0ba820a3b5b5761915d628408a52e97fa9f05f99269c235972916f8f21a48da47d75ac2d67449ae0e42a7d92893484a3a135139d17c5f1a2560c2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5f3853bf05a61c4e9b52b6ba654416f2a051361a696fa1190eddc5315844cd0797760f2fc6d3324ad7dc98e6cf2c7a85011f64645457193ba522ffef6293a53e11584c4285665fbf77153b94a04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc694d3e2d5e6ab6adcf4951a36557452ad6790f9dd096e4167992d301d4e2b89cecd590b6fab5af21a5b6ad77ba4cf452bb109d49ec6e699ca627e41a4747c8fb43547fd3a4d091744c7ee762e8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d481e26643ad35918167951ec2442de3f34d71b7f42997a3524a56d9ececfc281ed025adf82fecab519f40681f1c7ae6add7178a090a1dbbb43b22d0e7d497a6f87d01e1997ca95eacd5fc17dfb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf52abdf3282dab075bd20e255d9f44da1f03fd3495b093e3db9f1a13fad42421f53ebae2290d1ce849ba9c7d2721eb11e5ba269b196b338161a7cd7e87e8fabe7c369a95ff188c3fc51837a5274;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a877b37e3a08ed767863922edfc1503e45a36451ddeeddd76c740712428a012fbf59afb8594a1820f044857c932874a965314ac7c2f7d8e25ad470056d450a1c96e7233ba1f93331e2554746cd11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1485857fe70e97230d09cc13f2a3cfdf2b24d3a3f5f05a4d808bafb969b15cbaef2128dfe5ce10b2d96cd80d30d638d352bd71f4408fb5729cfb1cf42564c1d9a1610002117ce0e5de6b4500ac179;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb720bb10d1e191e4125bfb57aaad6f343418a2b890e9e7ca45f6e8c68731c17822978bd03a16c5ac1f96f91052510a7db88e6c62c13257bc7ac07716fd1af68fcae58ceeb9361de46dbcee7e5c7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f39e896d1a886820bd1a58beee27de38356a8a96dcdf0470f76656be76e5d5d245ec5d33d26a626e9265bdd6ba7b6a945d925cd361a0add874a719c7d464f76437cfed1ac517e5d5ebc87e3047a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b3d855627aa2013b5e223e462c6f3fdcb98cfae1e0aadff1a9e65326a6c4985dd8aeff04b35a12261119e9e98c7633a8b963e57775c3a46f6a57c6826ebe8b4a6599497eb904bab1a5bdaadb467;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b248b7c179f28f08b28ada19359beda25598b7c0d3905a83d3971f21d7a254cb995a8730b9a182673af486585f0013d39ff89ec80d3718e36113dc64d5e664bda40d843ef94ef5b11cad6a5bf80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1888299ce7c4ff883dc145f4f4d699c936048d1d8dcd29aeba92c7aa92b4b0e93f34bc80836c904cd7a665345a3a4b8c6631217a76951766dbb4312c2b94a236f0284a54f5f81f213265c42024000;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d5ca06c66f6301e26fc99d435d0583ef470f53d8aa1b679e10938dab0fb438360774ece6565a8c1855879b3785f90674388ccb293b6d02c14461cd371227c9f5f569b4ca6628d6bb2990d897265;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb3cff527258a57c269fb9d6301850bc191824c5141ccb95f25f5a2379550e32a41fbe9a4881f38736bb1116d4baf48f12fb6263b828155a2550dbf9b5e6cf392911a659336a9e97a6975dd3fb3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb0543648a983f95d4bb4f27dabebca405ad84642a8faaa3407b5b0bc21b6f9b55666c68233640a8dd82a1ea7cf0fa72e3cf012d42aefb06d5607c651c9f618bdaabb9c1dccbc9719a7386e1494;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d53e847d908dd7cfe73867bdbd4b2634fc52e9c528307ff47bea4d8fc996b1307c7e01aec1be9c79fa4630df566f39f0cf638154fca6af994eb66a8ec02fa56cc25f2bbea0b660ea0f79c2fc38d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94940c5be70a0b7eebec5d6635e0c0116f99f1f111a1c7a3d6919bb28b7e3e19fb1278599bdd238c707c4db2b66fabae69bf56099e9ecfe3df5577fb6e98c33dcb34b404e985a8356820e6dfaee8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce955f801db2fc9bf10ca730a0645a47c065ab5f5230311aa6aca738c12e5419161130bd2c75ed99f53d2eebad00914e7c1891e64563234dfc1da2931e9bc994cf528a91422e0657d2b7641d7ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h403ea5e6751766b1ca46e53b79ab0a9a6bdcc994a4d43d1d6ff808ee923557f6bb0a651bd1f8b70fb17c687220c04081b070747d91dac7c08c67548a925a4f9a01167ce291745832b2816d2c106b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1f84f2b123ea0eff8b10aa11005de3f6dae21ba618403cb5bc60171c65178a85b264e04c8d2831ce896269f201db6181f0426e98e45a7e57f2c266bc33d59b61f5bc8922c7fd4f2b7e4816afe23;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2005516028f6bc6727e1682f8a6768b6e4619dfa8cba6e7c98952d1db22d09e261e09c83dc3e78ac2cc9a020b705bd5a0cca2f0b73ebb63170cba267e7ef5ed8be265e4191fec216796be2604f60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c9035c98cdab2d8c4138fcbe2f52e635719c5c44a44a735056c9b1e222ee05588bb38f522bc53b150055dc1c8b0a70bc5abed7ef08e1ec24d13363eb324dd820fc8063d60fdf67815f2afe83802;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e0cb54e8b8deac90064a0597bf891e2b92b732edc9be9a96e9e997b5d7a977ee1316bae6c6d5876752726307cac98c7d7f2e9e5b761ec5d01cfcf655289b8b6f584a13f03fe56790d412b24fc52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h630a5d05fc63cd89fecb3ba1f819537a1bc33fff471a5fe848558df24ab67dd29943c300b30e91ec50cd98b5f25c0f4a304050cf9947a5d962f1d41cfbad3d04b4ba84a37b791513418a91011bdb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1c9c4eb576312c74002109167cf1439fb032dab7eb307762238628a9bac5c8d9acbe48e226472a38a7f7cccf002c41ff2a43f97af40ee1e62f80bc54275e2c9c74b031279831163a644a619d5c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha701472f6a9b50a8ee6e79708946f4f6c7d905e4dd5657a16afb77c34206ac42701813940ca3027b8653e03d031c01e53b1709a5b55b340928c01c7886081cd986659b6e8dff892ae80fc92e6ec7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5a242a6145aa7a6bc3a4b1fa8a26d4682deb33efc3142cb65a27b1b8fba835f926a7755d09f395a8d399c5aed5dd0c433fff2aa1a44279f97d87cdc44f22f13a819de11c5623c90cb8216f30156;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e6dcd4d074ed6f1f9d67a38174694b717ecf44ad06e8898f005b55aee3c3cb0f5bd9b1844b00f3547ce1e7ca5f53b6a0bbaf67d8339616e8efc9efc94c66f2ca89b2f19c98efd96b8e75162b336;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3df3b24d791e0d0621decf593bbcc5913b40f5cf7e85653ab03d9477a16f76414d528f3468bcfb2484f574bed1c95858ad6161123444d1c12f7897c80d1bb31d819e327cb0571c55972e1a49cc75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17298d18904fe1740598fa65802de96cd564ceb2bb3d20fd56a8f1ec9481b81d49dd684ad1afa3727a3ac9fc49ee6e7f0da0726b5e20744e580609276373124d74c44dbd30edf555d9bf22d029323;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17377eb013e832e5fa0dcf9e7962893a704bddac72ec56a5b84b4e6f615e5fcd6ed1f7f47069a681296825eb1f11b1ed9d4a4e258185535c288e311c7c05070e3fff94fad09a0b28b6ecc63f17f25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f70d96d297fa692a312040d95bb4c8b9bf3bfe1ad29c714b79c1617619b08ddc5802d0c43e0a9eadff23e1559ddafea7f341701652c3a8ba65645fd9037001a694eddac1df7b6977d8473be4c8d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137931a7aa28dea28c43dd63f216710035e19b3e4dd7bf696dc2f88eaa41e5304a70ad1756071574a2f243209752510f6b14b92961a5b0e5f72b7f39c4c405d7fd3dd13f07f9a0ce12511b131fe40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb324363693090a2896f1b2ac1bac4298d2135601c0b45aa099c960b21f6c1db15b577ed6c94b5448141782c1bccd7c47a61bc9531d7fd62aedc3671e8ee2cbc2f7a531f1255cc00ebab597738e4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb103aaf9822daee49bef8fee9f19d947c41588d928910ae3e7d219eb16feb5ca22c7c1b1cc4ccbec7303c136a102ba778a1c44427a6c2842f9f0ff9f983394196be762ea4e49f06d98c7c1f66f83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0e858bcdc6ce81f71c071167c8d3db3b124ec38ddac1f0f06e08d19f905d24a236299f5c5c66142baf9f66e6289b270037ec4d6640c76947979f17dad70725ac519825f9044f7d946fe50f4d16f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfddbfa0cd53ff99255a88dcf4461ce4d3ec2d65be2476b1dd0c2c7b9fe7c0eff97aba69b91baa7319b56259967d3383fea4b4dd7391f59f0abc4eaa78d61403b70455e5fdcb29a3d570d7d665ce1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1474193b171883ac9ae09f86f43c72d4fea635d2c55b1618bdc2cb3c659bb227cfc4e65929220be42c6f406da47bed31b62c6ca6dedd88dc3d751defb10fbe409a09cd5eb2f28b86e937726e1fd04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h633c632d2a1a7cadec5f4e61f68e70674f028540c615f4573e4c25b956b8be9471377fefce849914539800a37dfe75dd3ba5abced5d6f87af1c694d51a2aebcd48731afc34144f848e9d236af503;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bab32d378dac3f09a92e841d9b6fba4f88988b08d41a11d443a405fa31b17bde30144e7b9d03883c0b1e3d96418cc4c2bbd77e389c019705465ed14a5edc5335e3a72cc652ea4a78e3217ded143;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7483197c8c0e9bbdc37eca43213c165ebaac45a811b564c30a448c7cd737bed2c6ccea431ce0bab27d2292aec6fa30772773776613862b0528c3a8c7409f1dbf27f410af03c2c593deafe7fe67e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e33218afbfd5952829304a854bd7a266e58dd6715a490c2868299c721c3a80e25996afe2efc290e18e562fd799939ebe5bc1ff262982be9023aa8d117ddd70b9169bc1c81da1442bb60a8eb2a039;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7f825b9627f2b47638b687b5a9872d837377268ea0c95add813d84dc4e14dedd180003c63d7552c1c4173ab7471fe39f2cb278609bf6052b5887744e13248aa929889e20a29466fcb3feb631961;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42ebe761a33e3ec688e70e101f156af34b27c7e23c8a25bc2535127d85f19636a0e92bc6728ecd0a4d692989164d42852d6c1a81da928ef046cd016b88413d0c4a865a967fcb156e8cfd58a8894f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h270a56ddf4dee3c7509786b45be833eb44c9180f1543e87e2659e339e4d9773620d8a6be587519e35791de5ad24d521d94f9ed44e37e620e58b133a5b611e084262309e2c752889a18c1d2c3c1da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36231c9fdcdee10453612515704900b1e313e519553c430814eb2395ed42f96a902a04bdf015a6b99968582c7db353add0c5e2845916f543846cf79385b5a9f5d833fdbd1c8057c722451fe1b137;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92a1b18b7c793b527825f96f46bd4b305947312c44ae53cc32dc65e99b4a257e7a952af676c68f05de3291ac4831f8c358456720e5acec89686f120039e6d512a4a34912ec88f89b4ffe10681fc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5236d9eb55bef30b0511de443e9107245f0bc8409e62c90d8f57f8a20bd20a1962b592b4339b3b17a2b0261d7ddc189d18c3c01fe1baec32ccfacbaa2ef2eddd24f3bf7e25650e6ca79b1682d64c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e7fdd914e6f26cf00de7f3cd2e11d82ba6f1544872c053a61bf36afeaf468ea48711bb14b2ab8ba79bf5eb99ae0a7efa4a2400f8684ecad5babe163eec508f1b55f18ea60090b3444eada22d70a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4d00e8407dd7bbaf689c7bc015c6a9bc1238acdc71356025cf4dbd2090ae88d1674dbc08101da5dc22836b5f2ac63a2619e48e5202ecdb8103b4fda85dde6cfa9b3ad1b592b03b019f00af4ce4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163b4b16fc525b2fbf35bcb607303315043dbde1388947b2f940656c5110224a3a704bccdf6f3fa7a7dec26d9dc74b201447e7aba0a28424ba713599f17e6484cc31d5a7692da1e50822326ef00b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e6cc9e3afcfb0cff0f24cf5ad49611d38c68947cc5c01fe3140158995dac09d1703ecb939906b8661da98d5ca24680153789d855783605fc0703335f901116e96aa21577622edd54999ab4f9bc3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb723ef3c527c6becdc27186e28e85b5a1c193cd8f449b782b3165960e29b1d5d8c0dcd9a64ee54030284d5c7b0759980b6dcbf82ad64fde13702a888f12161a2b81ee05634cb20a7b6ee1f9a207;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13413d1f3b58cecf29d82e0bb66f395a32c558630c223634272d5e638cb9dbb38040e2314b492f714557293bd3906489bbffb99d4622d6c99fdea538483f6513a7e9cd507747608f05e819a49cf1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7732107449af8d37b49e4bd1c3178c49b59fc146ac212ecfd8adce9e6b9b1fbae7d338b8c693935dcdd14e7d174e8f061814d1e19f59c662ce8ebcccf20063735cd892bd7b27da31896a5c055ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142e046bd352480e1b779afbf3f8e155eb7c2c617b951613e292e7dcaf11e4cf8ba353f18a4267ece91a6c38fb482451a4015c69caba751dc2e0a7208091fef9cb713069f183aef222ad25d0f6560;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa5a7c9ae7c147751a45c616f9c6890b12f9a0a6ad7e325f067db39420a3ef638dd84720b3180369d301c82f81e4e5c42284cfb3668cec511cef8cdb38a54823e2cd5a5ff560269736f672bc67f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102381f1d5afb6228f85cf795ce1c28092768636ed2e6d25caea33b0196bff252676d649d7fa40309edaefecdac3de51def1eafa55d3f386840aab8f042238a1808f76bcda6e83fd1fba674827dca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6fad7f2dc0a8ccc37c635c6a45ca3eb805dde5b41f59e69c0a91fdce730e5e57961afeb242bec8ffb9decc1c05571932200fab7531c00fb34256d3b57116ebf1a222aa401e43ce1b5d7e1608feb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130aaca8600ee1db16f9ccc8adb65cea0ffb40aa71071613cc54907257d48c8db3001fad3848ed11773c60879084ff314d223f3d67ab9bf9c0757000c8e7662f8ea118fd6703de42141fde10a9530;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f178f6c82f9c9e81f5628c35ec3d5b9c576295edc9e5cc989aee567ea92ccf4283d7f90221524a08b604ec00b4bfdc8ae5728812d4a7008c57d8fc633d84489d7081bfd6b0e95a778bbd917b0bf7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22ddd8b462fd4dbefde28b97fe10960ee7af8ccc033737f813848eccaefcf0c2dc22a20caa57ae1b06d2323ea4b0dcdd55986604cb58ec470e800dc808529c531e9de07dadf2cdfa3fc61accb500;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df26b917d7f0792a7309aab2efdc31982755d2faf82613b273aca7fd60d16c5f60f51776fe865f60679635b28a718f8411f57007f8dfa6dafbe3b4478e5819fba503b17692d49fee0b9350b9a876;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1461944c38792524682f91934dbfb4bf6f6adc9ef752fc62f140dc0da52f543e44a419f0ef2faa1fcb4275208e90d7582bb87f8aae5d50b42de52b76b584eb21965456deecb1b7bcbe9cc34b13c83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha542a0a22526f9a928e674c9873993fe6ec71ceff514f797ee903e0aa6eb77508cf872f2e7e44d28353b1228989b250180ea4619ed92426c5792880d0c86ebd85999427f6aeb6682bc8fe669f48c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112aba68f178bdd7a157f74c00584903374fb4a74de285e09103bf5324d4066bcb7f2ea6ea671782049d4bab0829378c548d2b09412c3840d1f2d2794af1090a62e7f13f5d70e6baa5077ce29f360;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b1bdc7c325d5e8706aa90c6b8fd4f05ca9539c944cc60827f20b23f0a443f16abc75ac1ac420234ef4ecbf5f74c13c03f21ac6afda9fe92f4802687fe219dcb9677310cd174191d06a52c8b7532;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha45acfaf59c03b9a92b32272e5e661139dd9bf4bf067454c05e3797200036eaef90c7aa2c59d06c0df4c057ba7a8303eb5b43ea516e70b2f436e35eaac7ea25e40ae6db9dc1254630739121972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17eb7d3bbb9e9080bcc0a04b2a5d6eafb29b4d9017218712f798b94e737b60431bacae14ee2f51157891c1fab1a5304beed369115f21f9f45e2c62ff5b6a3ad6c38ea3f6368bede56a3639c063d6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha39687a0154c19052378e94f95064549636f0d9f3109cdc313d4cad5913c411c08bab9b71a17f912f70e266827a0db9535d1c1b0de755f6ea7e53d58a2e065a7fa8396874dc0f59fa6526527a43c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27e00e723a392c98ade8adda62e3b99149963ea101978f27aa0833f2d4ed5a782af1d4c044f9d6cbf31cab75b9e2030203a6eeb796b2e538754a7dc5ee1f704cc9a52b126cb2939856d0c044a072;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124db01520c0149feb556bc0c98f5a83689ffebd63e68d0d4955b6a645a7df01891e34d729afd62533070774bb77563881d1f6a143703e52cf234ecbb837383dba6ed5e009d7b020e969cd1052a06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21bf7086f3dfe0a587499b57978c930c60ac3bd788acea54b49654f63e8e69ae715209f01fcd8a259d60d9a0d02b8de0259f6145e5c286324d74a2a6bc1c25fd6379609e262f396e5565d75d0edd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed06548748cc3de67836829dc2ed088cc385be5a5533496f2104e4f2d3b2c1151e7d84bd89b163c30d177faa1ae1fdc00b5d7f55e96cade415538494828ccd584397e30b73daacdff52d8d04f649;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f59b63186713918a6f452287cb0d8cdc7eb1145a6960be7625d4ab64904ff8edf069ccad3e57298b4e0ab95e8b565fac0c3f4b6baec01356ee214ff51b0e54b08ae58674338ac13f0e5f4b0b845;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5707ed2f934b3d86ecabc31b539d046f9bb72f26abd7c3ee77d892bff7bcd9905129400481b684d852ea9a72160a905621fba0277e1a3f498b12a02d8c1d2978042be4603cb396cd271da6d6a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccbc83eb25223333bfcb848e55cb9f8a15168ee56ccf139c3332cc280d1ea9b1276277a09587bf110abd2308aeecf402cf61f69ee373f54e52c8858d7787f893a63e57ee8cb189688b48a7d31d2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8ac317ed4073a0530d3685483f691aa36c181abf29820f9263849e224acd96648a289f502c88e8bf8dc1592c5d2b24dc853f850553b7cd954810e9f6d930b4f3b6047b06c74f564b77a24869a2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f7c5965f0acbb4bfa7a02c9eb360f27cb0b2afc4466f40ff6aa7c90f38f9c1d13b7b6475f12e5e3cf11dd4e1d761f8813216956c1e4e71a753917216da1341d9eeb1e86a43a596e73d3a140202e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc31f8ca2bf97c57898048d0ba6165c771b889020908a2965aa4b6ba21f1d5833ba535e475b238b7d3c28bca7e3f81a5a62108dddc5369c95e86c8d0048609ce30103742671865054168a40b72eba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a5e0e77ee1b738ea650f0479e889c9c67f801afb7df472d5a1e54fc4b46a54fdff86740771f8847c54e320cfdb64a3b1912c7a1f148ded48e931fc25c0ad458687d1a91ae57723f1a2e2ffc503d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14179df719abdff478982adcfaf246ce9054130880d747f2305d912da4a9de924a8bc41055199a2e8e9a9b0ed4bc14102a8ef2d82d7aa9ad08e12d279f194e56c3f2049a1bba5c76fe8de54099ba3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17aa39b193744461ab4e9d45962bd4ccb27e7ec73b55835ffed5b4cf054597c4988fecb87ba541334c5008a7b6fb37d9772946ce30c383f788111be3f571bfccca6361b3c0ea18c5dea42b4134afd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103e009d21d84f04232e3040c0597c2deb5a76f10a095e136820622088033a2fedb588c7b1cb198113bd0564114b35023c29f9941ac4a89a4df52057de5117aca2c4128dd1a9ce8d41da19b280351;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fd4b178d3604caa5ae35bb9d60c93d6a5aaf61949d7d9c6b0203db854384f2e79e0c3c14befca118d9655c96c5caba196d4255b58b600a46aace5334d3e92ed6cc5f266bae620d2e1ae1c2ffeef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a8d07c7cd6f172a129483b0ad452f85caef886707e691bef6c2a2375bf58e8b88fbfa75799e10d255c573b60b8a2e8f1c6dccefd3dfe7958eb1c759661364bd2029746fb6f98ac475596f6bb219;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca2dd3d0712d4955791ee6508fffb75a853ec0ac52e458f59015091957fd526ecb4735cd646113fb46bd0c1fcc6a84be4adaa0de2ac881733017781d0cdbafda1041ff41365e69fd7ea3792acc49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19273f5d9deff55de6587b7c400b631634d4271678a3eae97075fd70ad0f5b38e4a66187d7bb587e6d4d538c6a4bc423ffa5935ca016db2300cfa11cf236e6be557a1a4dfc3453c15d603362dbe8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7bf13115d960cd87cefc8fb417b48e6060db6ce199e8f3d7657f1f7e04ff818d03a0aca544dd3c086974fe2d0d1b6cd0d5018878589d83b404a1aff5afa5fc1547394cd456d5494e7e0e8ac7932;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5257ec095c0d13524584cc77cf9419b9938d6a9cc5b447106aa7e9e1b8947ec1b3628bb66100da3d09e829351936872c695217b5fedfb58af511f182d9b4fdba913bae657b8dc80d4c23c97621f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c013adf0decceaa064ba29d1d5f840890e94e2fcf68e2f7c18b1f200a7a7df19f9ab288d44e2b85aa2c14903fb9c012a00f9e204a18f498449b52483b8f3b2df6fcd996b27beb342e049ba9f0a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5d3b321f0c958f746ec40e51fed495ef2521c8ff2425d43012ba418cb115401fc61c51bbec58ad57443f2125649828a1e0b6b6f94ed269e45f85ecf3aae40147aff2349b09225c745702ce60041;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f04d25d1b4fe361d4bd2f7c3578604154d16dc2b00656efb1193c5345dc5fd8d543ea7e87092fab989e7f65f61d0a73b9efcb70ac5b16474ad2b744f81fadff6aa8dc218b02d67c759a6c758760;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1213ce5dc546126805a33429d560b95e3d32732f6f429880c0ccf9d0a29ba78c70038042d6f3e22bf3f551de6bd2789f7d6bc49a9065b4bc02f7fcec688a12a8e66eed6b9cb1d009549e011ca7f3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac548f9cb4a52502724b8282bd016655e396f99acfb75fbfde95b7e2d64701eced6b44a6ab5eaf1438d5990f38dae12fbe71ed611230ee3fa3ffd6c98a0da715967bfdbdcf08ed3dc8732a91f6ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165d4669a31ca3ce73f816280e4f89ad4c2490e949d36764f9c7950f24d110db0d27bc9341345d9e9cf5a62cb6a368194617969b6f960a7f5c3d0c38a170d3fe1c774f3c0da032d469b5c9ebb6e1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a330bf6cc1357cd2baeb768bc53e3f380b2b77f9802741724f5227457241f48772ece3f9f4f872726e905684dc8bccd29add8796b0549c7729f7b1a0dbbad89eff49577a8b7f4448d03710d4a619;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2cb8030371ac75199df0b588673e112bfcb17dadcc687d6eb0e4194237bbe72a45ae31a809e75ae3ae474eb88ed594e0778c016a59bd6466316d5f57656d26d576e06377242129b15b5583dc3ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ad50cc3dc2d677bb744a14df370fa81c20dea5003aacd95b58384f54ef9624fd42ff8cae1205760ddc464f7ee2d1125e3a5b7916ca97cf87621094e2132dc78ecde87a2f46a1848a3fd1e08d7c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10489d33aed366064bcc216536e5975ea86111cad1afc3a262d125577f1c4b9582d495d9f2f4ded5d1383f88d4a1c6816caa62b5d56c1d2ef96454cc786e4687990384cc96831fe27639674ec359e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ba7fa8a3f8336899e18dac860ee4b6aa9426bd06391d0875a50c7d9806fb25b0fc81dbfac1a7ae45c674b4650530bda0f7ec51366dd78f3e68288d145a32a9263e76dcd388a00ffe7d6e6a9e93f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0518362d598a7a2ae286be39d89d78aa11bb4e29e08940f3f2d7ec0934d47f79d41247087437668ab1c024cddca4efc1903d37d664ab3802ca45091fc0ebf9dd5059391cd369ab57ddc3773333c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37d2f2addff46b6e5ae0f2e6713e400f1f6e3b302ee432b37ccc29148941a16e18e021fcfbac0ff96264f091c3a3d2132c48704023f81385bf752c9d5958f220a4c6002c7d803cd93718cd244cf2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ee6fdeea2e5a607d6d1ed5752dc6c813093507612a365996b21e5e65760b5f9d378bc0fbb95133ee6f3f8cc5534ebbfd2e838723273563e4d0595b47df798454acc02ef1f7d7b8990241315dc21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd7221e2f1bea1135756cd5ba20c0583b77b63bc6f97d9ea194e0f815957781a657f7b832c876d2b04f7ea1871955062b929827b8e0e26da502672d957b46c028fb2fe558ef43db8bfd7b52019ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3780fcc92dd5ebf24cc3f976240436c9c92aabfcdac843f05af5da253e5cc9686c450466b7207fa1ead7d0c13a5543fef09a9d72ae8e4739e4267f8d53d2106b2377834f3c48350db25fe5bbb74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6d0e5ccaa7573f2184c88e7377bb217b421c83fdf384119cd4f9d0319577be51d2f741399b3afd25bccf8d3e0e0ae913b135dcb6f31b5d368bbeb9508b89c3cbdf587d10a88af773104a384aa9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11211f06971b3fa02074edbec6f0013efe1423b217568725e8c3478fe3e0cc43281c96826175c7b56be779f4ac4ddb5336bc7f1c216a70aaa71862470ffe32f56dd0e9f1e093ca280a64c3fc6a75e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3069e5c28e0d648a9bf3ceb5e117877bd442926c039b417213bba9a855bf405be5471ee989512548848151172e24cd70576266fe43efdb42a3717521e307af0a5e4d11b8b21934a359efab6d25f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ccb345945fd38ee7d70c4545c3e9d086520b8a51801d3e885dfadf07c8129f7fd1271600479fe095c6aaebb9308ca9d6c840d4817e6d318714a66b6c4c405e3a4f8c8ff1f73aeae59218db212df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8a336ccf5d4118ac4db590f4d4253873affff43753505de7060c78f18808488c1574976f825cd541be50a535528cc659ff6697066b257fe5068cc11d07af6cc32969ad652ef5a83c3e5a34e1a03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h932458c7a137556a309f6a98f9404e1245dd1d290a126cf2827228526063276614d2aea0c515b637a868ca50a96d4028ca0c600bf75d865e5b3abc9b6cb406486c0e5dceb325763239ad981519d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcaab87ed99b6b6770c6095e8e8ac7a64cd895dfb637d956e6f77fc2401adc5c699cb19251f0f9fa4c5a623a68374bce5158995698d9eb6e4aa05bd599f78b7430a6c0db603d5928eba9fb22d9c8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c867f49885379cf3a1dda9fef1e25cd63f0c82b7a68c45d2554494ded42bcb7277f7b334ecc37e12f7474ce868afd99e4de3c9a5b34d0d77b6dad652c0ffd411adf559a9c47fd48a6c58ea1868c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc23a7a3086be021507751a0952c2bbf69e0085782d6c5d4e86d514e73589afa1ed70d6ae5a2116f2ee61fcc5d754e4c93862c7893c20294a2d3dc2782e598a73013c6be5fd769f1e2329049351bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2d2d2d2c53a40d46e338ef22d21bc27fd35165fcef70c6344bde54157128cd061671b88d8f35ef35c66ee1b1b315c9f0bb1c2edf04ef622fc448a33f015eac91a85b12542072602705428b37018;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58f4b6484981b667cc39d932903d71e99613460de102a72bb16ed58d3d36500ce252ab821a16f5326881facf157ed3285f1468d6e5b5d1c2012cef713b35a90ee68e86b195e43584936ddfb8a7c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5a63387f267036fd94c6cf7a8ac94c9f591241e0da063b1178e0589fc1d69ce65f82d95d1cec9aa4b91c34fbfcd3e80967c1f7fa3261a7f4bcfb82cf7479c73037b455d767014762474d539d49e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c12a44294f83a4d787ab1341cc258dacaee378766efd60622cc28fbafa6198b790da7c41abfec9fcd83dd9e1715f6d9549554074d47ea3d78bb1c2b42bd066d31a08b63a98b3046d8af1c0b89cab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b65fb0b62b4238e57d54b231a6058d646d987d4dc074242f697996f10e13dcc35a55aada78b33ceea11fe9f77624aeed7261b892f1bb9c4279db1842fdd0e2b34213b0a3973621d2e803ce1573b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2940359464ed14254cada5056c2e5945f3d745b23b6dece5db3ee8cc3e6ee4411244cb393f53f98b9a96bb3521bc54d48a124532b1589408978580ce1b5e00923710e1df4084fdd467c36a7b16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf69f2faf7219eccd0a344597923bbc232f21385b09e0170727238a219ab49e3719f06f14b0c3d056e45facbace55726e291244094427fd4031fd1c597c6300e145743a4834b12e051d6bd9741fd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae537c97c37fb9cef374477f8c8b29c47cb0f4083304a87209a3a019a415f4d2ecd6667085045c18216b2a5a27b600f9acc3d8753c9c5daf7cb4f4a31b60a9f484ccb665958e329e787436bafc3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181b54148b753c17875148e5de6892945902d4e10fb796c21146650c034a9d14ae9e8ebe49f55e09d0fc17b8d4159a7fb2aeda7c32a5930a2a1820cb6dd6888dc537e42ac2f482c021945a3a9b4d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0c3de8b641fd938aac9d4693e01af9adddcb880245d9cf0a34b57e7738b330f0b3094b55201ed15309fa31ae8e7c33d01521d4449610957227299d5b91a653caf9f257058696d77ee36c829ccf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9f93b1a48fcbdcf66ccda6f7eb2501d38ee8e92380f8c4a76f23acc5f5e34a221b7eb77996b03c4408c204cbff51bc0f1d4785c863f25b4aad8174f28ff2107fa2958f93c020deb5cc9e4ab1391;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128fd28b8cf68dc7f180ce7c1164f8f3371f1d0d263dabc83198cebf01eeb5052f02d7f65455b10bca9e28edfc308622834657fcf37bb192062f527c6e3325464834ef3f7a6306648a1809b0660c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15169163824c07788f063e748c1b528052f214b94828e8e908710d805d96933219a983492a28f294539e82efb89cad6e48018f83b85d9804030069fe4a14d6ba8ed0d3c7c13d30f0a8a82a8ed94d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197b9422d4b55e0b61ce4259525eb910026b91db073ce5c52d9139424ed98e8753d8a371d9a3e5723fefeafc458a9913c4b69adb1d59f983524376aed21c163e16437ba9a18192da155ee740d5dbe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196cdde2dc3d37711b12798c4eb5c47c32939689094a125d9f30499dab36997774f144f11ef42faa286e4b2910e589d421ed90256e76441a806e1a20ad9929598e18938f327138443f36fda66070b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27fcc0bf022121d54007e888ab890bfd1a64d238ce4742216caadeb3081f40b1cb81edb44e17b67415d119a22bf5e69978018f64f8fbeed41fb27c1f80d513e9e9d2a4d036f4554e5def6584ad68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3c57e3ed8e1336ee5e34fd0715e209965e898d1a4deeff4fb1465eaa1a644a99800453d043677d0a563c6ff8585e4b14cd70ca3e40cbe429a1beb0833df8313f35491b52b6adfee685d18559f4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176917dc8def8d30ba96d9f269ce5be0970a3d9b98b1f31b7f5c2e1f82a23ce0c6625216ba6f09b0a856c1e0e167a6a6a3254e3a9f59bdeed7d05b13c15bcc3faf7cc57c768169a1e19512957f5b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcec9050c4977ec1225c600a906169399286bfacbeed06a3ce5c02d18538c1dfc13ff86d7a27daf3cc79a6395fbcadec9c8b994073e584e8ca1ac3dc5d16c89ff41e3e11fc4e2bbe84d19762c4612;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106b85318da3c897cc7cd1222b1beba2ced25494ff542f8fc6c6456ab756c6acd165117ec2d9b240844196c7afba8474a027d6a403b352c0e63bddc3476f500981ad7cdf7417d769a5bc6908d515f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f9b585a4cc66fb91dbe0a1e595803a5322917de9fb9781f0c041abdcfdc881bc3c628e1bf217ca3ad4d2795a55a7c6fed3bd007c8b26d8a2e6065f6465e780dcaa3a5b118ec5959f7249af3c20a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b27ff1320203767a89c0a8a622b3cd4ea15eccd22ce777d4bdd394c598100a65c78b07f6a0001d4c39898140fdd0d4a4be99f760f8a9255b7acb43b9c84e18c552338b5326cfe38a84c0fe8c70b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1a335efed1473e72071fe310b27e68b8229876933fcfb7e91f75704fea1274759c37d3c3bbf889786e1ab746f1dad8730f3e011d88875d10049cfcdb23fffdf0cfcbab5ee17cbb9a6cd8f477be8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce67498c39f199ba824b423db1385a0cc9e3e33520d27f934de3a8e17aba6e138ec63f3b1656fd520946ce27919343fe7955534fe4b722be2a48b8b134774751f3f35980a082c12d19b0ee72b109;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf2c229ea0260de6bfe6dab0c4e9ef9d6d3328b34c2e6eb857ec7a618c7d6296c6381a018ec657f6a103114e17a45adda0e68074c7c9f8f32cc4c3f8f25b70decf646257297b1b41b30f8e8067cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86035a070b1598d7d9654dc00ca86c314c676544f75ce83e8b3aa4290a45d75f1444ebedd2cd8c824cd53fd4e12a86e5ed528b4f9108e42526a5aad25bfce30c6777d9c1d8c46b697154ac4b01f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189f3afebe2f769dbf81a3197601b53a226e08e06f699f7069c152b814bfaa0aac0e8bfbfb6bea1db30a216596c1b9fc2e257dee338f6355e7211d3a1aa9f73ab2873d387cb27d382b5036773fcd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7f64b254c9561c69b2400c0bc563d7d3ff9d0dec8571dbe81d065ba6f99d16988556e9cadeae4f4b6d9a2e90bdb6621f3c10cc79232d5012a1dcf4736defdafebeaa5f19b83d14e3b7bc6740dac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e95b55e32feeb395c1dbbe015cbf6ef73cdfac6dce01dbe44d9fe00fdbdc95933e57a76010389a996eaeceeef2fa5224eda1dcc2eda704ea7713c5cbcde97532ea1df1b6f914c4eae49e2336879;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107d063f7d84ac26064e8f16db7a73dcdefe7cef3be56fc991febf74ac11f3516bc6d63e4f1ef44bf90dd9ff72e4b45af49a2082229553661b83331741bb751062f21e79a91e70bf21d5c69cf11a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd9a4098d473eebb7041803d710221829db1267b3e680008a8eee374c8d5db9c046a5cb92ff731e53ebf848837c7e943d564072f8d35c7970dac9fa543e818ece51a3e74b7e74d302ef7d26e72ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf650811d5ffc84f417889966d2ce0071f43a7c96cb713c7cb052ba64fec6773cfe8852b53ba7f0321cf3d4d9f1bb8cc59692a014c5c8a41ee8ba0f02660c954943d1a829f6d9c910197893ed50fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1836f0c6d177e72edcab7b619fdf4ee4fcab819bcde505e43c4e824ab8c7fa4217d06f178a9e46e325da0a52690ca76f24b86b6e02418516fb515d28a9886ad1c726e68c2e52d51f9cf8e42d4e906;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b53b301f0ddf9d165849de12a97f324646ed7132a7dfad9ce92673c61ceaa6a2190f5701dd68c60c8182b1dbba7b3b4491ca1e0c1efeb182b61a4a948e462329aa9842a6bac2b3d3cad8cc59020;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109d78fe76ff9fb8d0dc9e6831615345309e7031afb201b9db8c2875eb0f48cbacb814e914d99febed7eb80825ac66f1fb2009c3f2d579dd7de9f4cbae6e7caa491b7ecdeeee896585f40050afa4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140bac5d3695771f23f09695465ed8ca5c29e6431c67d762543d0c3c4a1caebbd689f70f59e79691ecd62c3ad85240fd4b74de070663f516060a061ea70640a0973749f65034258778b3a8f90a00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1926794bc414069736c745e26f379cb8f8634879b30539193ed216648cd85ab8b703ea8a3cb97b56903bba9727c8e20271025b2012cf9a0ed752e654fd8b997b639ab291a742420421ce9a2e7a115;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb75e6006722c00b0f7da7e09fe9d1d6b55030461de6b5c8b3833e5fe07c74584704c887957ca7f5bc1eac37414f8fc9c7cf35e2787232e36fbded6945d9ba8997929cc55b5813c57f9884feebd9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd4f821f57a4237474f0cf28a44298250f10eba60ab148a445722b6f2e47d4bb5a362d2aad3618686b6c7138702d246b2813ea09b91310841507638d4e3d886301bca3ef467d6e68228a2110ba93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda0a3f78d5091b2f3513f8a23da645bfc09ffa37cf7994c9abd2488c0b29d96d09f5d2f60f4bd086032612eab32a96b1d5e7c4273ea86e6285d34c9bd8085411d0286c54edbaf88fa3e5071b221d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h599f47100e1ac3cafd198106b4b96a2a4117d91cf72db724f4e72de4faf66be169f4a222268b1d77716fe131412df8ffa7ecacdea61f816ca8c0bda16c965fee7705d671080a5fdd749b4f3f799b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d87456352ba62e8c7b71aa829a3b9b2a21079390d816ab129db34e05046e85d33304a44e6115ded92ead4f543ea6a5950385718420ad319c63b620f31413a65e9985e2339bf8d7d771c8e7e05f6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf99ad4437946239162d24b367f6bf4213f9835a092fcfee4c6c16dc382909c671680da68f008016e227a520c8c2272952353fe156b0bbf49ec748bfb2dc1811a9d25074c6f312fa316f57355f98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd5ae11bede517ede6ef8bcdd697e58acc16d8340e5448522e8372df22982cd0e7a90a81a304842b1318a4ad150ae5a9575061769b6ad44cc6d51171f987c5ad654e1f46575c0673b18813d51f0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77fe045fa6667f88f41602d52a7bcb694d1ad8bb22b5def795289bc5e1c2890bd3d83ccf356d652b89d64e62d91d303c627e0e34dfa358d17dfc0c5e4d6f0544d29d75cb8947d6ab4266794ceea1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86e95e86fd45a5ca79b839ebb85b39d4d6c32092e8fbdfaa09400976f5261900f17c01e3ac390ada94f77468c780f7d96d58ebe5ab39dcd288a25b45227dbe56386417defcb0be7ecab96c5ef247;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cc345c0e5c1e1a4cde20f320ad8728367809e6df658b61660ea5f021a3b0194afbff62296cf617e3f4bb75f38be68d2a9daad18b4f43697147e1d16455be9d3317b6827de4ca486e007057a6ccf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c7a8e4f3ccba2a97495f86d5b1c86c5c3336fb3c0de27951c8b2b7061d6d303786e7fd23a0a48f7ab54eac008d9e32fc66b466f93d29bc7b3f394ac2cd9c9df729f336a3877a33e7f86c3dfbb10;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d9343a47d4d91eacc028d60381ca424fd258910a3912a33dac11eef27c3a5cc78bf86f0fbd88a31e4e5fb84f3e9a772048196a8c5a4f71f03a629e2688e57cdcb0e693cb3628324e2e56429efc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe686a0c15f54a59284ddfe285109d570ed9ce4861adf7ea42c121c31a83501f0aa8b832ca3a68fb5b6473b0d717a55016a60a433bf56950934ff1b6b7d8374361aa27a97211a4507c1144584800;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc91f8ab0a16f6e1e813b4dd4f50c4eb4ee6704d61fcf0c216a8594fea085ba190ec560ffd951bbdbcd1351176087189f585c3b2a9e8415cb378a3c5afc75d1d439266361a018980e4d66129b18cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha19f4b471c884bb0da71e5ee00ce7d01c96323cb2281123c3a932434ed74bd729e676733955e100f6efd02ef0b9554d676afa11f499e2a5764a68c6aac97b7bd31e26c83c4dc4afdf00872b7678b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbed32151b23e9a89188fe2d65e7b3a3de45b842de7a4bf7b71ae0faad84909f448f63e978c034cc5c361971503353e89d5f478698a99d3360b08f53103faf5abd5498d3cbf2fafbb9aa8e5fe5f98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e38f0f11b116ebc8473ed03a56a3ef65a4261a4ce975702e9cbee7858d2e46c84daf3a9f24bf4142c56436b40cb982bf62a87af94f18e789ae4bd5c2de53cfd4e7d77cbc06a31fdab56d497161dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfde3e509ba47c8bad24a799d32ec5f896a403c4d69dd3fe330ae44590b24dcf9212566d009035de14ae06fd8523c09b011fef0b73959f800384904be37d10745705aa20bbc77d2aede608146dfe5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5b9c7573d14a87777f25119520e759a38ffa61e28a87baa97f2b8af1c81904d4a464d27218546956e7ad9030d2ee177c270ae9d49ebe3c33f01e0a51753b8bb9a8ab1b98c38f332640e42b4a39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193cc7d7c348f1b3b00a26afcc2353d826f93bbb8ac11772ac83cbd6d91fb579858184cbebbaf963f5cb6409da4dd18a37f00f2be85aabae0642eb869cf15554f0e9dae9698d42cf6518404fae283;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e395991df6c815a0c82add525e950c1dc08bb4cb558cee1ae5f67ea0466b9584d8f37c71e28be66104d03105263753a74326111afdcddf877b1d826b42c91f27f98afdb035ebe5c8771b2f68a7d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15500714af6bdba426155a1ee5b74a7f1e08599a54887f90dd48248bb93ab21bdb495a56d568f29436ad5034459c4a4df77205e114cc858615df19906e4781245106e19fc68c6048619c32a0fa111;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6cf5b3c2b8d88483acd4a1b1b0898ef94fa6be73ab3b8305a101fe76c20ef1c61cc06a4dd9a13aa5f167066ab9fd624320f22404e48e45c9449e728db9f5bd0e2d00113e9374a331b511a9cba55c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ba157f4cfd5557dc0a44ba7342aed2e72a35bd8323794d4b025175ed4a25e27c38a0d3a93d9bcf609e17aaf58a1d78e33c756751173b6ab52268af888fbc9ac51c43fc12b1292ec4229aea2789c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6cef471b641712e38632834541676c953a323021ea07de8a63d24676c37a5dc9fc08bf0a528d7cc29d2fe6f76ca76dc1ad295b58b27a64d92bf33613ac1b33775f7a92ad7844ac36ea1ba1c6ca4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ef307030dbe86f9b55c7a2ece5ffdaa91c024e1bdc9db9f7f78c94f622f0f0fddc0ad5ece8e7936ad70963c2aa43c532160264987c23a471a46aea23f15d6eb2b0e87296291d3d8cf93976febd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3797eae433a796af3251c510a2853b809ad36ee18842fe07d5d8b63dc499c3e40ab87b7766058ad7260c2b1d0eb5decfb55c3c2bcc5df1484b4cff79cde60fd488d4624a97b27a60128688e9e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1160019563c7af2641fd094f6b1568ca7e367a4fa6ea9027b69866d6900d30b1c845d764c15bcdcf188bd9e32e74187fa65f97940ed6775d6d76ca27d6b4b8e616b6927e97098962f11f4089a7047;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13027f2b3a98a10c576317ed9620555fb4446f14bb0dd1b43226f708c9ccb7972d9a3132474c207a5b31987f52df436943114d6c73668b61166383693f7b35dbfdfe447118a7bbed1cd365a5d2310;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f6b81345908f8f098495350dbd143748e60723574d3b10eccaa5c5ad7004e4cf7861b7600f0d9b0abd0e8f278beda5a1cb56a305d7f00d1cba12062718529bab268b21aa6baf5cbefd4d0e6518c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc96affcaa0293a5a45760723a6d78560d6b5823393e842e4cb4d07e41401b387aaf4e59151ce6166119b44c8d408392c86e772801539afc3f70c17f4cc9fd1901561f376e0545405674d207e53e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f12035425946a97cfd0e39dd8e84bb13a514fa6d273bcb209797f71fac0bc295e2b4a58738f834423177d9662c9c4c81419352613c621ffe18cdc05f4ef9a14bcf25220a5fa4cd4a1cc2368bbc48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf0a91218e6b30dd58a7313e71fcb009ced646590eee8585a61643470a14acf05b5cc4355821f60d792326afe856bfc7ccd7fb4ef0ea5d8226186253bf5fd2b2d9a84ce4491d32c223c577f4c437;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ea1caa78e63a22614210558a0375ce1d6f26ee876540ae5bd3d56e1a3b41831524239b4dc5ea2d71ee86a57468877c66c73f77fe82ec3395151fe37f0ac35a689c72ee8c60f00e5f30f466fe2b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32c2b4cce2278abc9fd2791246a0823b2e9cbc8c73d5f54be5ce7e6e2e74c292ab7679e624fd4212981d19805aab3a4b4885765deb94060b0b1d2ec8d9a2a5be98fee458fa09af692d2626a51919;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c87ec77015286238c17761065bbfd29f66688cf54868ed11b6ec4475494b303b5963da174b6f4cbb0c601bd6ce847ff720c7b205020caefe3ac5f980d29d6611c7d755fee55d5e7da4b41a034f0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12358c301d26a505ff6fe29a4b892bd9f0bb965f370e53ddd967c01e058351ca523c2bf658b5a1d32db1fb2548e5d0535a7fc20677e5c1c5de4c8a0a8cea493df7739077604e1af784b56a0d951d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1166de8318e7bc0dc21bbd70d966fc06d4eab99a587225eb26b238892eaee94ad334b7c02a0790ce0a058e28ed058b0b4ea9bb9280bb26c6db41d1e76b87e439ff18e0b892b83ff8f476e8c1f5ff1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d8cc3a39ec1ddfec60ccfebcb3dd534730acb9b693863e0d7b20b7422e25c517219cfad565deb5d40c146ddcf9c85ee9098fe2fac07f0db6cae8eb416e63b3ef09742a1e32b8b5f509beb61e607;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c435f4ad7cc9f6665874442ca48a060ecef761b1928c9e54f1c8a0f6151999cc01372092704ec6c733a0f3db66ec0d332eeae18f0daad94b52391c9a6e9d2de662395cd41385536221533c70d0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196b65753f396dad3fa5da0da7bc2a9ba4c7a3816b6d69fb28a4d3928e1b2946e5a801545054eab2605325928368a9e445394180a60af47d549c227d51382d138c7eaace07343db9eb3678e6659f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5bf0fcc63d9a5c617deb3794b2a8c8a234bacebb1dba44ce1f0d9045ed88e5ae6a7d8875af3cfa4ffd5865bed1cfe85f0b067511a8151cfeffc0b33c8faaf7614067fe997812443d73dd368ca5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4be7b2d1a220483a22deaebd0d1b2292bb849a71de54b212bea71c99b62cd90eeae700ba0a0e3cb4698e3aa0509001decec20c2b83ebfc269fa43deec05fd0921618d72740f14c0dcc500578151;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd58ab41e0f5815ccaf5e4e53d3d7a6425be1a844d75782ceee123bcbc911bfd9700bef3b54ed7847373c2105beccd313b15024687577b8d4360e1b99a3d4311e8d0752358f683030d00163b94533;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f6ad095d9854710f037cb745e3cca647d8d4e78609d0430c72405f90512352211932af0c5ac9e68d120e988093db9fb2cc980440413319112fe121bab3a0fc21ac8aadf9489bd33477437c7904;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h493aa9b61c8536008f209e9bdb00f864d98cdbf327dc69b5da634e026120758c1fec4cdee4739740d4eed37c05bd5ba129979f9dc3b11c9f576171817f5aff57484084d11c861757417352b43e89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a835e2258f56fe1f049fdf0a1be9395c68754aab9d33d741a71744b01a6af0d0191fe198255001582fa5c7ac05b511960af0770c093720c1385d0ebe60f4d5dcdf403e6b62b0c990397bf008b1ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1665015c6fac55193e8632c4f5692956a0dc6e52ab713b97824ffc2a9b364a5990074c0399396f047f3600e36bbff5a5da775c04c9e9b5757e53223ad43bf6185c891a5b9dd5f6d4e0e172d1599e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f556f25841da0d1e0707bdc08a977ed90daaa1e91267fe085a0e50d5c97a747d4e27369ea61d41e1d6de3b741926cd1e3fee03f7cb991c14325b270aba5c06e34b735f2ddbe0e0bc40d6bfdc4f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cb345604418ab23bbd973101c6b71261f79c8e80a7d9b73bdbe8fbf24f719af2a8af8bc81800e343bd72bc3c43eb3bc5b89933d327e8ed5377ca5fd95e1eebd145d575e0ced41c4b86c4a53a24f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc890e7e08cb6dc10b00c50a65051cd6a084b46dfa485c62db5ef2137964e808d1d7fd5d7870306d70f6e8171de4c7db91d1220db0f1a49d50f072390eb16adc2b28873349b1ad811daf5a6f767fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b4cafef11cd12e99b20ab96e0c6ae86f98dacaeca8a90ed3ca6857c793fdde066fc362dbf9924e5d13567f045dcb091d779a9d3c142ab018abd4ab19c2998c6c7a45483ef982cea62e76de092a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec80a4a248637cde18b3be1ec1d857440c8e70bbdaffb9dd5d88b21f0bd8d33cbd5bd8a85489b6eba1d6ecdea8c02c1e1198be3f80b0dbc36789e4d3096dc0a87432983097a125ecb20c7ae0a4cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f667d4e3de7337966a2517b60a923224ff98f49d9987e11924e5f52c91097b6eb0d9f515c7cf264f6d26ea0d1ed2d1c63b86a61274a1656c7e68e8b6c70181eba10d299b61887a6ea970daabe94d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ac436b969d865b97d3f7e29ae964866122363390abc3b899b4076f8867610a6881afc7266c1968047c709eb9d10412eca23e1eee8e5cdcee4d6a53cf7f23c8907fb9ddb177c6783def350608b03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127df4ccd1865e78516774c1bd6047fe3ea140c707a6dfc249dea533797cbe7a32f336de199c2b28891634723a9ab15dd2e83b8fe3e54f5b3eb747734cebcfa4e74a26c667dfee7914324c7fa1c91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h686abbe8876e59fb9d02888e66107a9a026cdce5cda76fec434a954b12b645bca1ddd21628fb67c4e6188ffe3017e6ecf0d88a363f063c046c59e44a1acaa3f2f33b445619b61711861e31de7627;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191f3fb918db190fc405f57e48e930ff6fe944a0f4cc193487d987bc24c69a52d81b754dfc7a8cce382d5ad79420d13bcfa00a305a21ac59a5439e79e97c76c8b95ea4a656ec29caabb0aa1a36b80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161e6a05e758f8edea7423e239a541aded03328c82fcf59b39af90079a647070a77fc56e4e75830114bbd95749c7928c7db9c6563836a047629a391fdf98153c20b1a88075f488a11eeb04b35f731;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a07fcc88565e1f902909fe5322a963eb335522b0ae7c0d14a559123bb869adbb00ae5d61636b8eb5422927c8c40dea00e96cb0f3bdb63597b1bd643bf667d951c5f03f0cfc1fcc9b86b92d2032;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149ee500754db9e518bdbbd314613db8993d916f6701f4906d93686a60da34d25e1cae5106f7071bf95b2bf17395813af4b28afb5dece6a4b35a8e04fc99965ffcbe2a3da987861747ca4c0cb871f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10605697820c90eec8a0d65f173421f6ab43b99df0605f17d72045091dba10fbb76e9295a34dcfb6897062290251b5013a64fb592562eaf53094d5d72dc066de1714008abc4ee35c227ff0f0713a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107117e8a5c7d64de0ff638915d30f293dbd94a6a292f5e41eea7474ce8704ab635dffae1c2868f66124ae5e57ef72de79045e86b88e7b8f92260b2ec7340da8eb8e37fdd92626d50c2b4485fb914;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125c70956e9a41dfdf27ef14991ff111ad16221527401a5799d000cf67a082a405c77e0bcd5bbcb8db55d23bd17bf0ba1be2c201581a31948912c7ef73b85b90840d4e695dffeffa82da6a19a6f65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bda5076c77885c533376b35f20c00457be1546eace43d72a753d0c08893618a773df236abe907002709f24f6659c9a75e5d55968cac9ed66b536d472813d4035248eef6bf6a876d7c47cccf3bc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e22d536a55be5b535c3d4ba196707d442bdd8046e8fdd96733cd738d62e96db8977443a3c0ca61d79f187d2caa26f1257ccdfc58d7d5b54b368478886a3fcad96768eb8c9216b6eac8f84f54219;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f620913e038c8c9e7a857d1e9196b853044d03d4d71c0c23fdad9c54c5a14e9d0be7d3e879d5eecd2eb489bdf4b4918986de16987d9ae76fef292a99dca85ebaf1f9e2642580e6352362497312;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfccf0b2d0dfa1ed9a255bd52c658e7c269eeb00622a953a0e818afe45670ad915b7c95e1857ac859ccaac11f81c5a13367b828f7062ecbad49ff2a2badd91723565b3e99a4788501eb422281e25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dcb6a9c2d991f6d3e7725111a2ef858143d918921483ae0da781896a4c19c2d881f86526cde0fa99750684a776e895de41ee0edcb5fab449ab42ccd26dd76f180b768fa803f271d03c8f7bf4fc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1130d9166f8129350c8f9cccd4235f7a914528f75303024be6578935af23d3a49b231aa701ccabaa8a6b6066816dd11a90f3f6058689ceac0cd7bf5d9fc874212fa1b45791d776cf0b0f08226e87a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11196c94475350526c5e7403fa892ad4158eeb53effb1381161702db0ea34800e59e832e90a1406cb343c8772c00b0293b8ecc8e8ba9189bfc9a42826e21143c99eea79b6d73e4320d1c073961946;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19939b1c193b88368062cf62a2b04fccc71da36b9125a940cf877bef8cd300bae67e89bc42bc257e3b0b3d5b6e3748f4416bda3d6fa813193e1f4851d4b3ee4c7e5a6cc084f74e948b6abb090e8e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f374ade6eae34d2b38a01ad66a40a415c8b1a331a681093725d5a6a9149a0709034b33e87695642d09ee8da61c31a5826bc5bd3e7c4a9f99edcba6203aa377a72dce6d642be8b4749decbdaa8648;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d9d764f17908bdce08c8edda187e856d2749b84649aa4b4c9d64db0488ab68bb0072baae6a3f6170177c7ef01afa9e62a7d93be9b9ca56feba8d9d3d100416ab8a1c460b3ef1305d5da39e56b77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h229c924d52537f82c713dea2d40a45b394bdc5f89deea663a3524cd27eeb12d2be6f334b31a40ec0d47e4cf4eee95aa9d3da8f0e42cdd900977fda57d6cb7d04dbd5047128c99b042e07d5c68817;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9189bfea4b9e7d202241d60af5cae7cde2a90bc8eeabc0b997eec38eb71989e962227992a41491f852200eece5b51bfb9705c433905ca506007cf47469105f97ab91413056414588419a5993ffc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0a83186d6512aecaa6219808a826b421c8d55829afcc76a40ae2383b45abe820eb16e4928402cdc3c405948198c5ea9182413b3f1dafdbbe8577b3d518cba78a7fd9b44065c0509f62c72ece852;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193e6c4f7796c30de54d3d875ea27dfb2bb3ad0ea668504096a16dfd683cd689393ca5041b59513633144ecc50239ce0e3ee968b2593a57a70d29b64e7a6445d1a55448883d13ef9042d9a8fe29e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19bae57403a9152128340562aa68204b63058d51436b6e7235fc588a72025738c63087eaab7e2295fb7b8181b66697fb69d16c909dbe9b40958a06c5f63d0855480a514023b0ec8b8586f5ee0dcfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8fa2c93c6131823b59fb9e4e40f3a8e17f9a2e2198374588278be7c606813045c04bc922702500627850bccb2081ff7d85e5c4b6f3dbccc230ffc60f95c858fb426b4b3ecd2afafab9a22715f9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9dc6ddc6f6191c827937685493088cd3114bafb3ece5401a4ef443bf10e86bc599b14458ffbf664b4271de6797fb96b4396d522a109fb4a957e69a5dee19553f19f41b64bb72e1355cd3930cef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17900b8f1e6b49f574be25a373fb6f451d2877ef0b0aa694be6d4a10169c4ed1c4dccedf412b74843aef51cbb3e1046afe57711d5b9760da4f623cabf2be5fae8bd1089f6ded13a2bba917ddd69af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41e169f0fe8a4345899438639c974306cb732502a4a04f40c15bd2931c6cc035d4a92b6a56b296abfad8061f1daee15f1df0386d94ce3f9e58e9e508eebbe541fe17c9a15a889570671127352f33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc86ccdf3b53ce985ef2373a5985139f4675948b48ac6d4ac268aa0eff7e67d737608f4ece845bb542a2cad5711671ac56b861c0d6ede27a388ed6031d538d7de9a07488b6fe899c5ed711f134c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139cfb4ce085960dbe5a497112c845e8d259e86d33307655549b4c118437494456f745ce8648856ed0efcff458507b22ccd4db53213e59d85682949c1328969e106abc2a54b6eccb72dda994c1cab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e514c0d85d7fd6ec29c946db7495574fb2203e75a23e9f6452483df6c1b3df864839a75a3f7925965611d99cfd068e4cc62a329c981c831d7518f19cb3a7a5d5a73d042c5f7801c573e346f6fe1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1901944d1b3e04539b9329fc3a4e63d5712c75bcd53538dd034a0633016c1854cc87b03949a22e9c08a4963b9dc994ce7c0a483b736a103457e9a825764978f84f89ad88a1d8e22e4486f14da04ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a1b03688cc5ac27ceddebcb00df8363caf62cfee206b61b39dd15afbe3d190d2eb7e052c55cb5dbf484a45c4c2b6a5f366cd1b9a5124c659f2de11548650ab904ccfb90c287cfdc331a538e76fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a9ab1199a319195c6a837120fb78c791cf722eb944622568e5af06a0e829e070e8b668c17ecdae640af53ce05460e5da6571e2ba3e8ab6e4fbef6829a18e700c765712b63fbfa45ad1e16ccbe26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h634c2d845ca99aa10abde3eefca2c042844603a69e5ac69b23881a90cf44fd201ff3a1391486e507fd69bf35ee3e76089500b56b4906fe6bf9d4a1c7887865a25c2adc257969ccf35be6cc9359aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b078aa605231b0b5b3526730a9e23302bc62d501d296ff88e3b5032048ed655555464fbc530449390a486f06b48c2646e0eb3540e1543f8b52cd2809f7eb45c9119ba85a330f260e1f084caae44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f85ac810eec9099dd6d4f399070d6bd3c30dbb8b8689d958cbc465ac4c44e123c6123e89adc93bf3043cb7d5db14880d281d6c1067067d5243bd5d5742ede387ca27139b7ff9a94391c5053f168e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6324a04dcf013f115e02d9406f481b6736eee2ec27d725a2a3243d748af41365a33aca1c23f7c190dfd4f7b943af0dee80e3359b23b325b9cb04e90643923bc29c0081830021dad5af66efddcee6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h51102d44827fbeb73bac4df994b70c7f4b1f978d5fb388841b79f990bc8283dcb73bbb7dd974db6ba03ecbd7bd0c0ec35ea318466432134f506640397b4e8748699db18a15b67c7c533460b8037f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h646ee7677d015442ad1433e90c3c92e67a04cb83d376f79f0cf07820581ee25203f35200d8e000321176ece48d8c6017b55703effdc46806534ba4a7854ea3be27e5b675bf0ebb5cf773d3192fb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfffc69b6934e7e2e652d55e93a5c05359c4ce88660b2c674897210d1ebdcd75d0504d161483896215f30a071fdf813655d19e2b581bb62897ec69388dcaea4bbac6e7b57e6f0cb36257adf08ce72;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6e5d61b216c4e0b10f9d269d1a0bd8745abb71095d99884b9d88413245c350370c5a087a0f6c98c792a2e7fb86959dfea0ae632aff3aff7752f65ebe64d1b53b253834296c0546982e0c9ce5c22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1051267016adf7f404d7792849d928d3d5b9fefdabbf6da22f59a55f5aa4baf84c2e80173780462de1d917f26db60743fc6ca13fc4d1bbb65a3e807745b10580b8548c640af18e228ae772fb4b892;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h948c4fa3405cc9c8fbc50ca1d3c810ef82ea8866cac6ba3fc555f1ada895a9969babb2eaea6eff7635186259a7e6be40acbfe48d3aa51ed17a061269fb6c84e6d5ca98442feca548a3ecbb9bce55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42662f9217789ec4baf4d5b3cd55bc9e29725a8535f8eb17249cb021bc423152e7a84c227df5192c3443c803bae48c1bb22e11a1ff1a9cd0fdb7b0eec1bbf10247a5dc837c8fc61307fd4fc7ea2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bbb42e34f5aa40153fdaea49ffeadc103d15a825d581dce97a2b6a0d3a3bcc1c6e79248815d070163002214cdfef5c369be70a5fa6cbab17cb7db53f9d0a332f8fa19e1cfda176559ae86a8a224;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15feb7b2fe588b0b52fdf068dd13dba505b7c255fd9d481d44000a961ae52bace651196262f04fa1f4ba9c29a031b179c9f73c40fccd62a8b75d38faeaac1ea242d83fd6766149ca7a34f37b858f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8000e7152fef7a80d5b987fe798ad49fa07d60ef5eec4c7c8c2d4115dcfa9fd9bf72e528cf92966a195b8f635df66752641ffa289e91c7479c4fb00e975f7087ac3bc75dc86195a9138013bf11e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f66348a9dd8fb2acc0c2e839d2b115b4db0428750450689fc4da8fda514b4d64eba850a9c99e21c7b5751775b9f6d8f42efe3e14b5204e8744c9f276110caf1b36dd37f58831d48464b64610b6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ba2c4f52224eee14af6f35351790aa7cfe7911a854dae7ef92fd5b943ff64acae771d9fee5fb322f930f81005b03710fd015572be9e6d67a5b312be6fb0bdb35cfe5a0676c9c7997b882f5de77d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1facb47b0660624370504535fd10c0544015711717a891b3b63841182d706e79dfcac35b0b026e334a5eb5e843319a08e6ab5cc7caf740592e3a5c84ed4aca747d36a5e9b5221ca8ccc69aee89d22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fab3aa799991b3050e780768de7e1f8a50fd67d713964535fc383e499f555755095458a26bd9fd8f48e69304efc7ca942a055715c0ffafc2a6902d97daed5d09f57a7a2c2c0e8dcb591de260d6bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18483c0c0991ce3c1552d516e6fc9bd5fad2b7f1bf3fc295941fb031021f867e9d9b50390cfba017cf61e679ab1801f42e458a9dd546ce22f385c8112840bb382c765c5bd3da332980a437eb68b9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a61c5158bdf94b393f6bce73bfaa12670ec1d37cbbc768516c3289af38573ee24f4dcf5d04711dabbd6e2e7af3fc717cb3ba99411af9c1a9cc2e8fe79c6622483688ec323eabc362afc9edc068a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180f00827a43414ecbe033a94ba56e818985b40db2d28c3b0b372e9d66153856a2013579d9a3c4e3330f36af7b9ec999d9cfab61fffa9e2fe50e5c79f134ca70e38673d47aee7e63e003bd97649d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf090ac927790550054c907f5e9aa982540c95f93f8aba507373b5d09a88ec24a73e86872d661c317e34306fecdfa27b8807b99c79a3c5ca2a29c50d5db92748124ac3333fb780314eb4a0d6a9e2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f03543676f6f8dbfc5da40fbfa9a41dab07417f6c5b30fb8ddb3241872ac65d1625d2bc6c549fb60da4efeb4128073e287651ae5c521cd04c84d5d82a6705b7d8e22b88adc18f49c6eebc1f9170;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7cfb03d49aeff50e371c185e26fe6821621ade3ace9c1f000a4e09dc15fd2b078a30fa8fc8520318be4209ff84f27ff28836ea5d43dc0348e107bbc7f3a6a3735bad2a2034558ce0d0c7a2cface;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a84cd43f34d7512960d61b787426e99268c45315a73407a7768beb48497eacded8e1f9d0da5df360f0e1b81a594e745e350b4a3cbc77182e3e6163a33dd937602822624d68800708071159b3cb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb73bcd5ba8e0de3711b171db6c5b968a9a0cbbc632bdd0ba53bc17ce64af15aaffbf13b7353fbec15dfd759a2f5a3f04f8c91738a7876ee9843aa809d68fac0dd4ee0ee27f12648c00f2ee4d64d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdec6fee926ea80f74b109636e90c8053fc7529b2e9cd421e6c23c356269b939b885837ef2cf4f5e018e31f8fe4222b91a9ffd812d1714fff9a60aeb19275e88093d2d468f93434eb65a7fda1be7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145724aaa1295bef616c31b89044f0a2d2616f840f43b6d518197c154406584364c26f65de0e5901234bcd04201f6b3496446e330c14d55d17c86cf3f950c97a04d8ba629ce889ff8eb0a297ed6e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdd46e4ca28ea94b721f2872aafb240129a0b07bf5a70d9106b89197613ff34d46b5c4dc79d34140046be14d800015980b2ec507d95d3a7820190f7cfba7a4687f6b263577a98e78ff37c46ef0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a2fb7eb0e7c70c31cf46494a75eb384935c7f45267c4bca53c918d7a8120876ed271e4fc415ebd806a4ecede7aad805139bfbaf1ba41038c8a2d71ec25300e8f9ea637d6e5bc1cc1d90965df3a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104096291a7ab2820d23e33f1f4c7a773d14e4ccccd748b9e2a5f33c5a73e9082a7aee5c15a860c6dd8366a269c41e40de8f9dc7440b5cb188c4c7462c064b33877b98e0fd7ba98fab7aa2451a7dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd940c7a395811372548796ab0ae000cbdf0130b4fb50820287d51f9d8d58812572ac8931729622e2a457f2b56773dc1d3ed9d8370faf70ec866817fe1aea8ab22fd1ad688d2e0b8614ae28bdf225;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df7faadb14ff1c4448c8946be96a8565d23d857fbf1eb38cc4bddc6217878a9703076f096b6c500d1aa341c0d78fb7b1604a04f7f05b5713def59ce7a39a64c2bd103f4c7eabe8f9fa30129bccff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14141c5f8ed97de284f5872a3ce0dc400e5f98e27c46ea58e22e8e78d54d76ed1a31837ecde8c61d43a319dfd0cbad750ce08b3c26b41376a571916b18fcfd7eb1f49ad2b69f049d2c0d2998f0dae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h502a59a9993a5707a63807df3044809cd2f43940237ac274778761c38e3b8db6de7a8ac96e6638d74075da7feaa361ef58df894c314a66d8c8e504ab326b7085e1931ec2ec200128654023307cb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heda7632c5313d12dce63c0007b98db035a0ac73762c4eaf5a48be92d73582d32d4389b68bafc11e3af6ab447c0dad8b5fdb022997b1e726eb7059afe5e03da972db90735459415aa5febd8be223d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158d26e9948e7c3ea60f7795b432cdc2b2fac413fdeebf8a8ecee99db7e46ba5a304c8d2136c8e1a5b5629645269849191ba2a494849508c2afc5a3523651285d8e4d00702346431af85e7ab20e15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h253d8bb5183b3302fc9f4db5fdc55baac4ec1ca60bd01278454de215491d18854bfa18f8653d2c9f08d2185f942545642e222992fb27463aff3bebe5749ce1077d17d390bff7fe8b7c72b8f58c89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hecf749ba33c93f4996f9f80b933cf1d67136acaaf7116c8e745d093ff328ba869375e7260762936ad992d2f1e2d8e675d789ff11a116bae342f1d1b71a483b712af8d3f129d1e1a61fd8fe7692bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16195077ba79950c920e8f8262f5ee13d5a8efc26510e406595cf6ac02e0a121afc33c592b23cb125080516a98bfb1d7b74360c597434e1fa6d3f75c05c216f87854b8ae2f74a07e1e9b32fefffa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38d9921d8cd043fe6e46ddedcfc8a569c3e59f1abf5ca4d78d25a2ab800be50b2231f5dca12ad2ec41a7e439f5a274005c0ee54cf96427c8d48cafd1286aafe32af45d2beb25cc42c950cf531af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h666fe5bb03c1f90393e2398be1a5520a6ca7e74edb41d984c99459267933cffd52c4d10cfcd9f84bd19302d5b1e173f4ffa95c55bd63215ac8b778f8b27ad03458d7ec9f99774ef4e00e58d081d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb8100a1f71b6f69456cee855f5e60066a118eb7cde6f14ff254463c7c3c22efc0994d93862be39f65bf41bb9fcd35b27ebdb7e225c0f770a05fad0e735305b7c0a92acbb7444d95b45ed51e2ad0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc83659f7f0e1d5d95085a294ed06ed464d031fdd20ee6823ec5199613e21938233d19a7e52fe32db23f91f8f7b6abeb6872c4c37cf7f649fda1f61e7a1cdc0302cd9fd9cc3fe034b784e50e39a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1833a98b098fe9a8fdf929c841fbfb448a8991bb434d790781e8f9ce1a9c0551ef0d510342867db1048cc808505c6dd336ed3da9ec1acdc9ea302e991b5126a44bd1e3640e58efb406efb9f8bf74e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19af323094614f47d1155bdcc0c478041326659e907c701b3c2752e456e667c702abf9599f942dc52a01e685dc81b7133e806d581b6ab12006f041fd594217e45574cf9abe11ab7f76bfbb938ac80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd8d3a87c53e6927a353448637e915a3deee665f6732ea0f0b1df8bd196e20e7f1407b11b419eeffa1df9f191696fd6ed3ed16fbbf71b7b497398ac454344fb0971ea553caba979930be74056681;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd0f4b069f8f2108a133070b91688de26defd95f68278e2b103659c6ec6092ea8e9dd734643417ffa4771dc666e2d8cbddb610f6d29dd45e1336d1426210ca68655fd528e61710bfe1162c19a423;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fb8dc6d1e70ca090e7d4cb070227bf76e29e0cf55d221f545d7efdb7aa642d35d4c4be59bbd1f42018d84106694bff0b4069339dab7152427b38b6e6268e69ba76454928a416fc3f5fe8acf0fe1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1006db2b9e0a42b078fe9c41b53745bcee6cfa7f020693fa89cc5111e539059e2e097f007f2cfbc7f82e8a2229e9a4e286510e36d08305868af0cea8de4e2a2a8d4264f40749be586ec0c00d57426;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a822803371b1264551733ccaf503cbd208c7b768003bad25283a848c1d8763f24a9d624750a3095239eb451f2f41af3f30213561219a2f43f71683d8f712423ecf88fcdc05288d5b88c9ceb61fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1379724d68995bdbb027aade72ca61c8b74f282a78c858ef451f367e97f8c4d2cb51445bcd9503585dc7005d28547b7042326083d6511c94a550502620e62c07050ff6d992960ce6e07a221f85c25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4e5ac32a61df95edd4894cffa5be33c14ad84905fdff8a29862f17c74c0cac5ad17013f11f42afe3f896955e52ddaedad2ce47627c3eb297deab42bbff4cf4697d144f805270026d2d102fe0e9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef51eb5a10e2c577ddfffc0cd4cf876d28910572af6074141da2a7c3b57fe951439ead58882e092db67a54c7f5487c86816cf12f0b506e7b523a621fe6d0dee9cc6b61b693c20e119955a6838b97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aef97046220dd5e4ddce5363ba26c9e6e9a85ac4b6fa6f0d9965f49148cbc81ae670988d5fe1ae8b78869fe07e92605e1ab916c3ed8890fecbc4d8932b00e39f6df9cdbfc90d9a62bdf79468f08e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57497555ec3caf07d81c2e5f3a5316ef78ff264d70260fb4d8d35af85ad161da781af61e6cd861ce1d380a1cd700290c98a7cd3a865ffe75fd5057e8df9d376a5c199c688e0c35f91e1a55c4d5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18df187f44ed2a2841503e2bb2cd3ab12136f1e1d3c7bd919dd772ee85107946d0bee0515708eb41152d5150a21067dbd7fe591ad6a03c66e8a01a59fcd5897898eb50fec74ed3b49a09076e1f7c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca8f589a164f10f0851a050bc9f6aebfd61c309cb5e2dd4fae3aada36a0330f3f29ddb76f5af1f591485e8d97649ff21cdcbfedeb63820d4cf68b0794949f2f246baaff30c6fd690edcd59eb99c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bef1ff55348068521597004cb0096185de4d32dafe5c929d31b0c8256fc01c97312f1997ddcf0272e04f49cce460da6635521248bde8cd37b8617a14e51c4c4726d1bc015fa30931c9f319395ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164f8d2af1bbbcefa75e73040b41f4bcf58741425263f668c9a47a2fa5f51d4ea7d655a6c84b46920c53cbb29766269d3af7f23626cee9a97be59f10d77ed34f8356acc1521366acc0a5b6b1d960c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e70a79a0c9103078a234e827dc7cc3be3079ed002b91cdba2f4644d50e019bc2fee39759cb44f4fda3ce90a5d5683b0cae5678ece800b7f0d5b1f1b09d0f6158037f7835f1aaeecb1958f8fbc25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcc7245cc595072cfc721adc1a65e2c5151fc27cf146e3269a01e30038dcd4c550e72ee7cd3227102d40f74266f3dccdb952b0205fa28557baad64e606d51c3111404cae396a9e9bd29999b5253f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122689af7fe570b80b75b424a13c86edbcd1206833bbe78423ca736e0c73a207d0520c95bfd7a335da120566cd5aab26fda44932892b317879e89c453c3a77b1afbc9b4c1a4a700b4c03c0fa3b565;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b3a2897ccaf1614ae1376ef9bfde75ee2eb797879b7011c024a011407e4fe5a17f0c9349875cf3963c7503e8f7220ffb347c04324bf174ecc64f0bb70e2810ce0fffa984c41d3dc64da7a63e527;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187fbc0c2159894ad6ab0a31a687d53edc852d15d8f54d99e276da681d5030c1dbda73423e17b429a9140b0d94b8611f8895241acc4b0c6f776a86d5b3d297ab6e9df490e403943509b2ed0b96825;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ee5992dcec4beadd7f2330390bdba7d420a7a9da5e0a1e05a14006825378fb5861303f658098fd02994ed3d62d94355230946cee478f33ad28fd24672838ca34ba0fb7ee047fdcd7c26b81d88fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a53996ce5f20dc707e61b8a063b1b2ee5e4aaa4343bcd71d4fd141aedbe5ff928f10897158ba48c06ac8a62f4f027657b27b2b9360249d90b6bd6a5621fc444ba2e0b4571ba9be1dcad3f22ab4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57c2837ead6dfde707c5768a86c0bb6ba8f19f1dd701c0e24b7a352881c665d4bca8699e3bec052d43d89dbfe14ae60d51eef0b1f8da56c8c966f7f48342a2ddb0d86a3d2e63037f7d88503efbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c73d9711bad7d9fab1cc2e3acdf283d056699407530a16adba6113927655c626b114c4013512e725e5f67da5b99ac82df1b2750f078f0aa22792fa6d1eb642dfd3a97a009a114bfdd7ec59fa0bc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hecc77d4677220a3b80b062a5c143f5c26016ef77568c80eec503a821fbc05593263d997c7148a403dadf8ec7ed5de97019707923a2ae695353b56a472b020d121ee5a4b2b278cd2b7b95136d17e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad93b9dfc7e2437360455275181fd29b592cd587eeb521306e81a88264e88d6ef01f42de88698718c720d156a900b979c247ce8fb03386f28cbc67c74dbf5aa2a50fd370d15b4633a66af5af1e0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e63ae9cc201cda952b869cb2a3406ee6a1c59f8e18ed53f811b3cc2038ffb03421577a08bc139daf7477a8cd5277b38ebedcce0353d28d89ff25d1f83fc6e424a372020a1276ad6ca01b3784a9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8e66a3ac64cbafa109b99cabaa344f3cd8708959c7e7d3df2fb2c0b655d17b58b1047a578dcf92c3ab9a3d29524ad4430dacf69147807381294abb793f116b3873e466513607d7f00f089f65fac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1788c435a2581866499914cb5fa30169303e04c2661ad1cd33d19166212d18f1836c9b2f830de4c575a1824a2899b67592a6eebb308cfd94cb205f9c90737dd59cd422c0227078b2caa4056cbed4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d91f0d65583cfaa8cc4c9a9cb93dd064b365b3839c43857cff8e988f814b2df188ed0dee486e3f5b64e14e713d1fa0ad142345cbae03995fe8c0a9dee5d9785a59389108037dcc0a805e11c32107;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4b3a96fcd2743621dd14968e8169fe5269211253e49a23c4c9c5e6e7d6bc080cdcff8e25dff486ea34bf52a6d0e3485d4f6a9adcde36e9e5deabd6ba4894f11fc2aa6f24bbee5a06dab06e7aa3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a96349cbb3972e5e05411b53f07e01108b97ee11283011915ea1652ccee3a875fd637f7fb20454e8be9bb792ea2c3b00629bb77c011f61c10abc96b25564dc9bde2f2afd520415d651c4600ff20;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c321b49f2ebd980e5adb05316859678c88eb9c8c64967e684b0aa303538b81d2362651cf0d0a31f0304c8fddf0ba7cad07bfdf3827dfffc120bca637b4a70b5b817ccd04e6e3607e7b51cf97f3d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88941835644bb56c0fc1dbde5e25c37b09120c209b43ce4b6b4c6e69506c8c1ac0db31fa39f3b465f3d1319aa652157754aca25e5cc30154d9b0f88af6e629da2a381d9084d2877865f56425f180;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb40652a3fd05157fb481d6ae50e4f05c8cfbecafd7b075b9d2bcb2c0c2832b03fd6a49d49c6fdec1304e0338098ff58f87d9a932e30ced1ed0a13ac33b16e3f982a74d8ca34e4fd66f1bfc0ffd06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9de297ae23dee2ec8d91c10ddc13feddf02091a4f25ad0e4dc6bdcb8927037e9dcc63cd959e345360e80d27908c51dc45bc5cd133722a0d4a0d315fb6efcd56f6c805afa72d17df769139bb3f80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaba380cbf8f51afd410bc978b93b8b919e3bf74d8c394fc77cb6c7c78ba627fa58ed24874c3cbf1f4291df87e8bcb2e066479c29fce0bb977d7c87f1b15ddb1cbfe2c6777ac26baffdfdaef6ca2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1025f74403d2fa3224172925d83b7bc076a863a38af083c6e184af995d8783e7c4bde5dc85c025e7fe75d4be8c5ae46ffe89b5f7f816683e04d1b8279dc0133a15b9601be70cf376079bdf22a11cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94214d7fbad06e5bb166a4cff6293cf424b0b9a2d50b78f79780ec7913820d225cfe709171331eefa4989fa0f00130948aeda4ca10bad4e65aa5fec9b5e31c78cbf0b7b64324b993d97641eb801b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he263213aa1ffc05ebc5765e15ad0b29f28cf26fb7e7a93195713c8db042a83882c311cdc21a9ea1f4233065723e88b5f06bd2ab11e724fa985475902ebfbd25bbfe35933e13f33afdb3174fe25a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f91d541a3195bd5e971f600d2e2ee58d7e0588d534d6cefa3c500b04f6ad5e5f467a951acc5c3e16214af8c521066b2f0075e8d68bb50c93ff67228ffed3eb1368a252befd819040dd84c55e9e0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18370043d57597c1411d8f5f554cd5a8d5a4e7eb06e0d99862156ab449c3763e1fe4bdfb366e20f53c307ce279be5bfc8ccbd457adbeb067eaff4eebc4eb42a8d6670e6c47954dfdd9e39ce86e368;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8635a94e1921766a414b8e23389fca6fa862733ddd4e348cd5d1b03cedc32006ffa14687cb00acfcbc6cf873b6c95072301de71215dab96d5234c55295c93fb3ba8dc4cca9eed58a6935dadd4b1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee99ca8dbb5076dde84a4f4e92d6c343f05de50d5260f0e5a917adb4db4bd44a51e03275c7761ff219b40340e1428246de1e910fc6ef1f3ec1ba0a751c1d33c496eb77afb07c7ec26386ba9ef569;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5b2bd271793864b7e31f61b9d93d2868900e10f9366eb10ca8d359f76e33b66e0dec361e036e9f4677d9c546fec1775bb8655ca59f36ee694119f3287fa45390ddb42626c4d9dd26d9dbe65cf61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8af2496a0130424d514c8b14f7aea354001f65692cbfb32e05b0976b23782695a3dc6df3bd128321628db3ea8eeaefc5410cc97afcd4aeceff18d5f77b442105916dedfe14f586eee9e990955631;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7f033932ee602fee30fcef0a8bc4ee5bb05a006df90055c5982f6b43308c7c5d6d49741ef881d16971137ae2516f9b015a2c1c5f245124e1fa6639e95f8ebcdb4193ead4679c5512f37b214086a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c6fffb011faf74a019cabc568abe0e8198ac4e3bb8c6d5b4cd82ad0ca911859c2972ba888e87b0ccb433e999f8f3fceb2801d76f789b59b23026b8c0b43e154fccffb563de9b54a0d70ef9eb61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152ce91a42bbcba88bc4a5e31435f3f7d5b3baafefcc051058d35d4699094e756a46a3331d5cf808dfe7346d38acc29a6e6ede517aaa9e5038bdec4b405515a05ebb30407ce2e2e9e7bbd5804848c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1facf7b6fef37c7c4c50ed6d81d61649fc088de57c92864fec0f442d06255b65b7b618035b035c5088ffa1650f37dd535f14c70e04851015c5269f284aa15a6216dcfc688884c7fa0a59e1f306cb3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7bf2a3035958d1563d409112f8491945acbee1ba88ad8da3be096c0adc254826eeab778b1b069f579684823dc60116ed3f5ae44eb94426f96dd7b1ee240fcbb26ad698cd983f52e08e758846439;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbf3f5739fa1c088fad6ea397683d4a95a5f4d77a340a29cc3986938dcfdbe30f953cd64033ffae9e831030d16379cf3067415113f57847acedc2a3ae043baa2962ffc851daef3fa2505c2328053;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d48bfc5ce09d9b2390755a4bca60856204979a2829eace067f7a29e11b60ce6333d4a055870ed68086113de024a9c5d240f99b0f6bb20968e82200b94b240a83f686f3c5c7a7714519b0f88f1d34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ea11911dd938d09d44bd585fced114de996fe273f7a5ec0da02ca24d64c856f1936aabf5ea3770368189f0dc9859702ec71b249570ed9ba19823e35182198d774dce660ac6e1af964480640bca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8c02df1319f3c1d0e14be31da61a9050c927129804299a18d4c553e7438029e7c16c0f355631a72b6c8954a3e18cf036d90fe62097d727c8b01adf474d3429f057e0905235646a958fca10f269c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h248c5031f9c7fae01348f5b8765fb4b75dc3221c79e17efcab86ceb2039f6ede5389da0f060c73fe978c59119ceffe43e00d2e98073c63caf1d2647afded597a3c029f9a029ccd43ad1247a5080f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27c965fd505731400206388996936340ee841fdb546a9a56726128865f89d9d54aa359fca439d529093bfd4dafbda06c71ce41541f0c3efdcb5fe8bac2e134091e860c10e3e38865a18f9985aa7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f44837bfbbf3e0751af256f4aa7743313f8e704b559ea1db042417191b6aae6635683d878258466af3e13506df1ddb6753181a78cbd950d41d996e085145b7d65fa540c37b492e6971ce8a9811ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e44413839d70ad8b84885c18fd10e09f18644cd989fe028e2c024e0c64c6d24dd239967c68477d9a6445184802bffb4e91246013c26111d49c89e15ac09c86c547c8fe6e082738d728bc53b977e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8e0776972402a81815f90df665497760d5d75e95da37533640ef3a38faec8515b82b956b065164a102eba38e4873ffc1dfe529c251d962a4b683dba6d5889344e19ae762f33d36fb03af6f9c6c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0c18d7d420613cb49e65239e58cfa019968ba9773d4700132c9cef599531c0ca4e55ac2c6ee1d539e8adf7eedf505ad89043fc118a8c73e06a45aa3c547fdbea6de23059baab7a7b19b47d16a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbe4703c3e4e0d6743462077387c8de2cb202d78fe13b290c939c428f9ca7a55e21965f73346aab067cce1191cb8f420afea91974f56ff35e9558e3f52b2d7eab8336c88795b8327a2740dc6e060;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cadb9130b37ca40c39a61a5fe676e24c3e61081285d1ce20caac334c6b1b246ec67269e517ac739207256a1c9bc94c51badf6366bba07319cfa702e03d09dca54c410e296b955dc118bd4376ba8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd379e21ea0bd535c9c1c680367c171757d85ad80d01d0d1b2d0235242680867cc3e8ede1f712669e8f85e847092c2713acac762f741bf0110798a60af6c1c947644d99d7cb5c83b412c8f659f626;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe547c5a63f8eedc424087a7b18516152964288705bfd728490f98a3d8def8af5c87efe26fc589fd4a84f6dbdf4323846190ec13321f84519ee72bece3bc5bb45f390bf8f6381403c1a5d2f76d99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2080e057c0aacb814584403cdc11d9bed5ce0ec3a05f67587623fdf64062bc67a58df3a294925406c1a7c62b236bfea8148ea8d3e28acd9481176f1ddf8516f7a4b69b6bb3ea65aa85996a4cebb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165c91482c3d47bea45ee9df6910fbd626628c6ed253ceb8c7f008c2c5d57687c4274d2bbcf00610f9a3fbcbc0648af578621f2a7b20737e4e676dcbcfd20417a0645e4beb92e997f1dde945960f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57b1ba94b32d894b0dfbc242db9e89d905de1e8f5b35c8e439e179c30139bbda18ebe74a6a465451c041fd6ff9687d8e6b5d7f288c964c1a9d28c7119d402ad9f99043575eefa201a0eedf8916c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1beac36f676e421a090fd07f76575043d492995fc4862985253644d65d5cb1335553e7e2a6d2dcc6d93e7652efffaf724b9e1683377f9524b84c89bce538fd4fcf4294d1b54c5746fb1587f45df6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda18f3efeadab032fc57fc348893c4afb586586665e077e11c789cce6ecff01209a223bc790e06e1d27b959526735ff4e392f62f1bad4398f6e109f2f48b84b8a807d60872e06898f0e8f738ff4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h641356a89f0f18995505fdd948d0f8739db852f5972e4c8f1ed934bc87e208ff2de48cf0caaac1ceacc5ecea9f3cd70b0dd97db4316e99926508edb570cae9650df01f2727ea597cc3cd85348b96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44f00858c6d4199d12b2e870f799ba052e23e9b9addcce5fe7432cf8f25952eb51b4a3506049bfc8764c2c73a0d0191729d5c691bc1d01c2e686df7e48a9ee09ca1647f54c88869521f5335f89c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0455ff7755ec51503e27713becd2a7d2d3ccd366eeccece3968f5845f7f034cb48b616741f1446d7decfa568a6b01f79aab998c2d9511bbb0b299ad019e4fd69ebff45288b278ca79e812c82935;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62ada6c537403b4f33dc40020826406808cb409cd074d4478dc834773b7076c37c1a34244acffe46b30ecddca81ef252b5bdd5db7bb10b0e398e32aa5519c5e596eca47e7412730d305010d8b962;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4fc4cff6845df20f368db84746a846aed95c9715f20388f593323ef6edcba05a7cf766e4753c921b24469e0d38aa114486f22983b88ab095ec15ed5a889ad6b99f611d91cc1ea81c426870dff4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32395e6302b9ee5b5faaf0727afd8d9fdf2407befebe143eac839a4aae9f1f95b7a61c5c00e86fe45c8909987f33472eeb13d67291a9e783192b0022b073f22dfb78c383c9b99a70e715455c8336;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd17a6e8a16e3fba749d762e82eb705cacaebac335d1b1256d71abca5c4851c7d1aa300cd0baee907653012ba7c1e8b4ee9621f31cc91eab772f5b7d7b3840ea23f6c6dc0d1429d52a0205e2e616;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0bf830bf4b656f247f2b23077f5d748d54c19419689cc36546fc16e2f7e00cb5d71d3091d30045f6de8f9c343af53c539e1d04b0ce3d38f28148883faeb053fd9020d9cebcc3975573ffb52cb6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1c09d17d07fcd4bea703eb08193d202c466f01218c18a1e086153bdcbc610c03b0b1a7a16a1a7ab6a40238947918c63edfede03414519c12d8e2d46ac0bfd4f625d4005292a3017f6584b95b74e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f3fc0f236a096ff28f6fd723717f0cabb81e48ad27fe00375f6fafeec6e4d2c9fd7a6169454a5007680223a55ca6ed756b88afa66bf86fbb82cd9081091c6f5f9299b48a51176b58928235238cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he708ecb2f3d704d45800335a3197e60ebbb1c6cd0ad751e4241b9da9db9ffe2fe2833f8eb6a3ed032ccef8d9cbb8b861f8be065e3898478fdf907b3507ed56467964f7494b5b1f9640d5f103fc22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2473d15b244e96260667ebae1a8f0d55c774a523216d01f1021be80b25b627e0a603950778cede53929a58300f3d20f611ad26d1c6c5ef22598adfa66b68e994110cde2a55fcb5687693858bdd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105cbaeaf3d44aa3e5c6342b0afed50df2931876edead0558a07bffaa1d2ad1dadf35df78b12ae861e736ea9b68a05db40f0b2581fa9b5f67d540a851d3f4227377b5997f2d1b7ea1986c8a6dffe0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28a3fbef1d7a4d1a8bc3a3b4375cf62c6848044f10a46cf6e3c469cc87cf5e9405080b66ba86a68f3ce13222f68bec3f7b9bc5c123a415ad9779e0eb3f8ab6e5f740d7ebf993d8fce71f720d353b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1546846cc1a7de66ab8682c4bd2e7bde32494f2f5e6c1e6d6800c7d44c1fa53436345fb2edef0a55ca45277af7bddd60ab8c20fca95a2186680939c3c19b545d3794fe36b303b0a4de506b17c8f1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha89f94b8a13f85a4c8429c9d1d61db9f74b8fe9fca27d16f163baf41901515325b21007bf54487f3a6ec6a753f8586b49709502d2b49c006c9063912f288bb9cc57a39878b1cae25809bcee27a95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h927b47b50f8d4ff10e2d8daafee6552eb7975d0d0026442797a2116b30524c9631d9a016bf10d99517e506d019cf894d6ab7ef89c083ea5fb7495d664de3311c156c03d55996ccc3c2fadb03a0db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f4799bc7032bfd60d3035228361ef3799e48d9ef69c115e3aaded22998594be08ba63c4b317cb5cc8f789f2690311197142962b78aadd69b0e03d4f4826a1c9c2bb81b47ced0e706af11d2eb63d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd5d071f914bb502d3f2f27f8e490f7c96c8b491a6288ef1978824775aeb4ad9a590db8594100a0bf8a5880409b6f798c57f0750964253ab97c8a0dd5c0811d5acf0461374c0355c361675d93bd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f7d196ddd3afe6f95f7cabb41b08c89aefcda70105eb353925adb31844405a61e6720ff7a4f63b3cabe9b6a71f85aba8f4195b742e9cd9da61706f9741949e2ffbe92133109ac0cc580f5db29db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133f00ab13043e3314ba2beccff065141c5a098abd2612c5ffd90f32c55215b0f5b6ec2ec55a75a474f02e45fcc4d22fb12ce3620d220b0d11193505cdd514f2b152bb9fd5dcec65c313ef559b372;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc81787e198d7cf6c9b1f1ea0d17b970ee9685db8c47e4acb6a4d15cb9ed413cd98ffc6acd0d8e804cca35c70434787f642efbbea141e0ee5e98c0655d42a92206311b533c72a155521a9386dbeca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h327a6e0568aebe1c405225ca49bf20c8b858b8593256842d666c4404a52edf1e4fe42e5c8208b1ea763adee06fd4bcb217a7ab138f72f4dc9bc16ab1c08a548cbf8f6afe973a097fc5fa132a9645;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb7f7a32e433cae054fbcd2e1c9479500390c3a2b3bcc6aa7fd52c44b73de1f0d70459a47c3f0270cdd6c87dd2a752d623ccaf6affce1fae79b441d674686cfe81039b372d0f3363a2f28fd3accf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1aa7c574d694f4b6f95b28998f558d8afbf4417383e209a7f6dd3feadc4872e9f0c053c3c2385b8e98ebe886cfaf69d3e87e0b52dcbfc427798333f85852ab74c311d3a8267b4810bd8d00314a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d07746a36eafa5906cb32c1724a70cc212a10fe9a4173ca8cc11b7d258e900b7bab863c3d591c8e6c51ed881d9e6462730812d5e4a3b52908d0aead9a1c0ad30cf3ba9faf8ba0a71d7856c4fb2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3bc10ffc9b9bb5e262f50b42a16ac9b18a91c89c0abce047fcc8365a0678bd450a7720db868961ab16142f80894745f4597d7b3a95544a5c1754bb64d58088b89e0dfa79a8d97ce91861a7a6f2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5da06d939cd3052b772042f53b40aaa6c78b1c9f8456ce9438aa7641810b6ba30ff22e0c6d355076a8aff68d9632af2afac5ad1d8a3243d61bac03da4981a0d5cf85a3d6d12045858669a294497b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12373e2383669c89cf2fc367700100aa123a859a879cfda616b11a14516ce22bd35797b48851b8357af2063e927b54dd282f0d8dc86753b0e91cfe37bbc8cb59a269b12938652a0e402093d58258;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b40420caad2c7424d18872dc52a15f609324f5111e2a3ceade00f936bf47adf6b543e47881de037b876f0962fc121f884d323b0a20be9196f76ed8086eafca3e9d25ea7b71499337f79f40d415a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e822f098fb00aaf1cfc9507d83154ed54b6eff2b86ea10da0d276ccc7115eef12bfa1e8ba8a982d6446ad15b658a26ed2ad25c96e83ac72f0920fb6655a47c46b11a38cbfd4e1b1ef703bcd45e43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee2023f064ffaaec203cd7544ef0c016a18ee60f85a09db04b9e5c4670fd7c03f748b42921c526bcbbad3f4b176dcc7f223f5895b980235d221f6ff0abc460235c7698ffb1b3c721a9ef9742dfe4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2d78133b9e7bfa9559ccedd5bc9088f560b1668cecda85c68254c8e0ab5d42e58dc13c8b75c8810cc73a2c0deaca0e1a1460aff48abd783aa9f16a87035260e3bef77633d6350ad5dd585a35bca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e984bbd5cd158dbb39d5aee73f9de7416f960b1477dcec7377f6601ea9a8d87bd3eb9a2d51d1edb8f3b6d101aa663fe043c80628d3e69531d2fceaa1e2f0286bd18365a3a7efa9b1dd170b4093a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c064fef9e6b9601dde3d474808ddd85f0b3def2c1e2324c2693b13c8f971d5f0547c58c209c5d4a2d71c52a678065b35a15764ea3f78e9a523929649515313c2f44299251afc6d441fd03cb84cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1062828125de0cafa1c90f3d3c27efb2486c1bc98a7436369c68b809f4771717c661dd3355502334ac9ac6404955d29241b428eebe8e0b1e0a244347b1c8c8c742b2bf04f50d7895626ce2628a2a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d62f2ab8170e32e5b5d835045397a27225b22bd8cc4b198fac5e93ea42f19e3308f19bcdfce51ae4f9808058ad4f0ce1d2015ad6db38a302e2c8c3264b157aed4bec68d0fc70665621ab930f2ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16163c145c01f8e4424067a5605b930faccc6c34149f286aa679a529a9d4956c5b680717fbcb95bbe0fa1851bc9b219dbef3aa0782786d31a9e80b28f3686ed0d59ec140b68cebd2c9116e5a7ecc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125ddbe160291398d13a539e9e0ae17cebae4127c923c4ab061c166d568cd03eeb26acf6290e2c345206c9f5eb7fd17870b81974c1a9112a1e5983738bc966475287006fab3f9fd1c4229219990e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85a6792ad9369cb48029f18ac8eae9c99b787427bfcb4eedac4dfec996e86c9ab2e5b9f97bee9cf4bdc508bd413e6fc5761db6ebbd1c08aa926ccf35b2421f8836206433458e91e8c45ebd6549a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e9f89e1a0a376771eb585c137d1cf8ec7158a3da5a65b602901668d42a82cf253159cc8531b81ee31a9ee87c9dbf8566a6e9ddca8eb108162168a4a22d1fc3dcee26c985ba85f31794dc96c7388;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10595c7d6c7402ff4e9aa5a81e7dacf94a671a1b82f3a5ac414e288eb23e7c93bdd28c6414b74d3c492768cb7390ba8b3abbaec5bb11b70b91a7c23baae63d3679085618a2f35ee98058012365ae9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc418489bc7e142a523d95a53b7339cae4e9fb9040d971782f551f7ee0fb7eb15d06035db344808c74e37d4291295483b2c3bbd2cfee2f20938841d51c4962041cf0f9b423a68bb34508ec23880a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb749082042433b4b11aa1f4dc62c944b7e8c10a315827c84aea2db295e1b721f345b919e9582eff54cf4c72b82dbcb32f6b2b281645c3876f4fcf55642fc1da9d782ec8f6072d439985775eedcc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bce3b9b6f57c8a6ad6d1dcbb37c36a956fbc5a3dd268a7694829c662d3dea4666d53e391802cbda66f86fce001545544bfbf36dccadecffd39d1b861c5a32aa1983f53451902bcd88ad23e2ca15c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31521e0906e54812f8d078481fe1b21859ad7c8108c22f4add8c99a2d01e9049832f97dade420a9319629a0eef91bcb32b8eb23aaebf80bcabce886e61dd086de0dd991a0e5076579a2f656f6d61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1130d6e6d53d7668286ac28a94f110b2cac52bf8126f386336c1bd80bbb0dd4aeaff5f5b0fcfff34650c91d31b09abcff697f8271275ba6d9810ca2d4924b62a6970fa53446c971fee6d41717487;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf326681353920c9a57cf9df9c01e6b29374d075b5f1340a187de7da986c907cfbad16a6dd8156da44bd70f29dc48e37faf2c7a0ddb5dc3560032b2884cb5e67b5cdb27d49cfac6009cbaae3d9bac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4ddc75560aaf19bae62eed67ab48d502d1aea11c9520fa29fca165ca4ed25efc453275a56afa80463cd1d72f3cae46ec4ab872de97f5e22d3edc15cc0da572544b2d1fa2b5ee907db7f8a7518d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1190012cad152a1cb607ae638f52a4e749b2486d8531c51503bd94683e1d62b729eedb5031b508876f0145ccf8478539256916b57eae8502f42eddb9372399fd4ec1b894209af836e65d2134d3316;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0efd0d6d426aab62aefc0bb628470519a0e43df8117a1997008abc7ab5a2acdd68a65d6e091245051bcbe10e388a0fc5c21c1c17eb501b6eb1d6e35292a5febd1bcc2e84c43c9d953c5d77a85ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f367a65545f5db4d2c44bd170f7db814664a868969511dc1e48067bcfb681a27829347cb65b00facc2517b0313c55d9455632fb1d1cffa28d228baabe4647761a87bf2cab67b9ea671f3902bc0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e63693ffdea496454191d2b9f91d124e2c7fb06b46a555aa8907d729dbeeaec9de48d82a6632c6db4abfe5a8aacaaaa6dc7d9dab63192cb6c01cb2b0161b37bb8fca1924c5aacade79a08affff8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc69cae2a3a4189d4cf47f7300ee38f8b7e1997f4e1fcee560f92bde8bbed921a40f267c008fc28241f6ad022b7624999ccdb6ca1decccd3c80b072b50d15a7d33a774d8ca1e969cf855945dd3739;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habafc1d611dc3024f39671af12b03779eb911238894dedc3d1ef876065dabb850c787ee528aa43bff6ec00a4d937a614d133183c3c4d2ed5ff9229fcdc87ae6a33cf199c43868cd0d79c664c0f67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89136df8e39f9dc29c0675dfc2c0e4f0ce14ca8dbf9a60dad2b4954463f7cae5fc72ef6ce8b5329f230e0154b3e0d86b5a2a4034c94c791c8bc705cabf7ff36fbdd576e85feb23870c99db8f01c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha12aeee2e6e9cbea9048a08e8e9d4f84b2157f3aaa5f62958df52bda6fc17dbee0d8ed13efd8a9907cb84bc4140401e2967bfcbf8123fe6c2d9dbc620d7e4efc888648eabbf8cbe25474a2128ca4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62aea14a1b6991374b718e9eeeb0d5f1c8855018e859250b8fd3dcae8c0c8de5840220358432b9041d997cb5c2066bc2a6483c6be06d7ddf8f203d5dac18418e660233be4bee6a6b18e543fd213c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1507b8c4d161a077ca878f17bf50f026e51b1b08c5a4b1b2dcf94dd815df84a92981b9b029f09b364f26b16bfa209385051833e37c84864bb0f597eede235bac5a05ffa2e6ddcc8cc2510c1249744;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19596f5496c9b693a6007acce838f48cb026a39c2c676db6143214a46d54c92373b78695507514df8295dc57e87eb24a5287e51149f82315fae22a77e75c31627fe23cfa2bb5791e65aecc586d139;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f74696fbe492b1f4213d4858aec8e217f5338b6afe4481089ea95869ba4df223e411085c394a9940029dd7e99c921db6f86bab12fd93ac99fb394b4effeb527ad2537fa77b9d6aa9e06e1c82ed0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16714ba475fda0a7fd1019409f4963c3d6f2da1ca9ef5d169724c5d396df50a674535880f6e62922ead1c9270b31cfa04e59a604f5f442507fd7236c4fece9b78cde2897ad7daa19ac3baa834bf3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1185a481e413a4df835d37d089e76edf1128a3413895f443319662db2d02e91b037d2e52af7c3b71a8b0e93cf9e2a86d3afae98cee068caef849db29b10581888bd44593c0f246e2f5178be1a22e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6876e25f2528734bbff4e9626349727ffb731da0b32e326b479a3b777c3e81a8f33730c3b5eae476f384cb3398a33a182e5cb91177f696505684ac84cabb7070d4cbf07e4439ee0d0f656a5080c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f49351b0405974f82ef6995b018b8f508de5122e240e88cfad358f833f35d333638ceadd2a15de4dc305914562aeaf28487ce7153ecf4fa88b57591b6a8f3d2b18cb6be43bf755969e0307c5ff3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187d5ba66857bc35f9c026b461669b4e227fbf1c677ab3e4f9174975be4a3d64b70f79594f33e7588f816bf7c0c9014f26a304ed7af135bb5327c6e4d5e1236c29a525a7591fa4dfcbdc97fd0e071;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0733e62a567aa76a2dd31ae3530d886e39215369c6642700e1d967228f0b5674d1b9a4f3ae483aacea7efc610c60331261a743c134e9924b6d001673ef2fe6d3a78cbd6dc0d724848913dbd9c7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c2205f1999caccdfeed440901f179882c3b2e7580ea6f50d2322ddf11e70b6ff43b77cc7271e3fc6f9a8b66ccce2b6f913b74d255839507ba6d7fe2ec5a08f97b6bc98f9671eedbe3d55b8d119b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1711ade1d607889c0a6e51e554407a0f2fa63640e36e2080a4a71ee962b746ef620ad197d8696e09fbbc7f42fe7951a66162828285f0d03a167e7ec23ca7a13796bb58c2902483355e0b69aff57a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ae470632689a35e9bbfc985e4f3909d467ae5476fd2c89b5364e82f68720a6c1dccddbaaf3047a15cbe0671b361b945345a51131ef502992bdadc61e28137ad5c15fc17ca9062425c2930df64b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175adb79c8e5fd7e4497e28b07fd0e6b710316cda839fed8f62bb01c72e3d7f7d9b8d516139a204459a963afd5f805f11434e7e133440c66b2db10a083b825115982093980f1db5ae9d06889316a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb73e3e55d9ed1ed149229139e794888c33bc5055f37b514984f94fd39248d3dd489bf6138a51404e00db8f8a4483df4f7d18bad53b462732543940e541839afe327fdcf449b84fc2650deb322c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h296575e671369a22e17ac36f6f7a87b0471d1b4e8ea01dc1eba8aceb77b80d0b40beb24f70ea61443bc22580f69da302e4fb354ab6042fd288eb6802b76c95bad11f54bbdc78b8a93ccd30db275a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13314e5aaf5033fa31dc16de2877d050f97c098468970303ef4bb6745458d85c151035eee37f5c1e8b739441e88e0fe529dff9565f8326f8fd81fd9f3fce6bd8a432aa086199d5feb02da418aefd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54e246245bae735aa6b4c9e46dab54c05c59618604afda23fd0f151cc2d7ef3ee1011f754bbe0f76aee1f41c6c7512af0bb2038400a8d98bd2deca2666295daa57e8b249c2f3da0973fc9b4f914c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf5eaf17e927e70bd8ddfb3ba219f1addd01377df972651da8de1ca591a97db502585572ba362ae2c2500c57373c04827a9165fe62be085585f67dd17f18f872c97cd419acbb6d5875e611f63302;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a43663afe7a16fd98ab6c23f35da49103c0a6b78dfa55258ed55c9cbbd7a0c199cebc8a69d8a5be3c40f4e08a64ab57d6152fcb1d4ed9834c4f44126d464f9daf1704376a0c6666ca41cbdcd1c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101b8fd29eedaec055ef59b60d6329b154f8108a9b031b1440fb34043c3bab8a47ac059690a137816393eb160b563fa90d7e44608941d6963249e160ff275abd573b3d6e917ee6835b183e6223437;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e188bc85d6f6b81a5f7f5bad0dea167902c7ff68ec6281b508ae8a32345cfd178d752ae226e41a84e81726ca66118e54f23a7f2a4a16ea47f2d5c495531bccc13c9a711bb814f8a8642d5303700;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e65b997e29510bd80022997ea6a7131544244acbf763c74acfe7b053c6cf75b9f48307f5fbdf2e5826c716abdc581d5b712dafaa501d934edd2925436dc305e5c5569f7c26aa365b3360e1740fb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e583dcd378c19ee5838ecc1eb3589254ef38ee866f285a63a57a7b6392be54e0e3517a50b69ff194ec3fb70f2aefa5699705d89d0bd55cd8df2df107b14e74ca84883317235046800adf58c84db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e5878a5d14662e7d0fe1a9a7d29151cc9cf1103d0ab6bb59000d572fe5aa3c91c35bf4819d62366c422e8f7e94b25c689277a7848ca94dda2db99530beb128c534fc24c0e25c3dcd9c19eab2fb9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3b839d3b6e180181f3efd584a028fe3dfccadf7cdd041efdee77a9e9650e3f15efb2ba3c5e9c6dcf30b221013fed9e9020aabb46e6cbf16ccb7cdbf06de6e9a9e0de961c6a6e4f8ddc8bf0b276f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e6e7ee0c6e824c8c9aac9c3e6fd80a0f04926c1d7f5b3da8174e3e98a63e538329fdc5df1896880f26a1e29e5ec2a359bc87b44dd0f9c865d658a12b55a98a03dbf0b5a89ee3941e2b858bcd993;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93f800b54cfa7cb24c11870b920e50d37dab533d4b8dd4a17e8899899c59d9929e92faab2361ddbbf00ffd00a504a8fb399a0a3139d5289c50372cd0a7bb2cfb66d8eb9ed03853b45769d7ea5742;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bd7c66d4f12880cb20d3f2dd8cc25976413dfebdb99db35625d1cf5145b2c9766476adbb95e85f8d32e9cff4b5a353cc431126222e4a2eb81aead9995c9b2701e909e3305db40596aed1941521d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e7837306f201b54eb387d792d2dde85673645fe6f1722f5975ed1698ae26f0bacea3494ca42693fc96eb0827422cd455d07eeffc3b6fd22f067ee8722cdbe8d73979590d33b247a6bd254047279;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72612f25cec00baf70fbba0f3a943d975a35bd8bacd40c296a6a70b417c2e068d0fa80f3285c48f6c869cca4a983883aa3d4792fcc2778f0bab7fb17d4b9cce68db63358e35a7b7fc29f5c36d8ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a31da7eb151176db5a0bbcafeb60400c0cc7f4c05c0240f756f89cdf823a69872dead940c5ec2d4d241f7a85a21ffdf87b0e37d3b26d7d588c7e6fd6994a5253172e392cb4f1d9e34c020390442;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h440b251b4dd42ec231729373564630fcfced3f072b6492113c5c76610f0d0ad5332eb15889f0650050924f7d5b48977a11f58b7fcae1790badc3c3d65d519d885f142292fd5a5d7c1320b7d326cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0a4dcfd769a6431296e587f1c44d3cb99fd36b739f43f7cdf238abe3ab348d440137957bb1432a6fa50079346300a61e4c46321bc5aeec3afda86eee7ec47669b98a968f01752844ca4b178ceb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h245244bb0d9de771362b493aed63ba07eb4a82bd8fd25de36d25c4346fa93f54eb27b6cdb4179665e47c5cf052bb84701d83091b7cffe9c6320ebdd16a36fd06dbb02a0dedb7af208906ce2dab54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c13c75cb3697bef112b19365c877417c7c3371441b09022d30ec3bfd845a990c8313e70687fa499e7bc922adab8fe006ac7435f61724e8a33c14674f5dea89c6250d3aaf978b5d304639d9d5289b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ac849a3702a67caab0e88769c61cee75cddb48c2b544eaca7b18b4d9cb27d596e4fd0178bf66377457fb3de74cf992bb2db9eb30ba7dbf0c849f66e286b662e7c442e266805e5de72dba3bea4d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f657d2c6971d46ae2732b932f470f0f6740ea548cd17044eb825144f1554c5a9fd36c06c1b6468289471c0dc8b967ec95d1887ada25eadb272a385d686d210c3044d60b6af810f30b249afdf35d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da985030e68452e31b38c2231ff12437f625764f623f60b3d241b47fe986be198b1a45ccb8ec7467cdfbd394bf176f9b38b3e5a35fed05fa7f7c05aca04d9884390efbeb9b5a32c83b5adea3e95a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53a00021a82f2830f677dd0b4717e58e0ad9b19ea4e432fa57a938982bd7a92ea84cd3b2fe0b4712463f71f1a3a8f7b863f70fb29bcb7e0bb57ab055020634bd10eae2a3661fdd9ccfca33472d85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae77818fbb41b78688629bb714422b09ac9c3a08a18f2503baed12fcbae2532c0ac996b0cea6dc8c7574f1e2fc872fc516c110cd90c8cc41e385e567a5229c3262978dd38b3caaf758fac3457986;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfffdf13797a73096731fbce72a437fea79193f2a67387ff916ee3eb73184aa3a4adc1076c4a8091b4b2d74633172eadb66e2d2899b47f9e45c64ef3ae02938365a8e7507e9df0f40bb8c864a5872;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfabeeb9e5b30e101340b15101c0edae1ab0ca6e4f8875c115b8b901a2950b4da7359343eafd9a0f4969c834a9f00cf802d3bfd65a79741e5330ca784369862b1f79c93e9717c4dc7d973f85adf95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e532e470da7ffe8568fa2f7b183cc307f4f462280877759ea18f580ec3639eb643572ad0ab31c385bf41b81ea73d36e76850734b7b5891975358e209a3fb84d3889d205a4dd436629a3faf7a83d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15eadf810db339dad2772209b3a888a541cb79edae9f12bd01bb854a141bb09af3108a5a1b0c019f647d3fa5da110bf1ce0199f164ad34d002247a3e6d9597e75d28c88389ccc1b99af63f90c8943;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1519f027fe8d190410bc7fe207ff1754ec48bf0d6be7b72cad631f1f2d4ef3843aa4c51e384e25f03d2a7c870e0fb452b308fa3677bb48d4b8b845726d9344ac8422bfb127c222e1eed3cf2b67874;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbbfe373305a9caddf88b40051a7593fb1e885cb4adf65298298a21d90becef9f5723da520c4340c85d4f17da2b7c922262d9295a22bf622db822ea5f5d09a8e713db64569983a64c0a130fbe37c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4dfd4a4ba230b662240fb54bb92a90cd04a33a50c70db0a5ec7882ee09db67787a2c8980af68844e94fe9ec6edac9fb0286417cfab3fde6bea02e1ad263cd88f07c9ecb99667c0ba2a8a0b167215;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f3029d7f2de58b3bd88cc0daf23fdfc933ec8dfdb9ebe36cbd14e66457942f7520aa10d540467056c1df9407e05cd32aaf2290395de654ed95cf03654ab35e88ffc91fd30d237b52d181fdb55c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fd675658c1f4530d6e4fe7edeb868a1cb86d9d925266550eeb3b582a8ae9b09e274a28645fdf60f4a7f6412dd82703ceaf7929cf7c552ae6ba5681624b1a5d3d7313606ba7006a20dd7578f9a2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130efc45b17929ea902ab499a082bca7cc877d668b7c681c8923f69079dbc8e2a9c3426336971a453593d4fd7e5234618a0542b1daea51cd24115bc95b3e35e69f8b773258f38a6a19190572ea445;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19619e104301f2844e085e970a1ec515889d0488d3e5717a0e59838a0f343543db9298263466d0162b19b4c6706003b72e90c3b098748e25eb59e617e796318e7e4c9dc8c657c9a8581be7ad5afe8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c97e615aa6349d05e92bfe8e9b55c93841b05fcc3e1c3e311c766001be65efc930357683a59f9c6206cb460fa34918a3b9a2fbcbe65d55397e4c2a4fe35ad3bf21445afba036bba9b68bac510b16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e9bcfe996e102d740a09732a43f3263361a69fc1549182c3361e111b43005d6184f64380d40266bd2dbd05d4b7b4e7042253e661cdedf2e3db98c36496e55dc52f64c579980bdaade254d56cc08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e20e83ce0e2a3a7ecd953979d0b93dcbc2cb4252893000148924e33e6e0f75f74c588c41adad5a79e3d433e42370d0d1c5a6e7ed08ce41224465763cee53f958bc975f7c0ff323e633b02d9d1fdf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8d0c63391c86898d94de0bf0095ef66c4d8529baf701f23a060ca814a9561f01fee40caf16d92feea00919b7679bbfd2cab61d6b19c5610f7244c13bee6b8e030579c1a7ff173abed54cc15b8b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e14be84207a1a4feed3a8867b0712e846fdead13aa345348d065d540fda703751ae0e21a5ef49e1dfd1bbf5dd82cf9628eaec0d08f9047562518b78ac89446d5ead502d05e38ff66f3986e384a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcb94d6efec2362deadf149ce2e66bdac808a86a2827ba078a99860e43f03d1a9aa79413a5f10a97d5a17242ffdcbc4ed83ef132f31271d62d0933adbc642d57c12118a6d00b4670d63478af50f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181f4a74c23f354abf11c05b6b3df7147aa937c4f1d473f550e925b62583a529197c6b26de7af4e537f3f949bd47db82aff88a9b62e859ce48ba4627ab08846f6687bef81e1d9849e5d242f5340de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebfc9a6a382fb7f1018e52f6ce64c9825afb9b775424ce34b9c274083103c4ee5f3c4102a9a5bcac9ac1f6b75065ef0604c057bf416d4f3683d760c300bccd6af83df5514a48d7a2192c67687903;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126492c2eff539e16d1ba8ba304d2cc3628754891af0f1df01813cf246e5108a74df0650b6fbf22a9d251b30282c330576ad09c4dcff3fe68a925d487b752f40e15d48212a908114637f920e678eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13da434d853f3cdf7f00edf31775ebdf52b24e5f00fc5b210ed841cc72aaee38b8bdbbb0ca798b12b7d6a1e4695fe9c1d9236449e47b8c81640a45f8e528ece9292f1a61640942435f33cca56900b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2962f48e67a4bc11371d1aacd52e0bb605c34ac1b7752a8930dbfce4e341f7fb6e8c7d2b6e1ce226ef88cff513108810cbf8c3395d523d04232185a51f8f13285bedf8d6371ca5f38a33a2efc94f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15aa646f9c2452dbfb04bbc9338f76ffe129de83f70003d3313950d1396342407aa62dfd5fd96f64c66eca42047ea5f83675cf982dda0e9d0f9f24d0394700ce91c664228a3924430ce6c442ac3a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc18d861fd344fd0d3e997b59f6a7dc6bb4e86361f9df33b12cf74448e9babb814c941b8ff47b19774ba77c82f35b7d7c2aef6c05fcbb89a1a626e1829bae62403afb07f3778bb622f8adc9cbf68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aec61f26e79e77a35acfb707cf3797b007c7eae5b323bfa2c0c1041796c5923eff1a688c44fd96fbd9806b77c24d7299574fe1c8d2873e8fea52611fc045e201a79146e0f8607c6ee9f9e28cdcb7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9922510aca89fd3c1f79a64e6c60bfbaadd4f086e2e94deb4ab73f6d6629c2a2a41fae5be9f0f07b63ec90323e3bb96cd7ff49689a648d9af04fbbd4b13a69e10c429a59be2b26403863b49d3345;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb86a8d6aaa6591df63cd1f9d8637f44f71d52788eb631f2039f5e8b18120b9fd741b6ce2db0e301441fe8c0e41364506f4453c6905e83871450028f166ca2872ed66cb248390ca88944bebd1f4c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb8527d5f93894253bb796625463987af7ad35d9626fd4fe5eaf4b9881d95d302c6159aeb778c3cee4912c9d91c84c075303837cbc2c50413a84b6590cba486214305586344855072425a80a466;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114101176121103bf8239cf74240e9231bfd00ecc11c225e232d50e5e788a8d8e89bb0b39c90871143f8743cf632d7bde27eeef6671a7183ce46f03a8f7f2e15528f7acc797e13998e03a3d437412;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16feadc8f4305f9a002a18f18accc2741fb0f50495269fb30e5b6be991af9231f29c0b23e87ea722de5cce22f578bc2d6f6008177b07eb39fe90d966ca097cf8b665b6d139be2caf585c43ba17db5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12798c90df563695ead1eb7ea238180fb8b64c805a21749afe56167b0fb5c18d7a68f3322969a394ffeab1084d6bada37cc0e1149340a8f0cc69c9cc65dec11d59c177eaa41af1bc1a64cec852c46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c93ec26f27b2473565ef41e092c82ff9f358e23bd57f80a0c0994436660ee7d65a93fb72f8924a18489ac547e08690b363fb4a29eb0187c34d629742b7117b13821b408b5fa4833daf116f459fed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc4db50941dea7cf0145267ddeaac7f54063c029ab95a9dab416ed7c34c6a0542fe8c8ce87927288f51a38389fd00194b256e234820703ce6f98733d6c0239ecdb5eb1d00ea7e02cd79aab88eb44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1620b9110903354975687aa6de0886fd6d6741cd09da48999fc107e029f745c6827308b841efa3c9ba6c51fccbf55a18fdcf9a8c489492108410d8565350fe7bb2051e0553d8811a2337847b9721;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7180bee67a36d2ff1f1ec22b44f83bfd507b266d93e191bde800719ea5d9dbb1ef94ceec22c8d65824d46789659efd98c16ab6ae03ab79d40c2fabdd48148619b69a36761d8957a9951f9c1975f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf26f778226c94895abc6a7ffa325fa5d08490c42ff0ae743f2a33323d009dfd6b65e86f31daae788bea1a6294e415771a52feeddb0ce6d7256fa7a25b75f83408202acd3b56fa49ed2cc2b31d577;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d7e0e2987cf44611622f0c9adcdb08e0786ef43a28d7950a4a92833760bb57909d869b60f69192eb65323140696e91b538ed46252cfea922d77d9f5ebe84a2edc20badccc4d5ce02c24f36f6ca1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfe2570ced5ae1a242eeecfcb4ff6e038ab0b500b29d3e5de0be9361c3f0f11683aad5a6375bdb570b4425fcc48e40e706bedb604a673a7014e344ce86d74d5ae8c8bc6911991dfb6a8845c66e48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1569219f7d8e23f711379fd8f505b02bbc2142d8ca7b1bbcf6d3e295cacf39390617aa6596496acd636f3cee0e45476dab5aea9c1a9314ef84511851a145da561af5ca01b560d5dbe3ee2319eb6f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d5283e85bc7913a845908e291722294c6ad393c0d9d67796becfc76fd4c59a83557d7538f2748ba379f6f5d47564641e60d00a73c46ca563d87d327e2dca7b343dd5e62bc93fac66e1334ae1db2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ee14160a87a12125723c3740b7688849ba1863f02f40afb4c99efdb1fd37140646a1aa6e9e2044f5a41b2e726c4ea18be7e0712efb12174b7d705bf87bc472fa3fa7ae6719f38bb079f63180f5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6dc53de73da2b96d8e11a95c88bb32ba6efb3afc21eddd856230bbd336d50368af19f143b9d11e7439c8d4eba11d0378b033aa33fe358ef25d9ccd9c21048c25433a6c2423c08bc90d01fbbfe0fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbef335ac79e82620b0abefdad427b0b924e183cfa158494793551f2239024e9659fc4d4405144dd2e578ace0f21fb64b69b66bf7e448e99a869dc0d0df9ccad1317aa453e918a9a592118bb18283;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b90a05f1593a89fded0efcf77917390708b68fadeb3720f746345427efd9915c78d7f07faf6634b09c6fb1a381ba94c1be5bb2acf6332a71d738541f047979b4042cf437ff3620be3c623e42cb5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126c365b05c68ce4d0162a49248fa6dac428f5c7f027d67163d6ac37c9b3760fb454707cd71dc97ca32b57b2670c4ce2805710591c7305dd36b154a69f116362362f8fce3314570e3ee872377560c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150645e675ef65b52cf71d967be9d6fa5aa55691e1b44ba2f437422ec4bb79d6d9020d710fc8c9245043c9418e815b196023f63eaca396bfa43cc6b5ef44cf0c0a48a97efffb5fa2b718cc50dc01f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77222ad7afc03662bf954b081ea0657f50ae2c88042df26a1536f2369bdb586978efb60e3f2294ae37c822019b0d1eb7b910708b95ca63f3b321b3ad6a3d87f06eac1737230be3f622ad022bc752;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ef96d2d9aa438a9a018b70aab9c0c6dbdc10d6c56246bb211d8b6afd7f2506ba017e71a92584f40a93322d4695f4a7fa9c54ed2f0dc98e1f6c55e52ea072c56aec10668c0c2909c9412697438e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea87c1cd30e8387f20f735bdcee37e7d2582d6e095307d7936c923a3f00fd0c85159b5506d1161af0b6dac379a3af96dc984c8b6100218944018e2a66fe0966906926bbf22e35679fa57d0e60463;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b633c067b4f1782e9eff6a1bfa9fbe97e9e3a74660974c7961f6dfb7a5776731a8522faa26637b0f9714bcc4596836c810241bac3257676b96896d7a720b51f2fa37e09d911c75acf611b6eb566;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1727a3d330588d9b8a01b968cef072e6301d141852ad80003cb1f5edb2b143d832b8667d7d5750a4384d4972608a4f9cd497ccddbf9f18a576b5ae52c5cb4c0fb1e0a5c99d61cb450c61a38633388;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb80b03d89cee2a73d74394609de540850c0395c12fe708c71ca45a98cb41bb2b9c52f8833c0067621073442ca64d5d17fe6ee91ce55c95f5a8992cc3d7d065c2f95a93b19d1b7e6663d75c299ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90af7f22ab0e0f8383cd42dbd7cc43bec30c020b4ca180ec2fcade88fbc227a9cc557ae22e3e96f9fa28e81b561251bf8b619042890f60ad80ac7cd9f89d914fa26fb6633ce08f81af9d7724339d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5867eb30202ea9c5fb62af90dd374e405913b9cb4874506c6cf83fc239252a36143b7b3daaeb70a7b1c4eb5910f962319b529a3ce199ded7bc643d604d2986515ba2f693b00d9b842041252261d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c6c9326e9becbd5823b39dbe49addf551a6895f57f5e03b875b371153660f30d11dc4486ce955ce53a77b154e4622e945dde636e12d101e5f6166677cc958e236293f62aeef35f86edd40fb3f05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10560816dc1a8694095f2ed3c62d47020c3e28eb2070d67a1365e9999bad34a467f60cf644f1bdc783c8def89319d591814ee47f08d43c70613f09442468babdc6ca6ff5fa5e694d6e460285fdeb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1403962874aa11db301acc02a1e4101509d922d3d843048ea630f79bdcb6103a9e83b9f70e04af0c73dc070fe944937ad60afa2d6f8f230c9e7b9bc6143d834b0f6e4dd1ceab389209f4de5efc264;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8f19d8cf93a947fb04f1e88a10b26efda0ee085ac155e949da050442adaf3a06928172063c525d8998b636ab9d12f8c5f0007a68a752478d51b27e86393615db5bcc98b840ae8a25bf8384e11d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f57c764a772f8a252884b34f45962b960abc493efbce1bc335194ae327cc6b8fa51a4516ce7d911508927b5a1eafaca1821feca7b62a28b6554d4f88c75075f248e94ad3b80df931893cffca26c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28de10ee10a717d2765bbba0fadf5ef70ab0734184ff36f4f76b011f67e3805d246f2d65191a24eefe5f4562aa35a425e3e5972957736b926648802deeefa8b912e2518e365298121cd0a0e83daf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fdc6193478147dde6c6221a5828d03693e05d242a347ec89553a955a879bf1d528c6de16b07a97bacff9cdc5dc861ac25449d05fdf2d396d4aa9d3fab99e40f06f807034f7d668b0d6534ad1736;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee2de27cde1d69f5f985a06bafd45ac8816d3880b12c7457f1cab5c84e2fe3521e729dddbe86aba3ade780ab9775e5d0a9a55a00381a02372e2000a6c44f57aedf8631f428e8a7759bd8481acf53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68c3eb2e5883ed3626228942b1658dd93381c7cda366d28b943618486e508e9bebd54e8bcef114a2e2e84682e7535d817ac38720c5c56d8aa36a3c818cac18649231a04d7d5dd4452fbad17987c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1473de406d9f618c324519d2d076345068ca84d35d4ef2c7bab20a7ee052c9c3c692a412b2bf2a2e1309d924b7bc40089e04977903aca9105dd26071170495113ebb019eaed17780695418bd3a6de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105c2c0ead491d52cc72936edd3541c0a4da2fe5fbf76c48d8da9ff245aafaadd29953a278c773c70f03c019f3fe790d00c0b333b8fa86799f8e795d750fd593ab27f681994e012fecdfaac5fbcbd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b24cc7e04a2afd8058bb5de123ebce543b9ad47caf87b6a368be6eec2d36d1035385974987f3d38fbb1cca5675661ac6556d1dd26a07e670bc85fa8440efed1dd4f3e1acada4943374d7795b42da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb78d16d3db9699e876fdada06a3236beb6315b6368cf413b2409ff646af8d3db11cd35e304b64dda4fa358c47c90b661338f090f8430658ccc89ee8e3eb1b50565ef215b742354c26bf43bfa5fed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c95098f26f9ba988fe34bca33e86f03a8a3017ef5f120fd4420db92d3446130bc90dcf14887f575596b1e4f946e96a1cb646339b80552af80879c244799220d527f0bed8b9921f72118518453454;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122c3694d00f883bb98ceb30f875242d49d118975373eb3d6663ec74c6d38b92e79b8c33f2fe3ba175af215e7f42e12b0b36dee3dc518fd3e73a5ae983dc016350a24f8462d3c3397b473660bd4b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1507dfca917504221c3eec9a449c0cba2e997de0fcee1d836428a3f22fd235affc6696bf3052230f6a207113dcce31c2400b0979f2c866b88f3ba27275b67da9af6f06c018f624462424467ba74b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5e163595a92bfe2ea13edc3903e6f858771592a674daf6595b8973ffa292de41ca919c788e359cfa5b7d1def4046bef5b0f490f3e0fb3b6939b71491029d41c0f2ebdabc97629883429be62af0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f50111abb6df05b55fdc4f718b3be1bd780a198f98fa9c1d4fe99ba32c33cbeeead22752d62cd49e126d33183ef72751d39db0e710eb197cf1c05f3fda3099c6d298d68a58c81da7ab71a0d1ee0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7d50c3e3fac3bd845542159a2d5a931872cfa1611d3f272c16e37065c161b18322e13b0bd1ed51ca48d875f50ef0be119c05a1514e2e420220030ac221cf74ae6cd7d775b1e541896b9c4256592;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1505c20a5216db9dde19691f2d13e1bc5d8e5f5498fd1ae9633a2b75dd72d2c36e08c4bec0eac872f9d944a559d4e4e2ca330d078cf54a16de8305f97ece90562e032c58acb74f2f2003f422c964c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78e90594cac58bf16ead40d33cb9b24d21794d4c2ecd08c0a64ee0b1eb3ad34cb0bbba84fa3c84ae3d9e9cb1c31a1c87b5cd8f0c2691ca11b283f36901737269ac3ec3cf1d213ac75c4de5af10d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78791376ac457d6d734f2a7c2a72d9732000f97c3a97f21db78199328d536ddbbd734468e83f4279eaba266bc14539a1d3f829599e39d7faa4bbdf1bdbb84716840449bca08031f72a6c9288f526;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8682168f0c4b861e5c5510ce98fc6efb4ae3ce9a5e52bdb813a58d72832d69bf19e7efc4ee48658e0831d6821fdcd7d0f393350d5c4854c4bed101d6ff507d02d781321ce7fcfc42b955d5b9fc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164afc64c261091244d76970050bf903faa9a125d33a8c2b22d44f5a82f326f5aa8ce826cc12e430f12555815eeac659cc84fbd97ea15fab8b891a482b2421ebdcecc5c588a1fe3638ad38fa1f5ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce89cf6cdcc38cb01a10fa7583181d34efc0c9b8464c716724c23e0be6ac3441272e954f77f42b54dbe630bebd85d78c06c62574f46d44a936aedc3d808033c0fc7c80ced6f87d249fc38f9cbfa4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h882cd1d2ba8e8266651f70cce37ac0f3db94d4529d8bc7190cd1621cc98c317a14b7b062c9407375136b6a172b2c86f07046bf24e5dd36ab987d5a032f9a6ce476b741b1ef833ea1ed2af20bea9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6218c37655c7a03c911449f2fc2c417a89aaf44f82bdfca25f7a6277ec293ea1d7567bcc165309c1d6af412982d86051b0132bce63f5f9d090b29f7739188258a5ecb563fb26f91c5f40db4d328;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b5eb46c8e7c6506898ca4ed102e025c998bd326380a1a06ecd7bb25f36b291f5c73a083aedf7f0d7e3ad80e71ede644ba187b21c8d4cd5ac5171df003b13225a8ad15bd7ff8375ef30788506c01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e005179dc5917b8cc04e964bc69855e232a1684a56dfd1deffc749d79d137f3ef4b9f9921312dd5d93f3b88f79db97f9d609d23fa6bb13dfcb414b1689ab0d23fc045358989d9fe91d533af0dff3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30aaf2b65e3c266e0fc7121e5e95c1b2ed47085026704483df1a30ad3d9d68a6c12ed39a8e1b2c19cade6a54283baced5a02efe94e3ce6869d05b5413b9880800ccaa69ba4b9089a136f2bd9dd11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119c0bc267a64a9268542472046e4906d4a89f8c375cb2b9efaa207719eb0d487a3b414cab1c08e2ca2f26d2a16ed5ea218ca13db394fc25795b0085a6ce31aa870ae1c161b1eb48d5a67f6db28c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba779ae62c279e701efb138f3091ab77a4ddb6c9d0263dc27cd1f992f0b4779b780c45cd4840b388e2a0de9510ecfe6799b4f253af7a6dd0188f9a2012adbb22cb71fda954fea83fee19d2f2b8e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1239bd7bb6dd32b287dfbe91e3b4d8d755df4bf294b1a5d911d1b6cb398e69ca2de3c034bfb02e9531c035e82f4887271c1cb7bfdef317b91373518356fc682e03e647b9b5686215f12d44d43ea1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38ece4961c4536e5aea1295417ece4865cbe29602bac8ded441aef21b2b70bdf032620703ce63925a70615647842de3f6950a6b1dfa77dd9e24248a77f8c7e82fed0e83eed2b1a65a69c3f45ae08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7574ce747f727042e0177ba9cd1a8a05ca567920f071be8ea2c7911f9aa4dddaedd645e08c6b226092b21e06e4795f36d5fc0360573602470197bc170ae8f7735430725552b86aa01fae1484ae75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b546e5ac05c1dce52745465f513c4c941e40c6525edae5d03cca2ce7572a6716323cda1e30a0545ee9d7d352760bf88c8a5fcd39dc0466a7cfc2c18a0263671d27d6f86ca55768903390b4eaa421;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb700e87f5e272b45456e75a334df8896afd4af13b38a820abdc55d5d8a0df002f25fcaf1f55b65c409304d81e91a5b2d3949a731c8d0ab91774ea4122d3d4fabe9940129117c3e31393033e3e85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd367cc5ae60b58ae01e80ae953f50bf2bf1b9fdd92c5d522fd93c33407aa537171e80bb4f3603e30acf0f2b5d992451b35e9ab76d6b588753358b3ab768f741d3b67fa98de49afafcf01c4d2e4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e7f4334d8d7ab830e8a4cad5febd8d870edd808bd90f52d366412302e047bfe566cb75e0959bd1bf582af6535a72d012a812fd1cab309b70c3a674f24af694af923ffeb0231f95c6ea746644812;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e9a36534937154930510d20460e139c156c40a4b7d668ef6cef4079a96b456fe6854dc22597d54ae509331e99dad8f118c9af3453ac444b878240843e1c613bd4cefd458ba4803b8a3ed856379b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d3f7e59761b1d5e5755c3b8341691b851cf53afa746e9c5b05e16c80ed6be9b1a70e61b2738b18e1a14eea3e8c848dabee4037b477cf10464188d5231f51e2afedccb1e77839da818c361975e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h697111990958f863b4887449586557ce2d3294aae81c308353b819ad343a62ddcd5469cbc88471220bc218db97937e2c20900e5d5d1384cde5aa5b54184fac0dd9792f80ac18fc4661c99af100f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163abe50813d8cbce070d41753eaca2b3e6b0a99826048fb27f847e4c6e4ce4ff1311e455e0c78598b9992299f1a6bc181f85b153c788ae70a5b78e8d6d4a36a4635a3fabfc7546e7333eefd6ddee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146da72059669fc371adb0aa76a0ae6cbb758ef82c71da58157960397698848f93d6ba7763429e06656b6976bf7a799a65736b116e90f0b1626849f2cbbbc5aa90b95a449df5658ff345ddc8ed4c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c9f048d4b31a1fbfdbb18257dfdf1bd690734362694f8ff14eb618d0b1caf4ac2a511fd1ee4f6d371edbce16a2af724c90bdc78130d8031af780e49760b0062d7734a854e2dd89ebc02f93ee22a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e86560b58d26221b59adb6f1702eb6708b06f44ae51d42704a4e68e1ddcd51d61dd3dde99ebdf34ba00be22f7b705c205f75053a602b5fd4b4e4142d4110e19172554552b0abbf6085cfbe8cabf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15dcbcbb108173e19f89c1ed3bca9559249225a54e27863cace60dffe5087e06f226d5f0f1e3a0782dc8afc28939fb3a8c99efaee3ae7c55c6db4195cde314d364fc17672ee8ef1594e7f78c2bbd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b38dc7361c4a32912dae2499468ac1cddbf3f183b7fa4e280943104f4b72b46395b9435b31aa4bd19a25c29b60be9db8fbbc7367622324a1d7e68348aa357d0a115b793ff008e3d3e29b70effce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12aa4aebac3971f0d16bc6bf5304009337590ba1cb128ae9fd9ad44f984b4fbd4a0ad250be48a5e46bf990c9da9401b197a288ac75034aed921e215c25959d24066b3c109e7681a0233b1b244ebb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba734fde99ecbaee1e545678c303c8aad18b71e84f322fc2e3f17a0780ab72e63ec61d857bbdf5326fb664e80da97c2e2ce698cf7a4e947e4f875a48b6dac46d54bd7d0d5f985bc23cba1150095;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd533c03676b15ea90c5472227d3ca5c07ecb01d848b5b93101602e81b9c6b6f3c5a50f7f5c45ac279d3be4d6b841ff331b5f4b42b70a7243cc02e1d5e9453b690eb924811c029c54e7b19f0d87ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21623e23aebdeeb845ac6d9d9c49584b08799926aedf14c44521632bb6a8da9c72b7e771bcc858e799feadd84fb7c5c3a881848bdf3ae47a308ece275d46e02ef74a65b5a589a4c58dd4bb67444c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65a0b1b7835808f139c96b00735519bd6edbcdc022ba30ac6d0df0cc01e58ffdcdf1f0819924f01da338582c6972bd77422bf1787089f6355ec4919a2214b4be0857b23a6d357d35e714bc841a16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0313bcffeeae495bfb52788c98ea579aab9e5e577e438b22cb5ebe51b88c50f72cc497c8376d3ca13832a879f02f1116fbd1788d990142341baed2d44320a9c97cf041d3fe3b8c1a585aa376901;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ea73d30df994fa9119cddd430b710bce42c4f8abe2d2ef691c458248b920acd1447a32eb494a904b3158ef0c54065529dd57e2d430e5430deb7f2bb9f22ad87654b9cce230311025c457d27272c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d7add9913bae32f1cd767a1da434b1ce36493b41387b5b31655271ff1056d8f4165f97f3f180cb9135457bbc5d1dbdfe80c60902033fb4193961b7c463f289d022be9c5aa322edcb883b54c8fa5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f3696e05e37802ab8224367ae3e33b5d95f3da934c8dfa1a7fdd30b79c3a991404d3e87317a700bca96ea84c84fde5bdfc5972c5942f899e03329f606887ec8022492062f4430ab35ddd648dbc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8db18ce54fc4e44b790ed5f2b5ac874abe713910da45d50ecafba8b3fd2c747e94749427c01382a7fd62bf8a4b161d271d6f29ff6df99a9514d44ee2d53a650fe2de961cb5e80c564874561e466a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b4d17d205b76cb17bfcd7e2f94f203835d56896a8bc716ba4e12e3d181c6d1ed6588b94ddd0f72f137b0c057a272da83ee60fdf397490d73326d7a9caa19d7d7d99c883d14f686aa6053bcdd519;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb81d9b6d2540c4aa2da94c058ce158bfc370f9a400d636269f9c7b55f7335ae88806f2160e609134c6db0b1dfcd0b4e542e90a9de5d6590159a4dbb4c1f6fb9f8a2e81d27b90ac516617cb8511a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117c98edde7057b400da3a1ba35aaea648816128b5e7732e3e6dc59fd4ba1578ac7ee323fb1d19649560c43b91f9e3b6d4817c15b56a7d6a1abf6ed90199e220ba79f562280fcb7d494ae51d6331a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131448c2288b0e0326a4ccd6012e545d8922ceed2c53ad601a0d873856df436510ac915ff6d51164172e72b291b4cce65d1ff8d138666ee1f8091d6227ed71ee9a9928fb728160a09b6e1d9e91905;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17cdf55553d4a8c95fcff90152858348793630f524276f18d35abb29bdc388714a6981d902a33184f9fbed9a4e2503a170f085aa11fec1f0a13cba8e67c48fab2cb29948b0561083aa949daba65d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cca0aa7d89e77c8a8d34c0fdbafb8f3b93a9901db8844fc359b11a9f7a65b8ec70a81e6f257dd901154aad8cfc836eccfdb14fc76103aabc2b4640d3a1edd108f821cbe9499a511ce7a775efa583;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1028cce25d5a8d85bd8775ed60d8be9760f7174ee210cf696ea78c41eec22c1d33f0efebbba6dd9f9eecd5373a6fd9deb5de782d70586374e4f68549b88f0243c28acbaceceab89d3c7bbd8df7617;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d97305ca23cdfb32ad5ddad48c84f5304373392515517103fa8ff6b682de3d44e39b378769bb325e755b7b378d79745edda250dad88f00231199789a17589db52f61509d41da35e794510080837;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d52709bf26f2014eab4b2e84342049a7e5e17aa009b20ac168123f883fd7b628fb11ede6bffb75cf259ea627b467c5e7bce6b3c44fcc344d9d156221950a157e40adc969f8cd9baaf050feb1913;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d14d8e8b50d994617736682a54e8c97cdca2895f933d7d587a6fa07f771e9436912bce5feed24173bcc99431a78a4649118662666a6810139704c84fd9651fd1ad4f4bf19c39723f41f0327bd96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6f3a3efc43c45f1073b15052d94bea538fac584d26645097db4b74bfba2b582544a347d57f54d944e687cf12015d8aeff02dadb48a2a75dc3d951b682e5a3301da44d87a70f325386d351f8801c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150961cdc3cdb8c1288c6406c91fd3b9cefdfd803f08f97f49522cbd94f42c77504ffcaf54ab4773a133bee373ee36edcb9fb7c704269f0ccb60fb7ef0bf6d5568d79880b3c797ddd4bd326073494;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hedbd974ab0df0109bb8f8aaa78f0edf6b7a17aaa9033cd5671daab9d4966df658554234a5fe8743c1fc38e0450a011c99789bd64c890bd4d72c29f11629f7ec6571a9951b9c5190a24d7ec12c198;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3e44a7de1db5ce99f11457f7ef69078ae615b1e68b67b65c1fdf230fd7601f4ca944565f69050b3bf381387a9276c5b72ac32a1969534373bb0faec52462c2508f1548cb156743f511025883b99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187f48c776e8b314e0c07d14b9e84805905b9afff6d88f9b0d5fcb6e1846f927e0f47122f99f4e71d5880a13d1b1cd4a24ebb4a86c1ee1b011068f4c01e522f1308c763948c9468748fe7425fad7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc15859ef4ec635b5f66362cbe27bd99fb0a1180f88d471675e1932f7fccc4d45149a76698c959edbb4a041e0488389457f3d8c3194daae33462b27efd5d087eafd6e0f14f577eee9f88b0869d6b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129043ec5322722ad00d9d3c61dfd8b4abcac237a6eec4859dca489362417fa2cb5fab96d6f2d35feaa1a63eff5f48dc6042f8ac4f59d0bdf1c85c5eaaa2ff7903bb477074ad7452fc0071d5f9555;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d74d88e0d2f81a48254d14a508f4904c89f5feb9ecb26f8744abb15e490d29fe3d4744b5c73290bc50ba1cecb6830aa345324fa8b001d991560cd118bb0cb15e6feaa52601b782993aac92fcffd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9afc0291b848f69028ceedf8d9b943311b8490a0ee62fc1f3c14c48d675003aa281656c93ff80485652b2475525fff2cfa6aab03cf3c4c0f697fb4fc3413b02a6f8fde805954b30abc3c3f59b319;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fafdd21d1913160c5a2aa3ed754c91618c6ad222bd780a8bd746be5aa1928e04a9b97541438c7508cada7d96a846ced475cc69863256a2bcb1ffb221b9c9a0c9aae602b07fc88292a5c1400c0a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27326942386bbcc0241ca54e74c549d249a835f0373fcc2d97db23ccda2433d6c8ad3cd4b60171dc26ec19eac34ddaa75f01232de153d3270253c7bca9809d2c4bc841e2f2e9bc90de0acfcf7d0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be8c2a6d5b58e643175651c66c173a03dd392c3ad847c9ca831b92df54f16782aaa9d4da5b7ea7aecaf2f9c1f5e283303809f3251c07b39f1e9de9c803e8d2d1389a5e7d5807872b98dfffe693ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fd5a85aedb9a55c33d698f72b87bfb87f966d70b0de8f1d2986035eab0bb895ce041936e723237d647cc996bc1699bfa2aa76abeecd48dd53d5cca504c5717f89bf2ef371f88a2b03df02e5cc31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bae287ede9755bb54af148a8b88078ff2c2ddf6b58d232d72855cce7364fb0363ae107cdc780bb8d553408964a45a4577fe1679622412fe526ec165bdafbb74ba320b264b91be2808fab9bee5d9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193c4551e05f46ad115ff69eae549cfa12512db7687c7b4d26e80560659bc19562c69d47f8826e94bbe1365c43df19cb51ee3653770869181b8b3690a645e84ae757e5ad3de407eff217870f19e05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0f2b3f85109b56253e9cb51d2d2ba3f8277c0735e140bbc8117b8b3af7ed4dc043951954fdc1c6e1e423f00f7b64baf476aeee6dd05ba710820a0bc2febeb67bdae197c5b7488a40a90362090e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e15ca87fef6e85a910c4e30dc6e5ad37d9e65c505e7d6a9efefc53005782824de1fb78426643de19b41769f9a8033f27da026753918a9c5452f49d529b23fcc8bed3077734cbd5bd97bc02259e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1815e91a3dfd184f205031bccf4baa0a2a365a81369e6244bb97a6a6c944d43de78f64bbd2cf2326bffb2702a2b11d0e0b6e6d602cb947283f73f8aac7820a954bebfd103ca0a87c5e60a99b6c62b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2349f76d7adbba66490c5895ad6f83211e30f98cbc7b5443338b9019b34ce918bcf900b86ca9c43e3bd04eb5c23f332d38b06447c54b1468e6d6e9ff6de204c0476115ef52e4c7ae650de7f45e34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1383f70a10a32aa26e5b47592790587b0e7b682641cec86d070a50b862ec25beba0242c60044fd68cec9a6e557188bdf90bea559ff4845592adfa3a4d2ac28e698a0f283cf0d3b2074648b1851648;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0964e2264441025619b66eb40ae81df8bfe7ea97511af3e14ed6e6213a090e52b5f42ae07f7884e781721c493276b953d635a28df1e65c7124821f075ca04ab2c786344da25056a42097923bff0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d752372e0059fc45862fed46baee5d5ce9b2efc26929fe01903160dcf1f8f966e2aa74bf0f37b6d4f62d23ed685c774e32fe53f16bb059c5b53f431e9cde5276106496a1d44b5848606b348a69db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80b36bdf68c6a0c8b5f2f1245dbecc6145bfe8de4624689b98f7f77db7ae4940ad0ee4fbfd54204a81ae11cb18d70a79685040a5be745e56e1eaa14a42e9b1df943f9abcd5b6d3b9eb59fc6f9982;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha67ccaa295263d7c5e2e83c72a32c75e0ad1bf3829be73f5bc15ad09fec222695cd1dc621fdee6777e8e469a7983ece493459f3c699d596b603e078a29370d90c93beb47288e5fd120a49cb9a484;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h298ad577bfa3e07371fe624ccc6fd790131c151003c0c288e73dc720add6ed9e5c596ce3f477ec3f67a9d2f02845a6370d0df1dbf72a51413b46a28e49fd4680bdd347e43bcecfe6218ea35f3436;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb99ca63ee869a0a9476d390df7c62783a89e42c3f58eed7c15c87d7303e3b767fe50cf82d571c32ac58d547365f99f70712ccd077f291e9115945cc72bfd966ba477172e0f2648a4d01d141c626;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182e530e331bd8d8626c45eeb9096066f10f31cc897a2b07f20d6aabd3372297b5748d8bc8d9a78dfa562ff74084c25bfb120d2bcbe1e2e25ba82d15edcec1a54a2c4c147c40b56452e3cdf9edb99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f823c0a212acfd41aad0b95b08054ce763859ae16178015684b91eafdc600e5b3bffe97f15d87642c19237f941fcbdbf2710973e2ccde7c15f03be871befc8b010b6d5a4af33f8806edeb76a3a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92912fa50e63832b06c1c2f320c0ec742cbaf31b00585cc5bbf87b5cc3a15954454bfba17ffc2a1211dfe4ff24a8b7dade50f8a38dae08d8ea64360a66a6f2351678b9f43c352df8993790d7ed7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186e552a680c0d85cae5d31dbf1c087c87325ff4e17a0ceeafe38f4efbf39487684480a11e238dabb804230c620f3eb5eac7c9aabfc73a98d15c0f720a1656a03b6a50620af8c0b1317a8650961a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a8f711d26d441c6b52da69273a18f54efe63714c88ff744739a86f64eb71ce32e95a684109641288b475be3975adeb0e48184bef273179dd1d9da9dabdf06686d5bd499976a9dfc48b3a0dd4820;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1819242441166cbe13772e74c2bad6c4db685c479047bae9e44911afd27e71eb3ce80b6505717bba4ad7e6e060236169921401e2e586865882dec18bf03b91ac3a75f81fede89c81282f9906c3675;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h420ef881de0f12a9e6684aeaeb304c095ecf9e220cc06a9bf949ec029dd976542b68aa73b8a6541493f066a34003a7611f43d93b8ba83a08ecced74107610ed260d8fafe146e3bcf4ac1e1b4997;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae491fb6f79973b3bc00143f68c3edf8e8927f1c4f60faffbadfd0eff15cb580c50dad8562777c4556e28867756ad11ca3b87ba48f9284a584926a033bf7db020880dcdcf6fb4b4a45a01cb016d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heae99f366a16f8b9e79d433546cd407bfcdbefae53a3518ea7860800156a548dfbb5d5f358cf16d46bc478349e9a59dccee078afc2f684f64aae4636ee8d78a13f191040da47828bad714fde6d6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h809c1446d9865828d7ba16012ad60a3d5645ce0653068aba687fc73bed65c5048556c26a34327f8863965e244a7d56f4f11b6407e35f1732ffd1ab5db7c2e2496a0876c684755959d92bbd50b62e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9da0581d0ab1ff78e24d90ac520f5a5718a8c56f8e09c0ac17ed2c8317a14828fc2be806f0f63dd2b6fe8e210f6c81b2eda82f355e85db21ab478e71f363f3831aee170461aa4d3b32cf776d218;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habbe7c44aeca7cb4c78edfb0af77292f88c238bc28cc36177fd429f428976fb92b3a6a55304a139019fcdbc7aee75c762dcba6dcaea4301c5eb5e5ee42881c040c3a673c91cc62948ef668676bd9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfac69781a27a34f49c2c7f53fe1fb0464b48727b4d6fa9b1b2e3bbef0db070f50f18376dfaaef4ec982336bd915e4d7d96477867408e9b8e3a099f76dd6d88961bcde566c84f47207fcca6ec38c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c879ce1fb9ee85091a21eb4ab6a1ffb5de158a4200357557e93538c64bb8afe1686a528fe7da6ddfb98fde69a5a8877730f027c73fae7416c367e6328b53cae2ec165060674ee5598cc92dba4f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a6ddb95e61003f2b60d4372cb7cce67436b2e09b7f94dc0db1dfc3c1dd063bca6f861fca5173e4c9ef6a8f3805bec19ce746ffad93b9986f2b2f7be0f144d3ce141289f0bd01adabd9ed9f8032d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17320bb6c9e07ccd2b7e376725fd5fe63b23b7a571513873317d2d57658b1ad4d7cff170e1c67c3010b859efb8fa21c606304615ea4b39e0131dc1274283823f7204fdffcd1b9869213a74cd81961;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18de24624a0638a124a646c15f155cac263a3e59636c80ec93c3fe37dbf6147540601b16d9326730119551aa4a4d80e29e26de3f8493549d2e3c65d803c72a7f6c9938d4fc0107f7106642c3b0583;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32c7fa6eb174be5e554073fa8a79ef2ca92252f4cbdb4c84abd002c534cb7c007c94ac6f9d014c8731038124152ae4375409886093caa117d06ccfc2a0e8f0f334f8817a2e3ff8462f6b06a3f7b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162cb4526f74553fff04d72af03cb0506472a25e15cc8aaaa7410a91bde7f8ccefaac13d3d6d7b533b8a3c4749e21e0b785a1e3834f286c724b1052bbcae2f627677b92e84549bcaecbe9d502fed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c752a811696b0458cc9cb20aa06463f1717057f29b7644eb17b5c6c2c43381714699a63fabac50b2a6003fe6c5d0e572a0017d102d61829c6b0d2de1d718e7f381e0cf07d8347be7c1a06f16bfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68735e14d96abd30c5b24688e2067fc13344a9254f43a7bedc6ac1840086680eb5b1b4846c683988371495cae99fb75eef4248a15276a98f63139fb936d9c942bfb3ab3d3db0b59a0f78a7630484;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120e429f0d7a776ce3734ccfd3218aeee9a5031f12304f0e6474b23126a1d9c65e39c7156ab63dc520444be668e9883df32ebcd6336790d38fa1bc3453e921211c5a53efbb34e7d8f4439dcc71713;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bf1a58502aece138d9bb68f3bc21723c19d1b5a203631588e1785e607784fee32f6ce72cfd3b31ab5bff3ea11555e885cbec032439586901a4ebd35a25744b0a67d183bb1ad43d081e366112e67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18edefe07b7c5d297b9fdff76f8e4f005e9756afb26cf9aed262b8975ff2956a196eb47102435f1ade386a4c2d71792c46dc94cc62e2b520964784b98059eef51ec5675dc02d29574aa264ec5717f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heca08826342b002a34dfd9a857b7c333e1503b142523aceddfc34eb43a3e7b902f53dabf8ef94dfb22916312abcfe30b0a817096c30e138b1e15beb0e4277d99addf57355f7c6565093ba78cea78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e542b3b98219c4eccb0a0aff203713a3a924b3f099533fb9d8c339269abea9eae9d33554d247aca5fa10afae6afc2a27aa2c21158e6c392869b3d1ea184ca9793f9173bb373ee0246f1d0c0c59b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4df270e8d73ac054c661d7e2dbaf2703e0b89462dad62bd339b4f7fd59b37de8dab6c378ba9398b93a677f23cb37b3f6bd42fdfcfbad1c18c3de32e9ce05287a570789143d9dfd2192eff96e218;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he40cc2473d71f89f4bff17ecca1bac8a1b9f357ed735a1243b2578b3af424a4bdd53016662751dbc6e3f33f32030c51746c4dc0996f4e0d497fe1507082d0bb9ba18e68b90bff7d7ff9b442b91df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6faa147445f073ee90b9888ac34471e41dfa34b00b4354e46287370164a85de11ddc6c4e6a355a510dcde14a478a419a55508e3e0990febef7f103623f538ed01e2ddeed894efa8c2b5e6e4053e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h313130be349d283918056725f7bfb7effee11b1621838afa72bdffe36044780c8c82d973b61cbd2ae7fb22354e261f12d3ac77972f88ecf62fbfb7b90fc3458f772c1b461073bd1776a7c3abe8da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27ea72fce1daa718889e453f3928048fb9bf04d93376d44235575bfb2dc43e5b6fbec80b3b616b542e339de67d8bedf486c0162447f749278b71d1feac77472f7b750c68c046153e6d58580069de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b55ed1d1be1edb662b40e99e37a398c04b415632fd109eb6533aabb9d9bcc1db121a555bac513e4aa871fccd3b4195bc7866337d956260e1720b0331f79f6cbfbb5ba99efab0db23b15ae667391;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffceca8491987aae00806a306124427acf5ab451493b1de5fd28134d55127f60fad06f460a5ebf64cb5a4cb939e6c7097cb551074174f712dbae2913c8cf4aebc8be966933bdd64cd7a98b0cba4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h380a96b0647c22295bac57e8e225147cb36ce5908c33213dcc6ba6476ab886ddfdd5b00376b1aa2031ae75da4136833abf095494e352cdb0cc1699587afa676ac5bc5399dfb4f788d886624c30a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31df3dad9dc2cf7444802a1f5e44470d76c5f1880be87d6fd36bcd32c1b6b823f3098f7e9bf673758602c335ae0eab3c4b3f169e858523008441df8677ac69cd86dcf6a84c0a6ad5adb1f717ac4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he89eff08d96ecd9cc39849a19705083e94584c8f46da403e5443a3c31e53e236c0dffd5b14750eab47e589de08593bd48ab2c8d8ec6d3af6adefb8ce0874a2d225cd593cc1cfe6352d2f66144c38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1231fa492831fac065e4d67943daf663e2bec39f818bdc6c5b26a12c7f1c7fc2ac35fedbbbe9c43678d6c208d4c67eef4f13c52435a93e11bc3f98216162c7fbd6b7af715e3a2ab70fdd22d1bba66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90e173670ef4b1995c388cd95be484d6326b06e3fd7a9ee7835676ff94dff6746e0deaab819ecf57eed1e0f949bd290bc5b66bd1999a6cb11101d7c699091fc8b9ad479073eb13830a97353e8b98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75a58055cc204d9772f06daa8e96ae6ffe6f578aef6bbbea6acc61129295624d54d0866e56df459c65c5197413d57f7077c64299a85a35a0d33bf41888d12009e3cbdd5469d628496e80ca74d6b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8100227969796966213ba8c3fded1c27d7dd1fa9742c32086ec65bd78ad4b688953c18e298950e76d6fb86609fad6f801ce8f0929c50005bb51291167d46c8e635b22945765622c2a4805de495ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4897fb1c547c910aeb5abf37115aa9b80717d2833178433ad6548e5acce8fa93fd738db9c77da90501ec7c22f9b8ffdff9c50fe228b3ca7d35dd2b72b7ce24eb7e0286823cdebacf25afa8b11eeb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16056e2721b9f6c20bd7ef66d8cf482acae78bf2e18ac992436d8b341afc4484255962838b963d304b267ecbff866071b2d10ffc7dc137f9f4df7d8d26f8c88f4a4fae469b94d3c231a5a107588ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78525eb9a51c965343b8189a0b314b685dc062c70660e428d0516ace57e798ed2adb189c5d3f7fa21f9908175be80fa47ba2739987d4242b897c46c29e1b5d5787cb0beb8c7c652d73d0fd2685d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16dd06cddc6342cf29032f4e6b30f62031e32b0cd3d1e1787fe73f33a4ae0babca7f0a86c19a61b3a10fe040a07c574802e888c4ebcbb38e4d9875a72be60a9a73691ab81ec91ccc7928cf7c3dbf7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h396422967f0a0e9b3c04acb8336fa8720474b5aa422e66479e107a13985b7bc9b227e9ada2613a48668682f0e8e4a85c51e0c0e8580a231a37a9527fb6a8667b4bee78ee8bf3247f0159792c5d75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h790e4470f649f653cb623ed3a3f57a4f747492dc6931ebd7d4100d36a13b71e51beb489644a1fbb6d4bada8db0f1cca3166149e2812d5baf4b1002124cef573a5518d3b42063fb78c41fedfffb12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6808d5f7f89f48ad6b57a7dd18f52712b57d39458cd91f9b2d84a6a476e181b80e55c157208f1df6bfaa9e708b6d4cae8af703950f04f1b5c1f7f879b14d99e955a33b5b9ee6ce2914dea3d33fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4240995f0d3adc9b6c4627f42964bc88f4c0219e8bc926824064285ac7e24c265032f17fb63179d1ed307d590cec9d202c12e49b3892427b26329f4259e5e0bedf2e3f49865e7836fdbaa213d6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7c29ebb9d1a793cd2aebec0e4ee00928a24e35b9c27a30f922315a3216c2982b17508845f77af3fd86ee0d9f8d5872d10aba37d065520304c8090b9e259062e209f61b4e5b20e6f26fa95b94e5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1018b9ebf4dbd89c0920c8d17d796f0908ec10e6c4d43c3185891e0248b2057a7632c065b37fa00e319155d1da61fcecfa3d32630a295fb1669306214861460ef25d1d441a0dcc96a179fe27a7a14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1220bc53dc4e1f0673b68495a23c459249eb9e78e2cf5be4648d294f886bb6c48500940aa932a58a4a410188f396d047bf78bb0650e23f7ecff1f7a78a923fa02c58023764db03f87085f32ff60a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f91c4827d9d6a77bc24384fdbc78775448997efdec0bbf81c9ea071b51d98fdd5201d8e8f73fcc65d4df3bd4f8a37d0da40279070d3ca4bd4af161443d50c3b221d7683c5d5070dcda95688f855;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c97d6a48647782bfb3230c8967d50d5efe9922d0b34071c4be5f34f9e4467d34a0eaa6a19b97a60020bb8a2b7d3f0f41c59bfb2fab2b1b853be33373f17e43bdafff5bc6945e1a545de72754aea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac21aea74bc2e4b4958bba112fc1af2e644d81bff3972ccaec369163e8f975656f1295fbaec2540c923fd54939e749e7000b721f594e4cbb00e1c166244987d9202c8a3e5b0bd70c56ac46221003;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a8ceae376d8bfd1d93e35c1aad87f229f2f0b0f7efb12df9c9557d77d43c29be1c56654203d815da1ee9aef9a7c57f78b22de678dc6f9b792a8687989c491ec20834a6374b8d37ef6acc923dd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d43eee92a32f01143e0b602c435bd7dcd6be606063c798d7f51e6313203462a38469bd6bb02af188ce72014e333e77821917b54382f66ebe9182f8dc2aeec2586f1694efcfcadb86d5d6736aefc3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc198e85ea0e0545218d62e34262b4ed1defd7b20844be7fd8b16b4d7a2cd2e3a4446e244f57dced8069a15486bfed38fd5d17813f8834c64fad21de8b1baf9bc65907bc1de17481ee3b96fc139c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdb7a871e8616e868309ef8997255f52b42aca6d89c6d608526bb6fc40d988e3b8cd050860b8d3603ccb8fcc881b2215dbadcd3f300f4fc8e9be44645aac55e3cdb42bca28a4fd65c6dc892df208;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93fc90ae09235ab8005a93fe4a9f43d363c3dccf8bfb5f5626a307c31d9b8cd1444fc9f9251cbff916895deb718f925c057ebd820ba2300330cfda4bf8198fae8c6412a0f12b2175fd75b286eb4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5f2fd38eb5fbbe4a7869e2f67d85efc64cafbd4a7729fd0b4f088cc0344877b06f40d59b2b45788acce527ececbeaa7b812279638584b9b5095e00ec4dfc7425649c8045855b8df092077893ea5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65376fd037315b814024c8aa076b08b81f28a954a05ebdd47537c5be3195cac7a48e2d245c5319fc92c810e6283cea6217bd9bff9656825ebd05511cdf3d5a45a40387f95aa5a7e191b98abf1097;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153ffc2a83366cc7ea47478b18713ed7b0c5891a6bae8e88fb8f9257686358a2e7269fe6f2ccf23fa8106a0e2bd12d846d95d7b03961b5f2d870de02b7d1f5d3ce82a77c4f04232bfb6bc59d2cbc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2a8afdad24b485d8f7cff29bac8526f35e7ca586cdc29692fad846401e288272fe6eb9b4fdaec0c3e2a29b651cef225e74c8f08ace6bd1d26488bb9efd5df0481b4d677d5de0202f90f592e9e6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde1c650dd28b8c63a670dc89e0671a952ceb09dac4d6a4ffd2f6df374be9fe6926b832f8949c4aecdbd25fc3c5ac6d4dc24ccc418c04b37bb6b528e84747232f49138eda8446cb99d4ed07163048;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e96ade66970c0e01e3936cf0dfdb6e3619502d01e9386a92bea0b82ac951d7ff627b62ea23f8e457de019fef820b2021ae34906ea5f7b80141f787673e4db8fa6fa844f3a4016916739891cb1c0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb6f184c73f814bf86375411dc9ecb5689daf4c8468244021b6084316ed852e07a9f405dcd41ed6ecf0c78767523a9cf2f2073794ac6f43a2099b0bb6245145ecbaa029163459cf723180b26410f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f9dfe4bd1d5792e065ae717ee130e04ea4f069fb8865d02a6695aaf2b2c4207c095387a97cf39183dc98116c076a011d9eb73c8c4ca7712f0e0c7bdfe76d18fcbc08aa1c81cb4fedb3d450307e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ebdc30ec64f18da1af183c82ffd6feb80e1fd4f75ecd49df49c4db6a9dafccf48b72519054c924b1be01abaadeb32377a777bfa5ce02281764263eb880a1d0bc9fbb16f0d102fcca0876ac081db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52e58b1d7da66034c09a0caf2d8944e82d7611bf54955ebcd52cbf58bb23456bd73d268f088b5d65420dd02d0a2788b6c8e12cace28313917a860f5c3c9c791d318021e2bc3f08346376401c6c1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6215d9fe199ca76e525465c6afaa2fba11b5c42852ccae7072874dd04b3d3111761dd57990e9fd5cea6b9629ca879e4e61c0f1769fb1410b0b7258135cbf233fe5710290972bb2deb7abccf6b727;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132afca033998ced4c4bfbe22e880afb9731fbc99852535f1b392cd8c63ef0d1568669cbf8ac853777636426d23a399e010534ad367055a267a25a9533c81ce7ab57babf0ba06ddefe0eed622be37;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61fd3004c590acb409b7ed2fc1b7313c13c94a67f4f4613718c2117277702c75afe9554d7ec7b6148d2cd9cf7f3e5f3d3a376f7fd76b7445880f77e77de8ee66f038765b0aad12142157119626b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1452e622a0ca332afaf21ef36c8a41685cee49d9ed6bfe0d873659afbcf966b77ce56eec1c63fb0236bb67e7e52671f2754d492e59097612983d3f2ba562b05ee15764d2e7867370864bfdd69c793;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167edb10e4fd26f581603ae5f605880c1c896c3bd5c12ab4ccad5d6a53585648491c2974e45196a964ccb706ec00628c358962e9a91d6bd9a1e48305658fc458f00f97ee609f751e1a6bbd7de32db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102dcc873ce7790e4c04f372455f27a3b918eabe70b2cacbf6a23776b057e9fde10d370bd421807be3afb9729bfeed3064afdb03ed23d63f3bcf5941e1b9db770e9eece89b084fb5b76e859c0713a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12098589dca335f8a46c192a26bb6dc5ce6cc29f27501a45557ffbe1a3aed6e93d1ee9957b46c1627d663b9b2145414506a1e005fd3dbf31e64c760fc28a25b85855c3d4fb3abc8503f6c794f26a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ec4159f35d69dca5ec4b2ed7889b958f2a9e4bdeaa29d717a5b650150fdbb68ee43e755153e715c075dbb60dfa2aed10b3e816ebc82b5ce243437e86b4a839850801a32e7b83b6f7bc2ac5503e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1511b437542bd3154f3c813bd408115393b0af10daa86c6ff3795affab120bb8ce5f683ab8fa28510da69c83f2a1423ceb2fdd5fa11025324c9fe8dd3b9ebc8dc3586c1890e0d769b686818892a6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18700436e3f02871e812390299b2ab55e73149d0a1f352a27df49e55695260ed36d4bebe57181029ec5c31c79983b61a2d8b93a07fcd6d174eedd46d49c71c2ccb3423a6f722427042a3b53290f47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92a5f0ff72fe558e5860e49b43397cc2bb7c68b9afec3423d62b96052ccad8cdbebdf5db83e0f0ce52426a668ce4340611bc7067999ac1ad407b41287f834613b2c1462f4de8ade72db5e29f0230;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h322a546792b07388e6613c9a79ec597fd5f698abb13410b797be7c66c382eb50b9618c1f143ba7363a67ddb9a907add13edb09fe9c8525962755210e52008e8706dac47d00c32b5dfc2df9ae3a13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa7ebafb016d19cb67e0cbf0139a6be8592a926950d8b86e27b74f720848dea8b9681ae6ab6092b97c53428ebdda2e72e68b4bdbf833dfd594857e1dfa1c7cf4cca976d1824e674fd081b78bfe91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c63c44efbf5ff3488a2f90aa731d8c12220adda6a937283fccef374ca9667480f3828a4b7524388201d96c0edaa00ab665beb9241e5d4883cbc3ba9e5a3417152dbd4c2feb8449d016cc974106d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b819c05bca58d32fa25b1ca523c302d5468dc269c128e41b4cdc1d5a1c8383f17f574dbd28d26482fe0318821a6fdab89290a985a2c7db9daba2c5a3b2b8c2bc543a11a4a3bb385d9ac1f209e07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3889c5231091fa0c974ff94ef4edb23ef5e34cc3783c66180e1eba1eb5818bbf6ce8d5d0aad773277baf0e2feabc3e33e5f8718d69dceca8468d8e092730a46e5c839dcae4c13076e684275b38c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1812b20a97462f2a1d2de928e15e16b0a0abecc1b053b9430a96ae657447f928d1c4344ed74413979c123944e8b8609cf19f3e9c8ab5f18399fa6dd106df69c93d0513b26d46830233d5fb1bb9061;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a43c688fb3fcba44da0d7c43ff3a2eb96ae0dc5623217d5cc76f27a833b3ecbebb3c36fef5921888d351cc5d70dd1a9a409abb36a49b89ecb2a431204730296ea1041bbf22558a52ef179208b07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he57eaaa8bdb503b596dd82143488a5d84462c5587cd7569f9acb3abeb918d1b801f018593e7eb2b520c22d560525727871c50d585731deaaafad2ebd1fac36ccc6a4aea47c0f7e6e51d4c492356d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db51fa8cb34a982e2c4dc968b9b6814dbc6484b0d09b87dcbcdc2448210562d8feeff3423ea2bbfd1280534af8c51ac84ae00cb197b5408e2e9758750ef26394dfba04d8cd28f2b673b98e16496b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed3e7c18d1fd33c08a75387741d320da450c0bf55a0d04f0df7e2d471e97f698b8cebca471f4569f47dd885f5ae09f91c04bdfcd352b416315506486664946197782bb61c5b0d3b767fad34889a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda98d6b44247eb3a30477acee4d19c52070e72bd7fb78fe31c150cac8c5b3b3e9cbb628d7ad287e0cabd4feaedb2353b408d2cb0cab32e0c9a2027fad8197bc2f37a04952188e3a24403809b0bb9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c800aae2326a670f13229502f10c944a61ea2c1c01e14c11e004deadc95219fb6e0fc7d805a87258fafc266924cbd448d47509081c3de1b34dba15540639ea2620c983650ec8b1b4475e3627382;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98f2b1232c955bb41c44092a66e939a0b50ae17caaf993aa7fae4ba2fee831a6d3465c1b25fe94307dbda0e846fab6ddcd22adc94f8429705d28b2c7e799a351c986a52e0a443d34efe4c8d0c6e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d67c0765678c1c0e8824168874e80267a75636c8c8803ed3298277967485a69b70e66427a5073f685b384f19d08fdb2b658025bc9859274e0e8b2539e2999e6c5d4e7b8591720800f41ee563ef6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189d5680049048c2cec777b141aa0da3fe2d2396cde8d96baba3a272d11aecee6c817260b5dc16dd778874fd68a297b3d82b70705ff0483f98df658b097fe47a3952abbd20e5601093014ccb62fa7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd8b331041acfd2190d1109b4e8e7c5b1e1b47e50aad6606b0b0a2c74dd44247f0f60c895f10f0ad0d0d185676fa190501fc47148e013ca36a0b6dc911785d11a264bee11f73df43539cfabc7836;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9cbf94a60357770c6525819a927c9375dff433cfdceb97159a4e871d6f137747071eafba732aa612d3c6d986fab07caf773de1a6fb862da54244f6735e9275b9fa5def52e594949f7e5dc6e9a3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145ae4a9cbce3c3679bb73f9bd8ec2b12185405e311b761920f4464a2241d93a7dc0435664b7a0cc62c30c0c7b375dbba94d3a2ca75b226846dbc2b0a75ff1c1a12ae08888f752ca20388d0a9f621;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10454a1a3d4a6186382d79d2d3147c45e598366588d99bffee2eb764bc388bacf1c87b1878f318d2a957fc5895db84fe79d529405a1ee38dbc734458f6ae2791773110a7d591c2a518ab29078500;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7aa7f11db463b7951f2691a40c642f448416d60b03fc1d237db915f0178356958f4fa0463bf7f7370e9cefaf667e60277b0b8ac71b46ccd2c24b0fab18b694265530d1530a22fea81ebe553568ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6613460340268c8c0dd0c76e762094661387a42f48f099d556b5403ca163a6f47e7105dff942892f0d796fa2d478b741dbc1743969cadf69459d2c757f8080d744d95f21c16f5ff5a5144692531f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1676a17597e508fbaab96fb6d3a0ef724b392adae11b3b6180dcd1a4b6dadeebd806f697403be1849acf6c214d4df373714d3941684d103dc609bf3172768ccbccdfe7aaa1ca5ee1a8a3eb20035cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145a5a5929f7b8977196d2674adc84fe159665831ed87395d8c67a9bf006fd5afa799be44a99f55f768d18405da9cb77895e09df9802d16cd6b4d832b7375469b349c4559326a58a9315a53735caa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h767b69023e359eef0f660685c256e5876493d87fb798a46cd3a76e901a49c8e1854e14e2d830640c5c3fb7698f6e31f50a3ea61ca28ba19df71c48d797d36dd8ea3f4e17e0fa745ecc2d2d36abd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6df6ffb406b727a80b942fc490535ecfad3a9508daf04c6ec193a18cf778a7d65a0ea775a57bddb0f9e5844b4b905680dce6b3fa165adf666997481cfea9626309de2a6cb6b07b314262d7e189f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1b2fe6138adfdb47205a18edafe69931357ce0205d6bafbbbe75f913d9a9428f02b6389654c2ca1288936ef4640d3b2afe320094915f61677fc3b967395bf784634d6b587c107ed784770236ccc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0b967ae25c630d13a119e8c44c33aacaf915342ca53a18b815fdd3c41996e51dee9287d66b42e187ba61839bee74c55bc635c12c6ce15126c334a4db1cbb6cf448d42ddcd13039d6b6e1cecf24b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66ddea66f87399d92d0cefffa8800aeb72e12275fb103326079f782e893e0abc58f215bf52fe42461ba630e41c608e204d93227fcbfcc72d92fea87d146af72dad754fe622470ab8d0fc8195488;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118f2b705a1e67114d557d66daef1fd969ef2fb1995b9f2e7c47c4bc831c556c5a1531dacf9d656501f8030c1b5395ed086b25a5a8677c78dbe89109f5118fca64a517bb6cb96f67dac6ab18b3748;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c35837e35eea8fc4061eca67a4c5305401d3a50b04247da98cb1b9aa17a078e5955f6bb403d57811c161f66a23e4bc7574e075b3ebb5cd91a61877eefb9592f72e55ded3488913356f2def1dc3e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17aeaa97caccd468ee21ffdbc18ab1370007a2689373e3ce3bacae6676ab389dca069531af90fc60adf265dc1a9b2f6f769fd9e3231804ec18781be39df07a8ae5b1c9ae29f4a1d3ee1e17d84b151;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h586b484d9c0e799a56e30a46f932231ec3bf2dab643a40f6b777c3051061882f989e4e9ac6aa4a806f989544b7be7389f5a93ddf3417aaccc679ce34fcd743ff416bf42bd2dab7177dd0b0708181;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h73d591b0f73242bdfabb5da8133b673b60d1ba4d741025c8a8cbf1826db6a1bab5f57b0c86fce55925c942197e700b21fa5fc23a9b34fc890f223c4cdc45e1f79cf46252958492dabf22a5dbd08b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87eb471dc86069c1d27b9f83723db5d544160dea07e29d5148bc25c1bdfaedf99b41b7da31a5d38fe74a089ec9460a2cd1032a4f3d076858f935a1ce87bcfe33b9a6722130eb8714f510c5ba930a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3e05c3516bf459a628646132a07221098f0f4229a85bc3523845e028fc144bd8a749dd1a5e0699d0d54fdd675fd7a8282d88373e9bc2d923ebba85b3a519905867820efbf369787987c127b2e69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f2df71938dcc9c20cbba8dc942e639492735f76494e6280ffea8483b375f2e13c6865ca46b9d3b38a6486e9342124c7f30500cf036ef38f144373352a087a290648566a24792dbf83736475f8c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f78b1dc5e3142bb58b7e2216e3604ff93e8e2aeb851428c09b32c4b87afb4677e8c7f992a2db893d3882eb44c054e000a97afc52eb0641cef9086f7f3e0e6b8e799def70002e338182c5c5a4e06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b4615edf1586da5a68a3e8db4fe525f22942c1f8053184e0d7db8b2eeb1447b48e8bce2c3a6e498821bff1e3c51ab1ee6b4625a2d616b177f9f9f69c183bde71c419337fce74769ef711781eb26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1125a2f542e6ec06875a6bdfae633a2a11970cb6d576ac3262289c32c53c9ea26c675e95f3406fe29f9c16d56ebab301b04517894f63985a242aea34fabe8231371b216710e9a338ffb2835ff50b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6f3a1669b8bcf31c4bc236f799b413ef1755bc67b1ff71868487ddd262ca3ccfd3b1de7009f405db79e44fa34bc55027baef907395a32a083a762318422f6837f309b232ca82a790b25b89ee5e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8a11414066f2b44637cd95ac32755e71c6c51177e2721d2d0d525b5ecfb2dfcceed81e6c2b74b45aeacbd442a7d96e65592be9751708a50e4f322a9aa2bb7b2d25814590b7c886eb2c0fc4c81c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11dcb8568cc8ca5d8d696294ffc5babb62ddc2c9cf7a8a22dd936805b3ca3f220081542f20585af10202eb4d9be61f725bdd9d18681726d9d59efbfcbb79bf03d121adddf78e2ad9cab6bb4bd32f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e0a7c2fbdf12c134eb5d623162d6ac6634fa6d64fb22c849da9b6ac93f954c7314b9b24ceb52d2fd584645206b6a5ec775e69eafcbb8ecf717f880053193d0f8b1f116e589e67338f1e686e6aed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h497079c9fcd017892637d332c907b3387c5636f780a512166d22d52fd0e3df3254061193b271f137c921eb4d858bd1183ee6d03357836bed9a60366280a520b3b631c46782df9ecc41607d9c6653;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h366050fca5f56ec9cb738469e4d9a5954a05c9727d9b096d0db97ef65ca4b9f31fb7ed281479b838d5550b68be8106a96bef555ed764c20b78fa22db25909143496b31b773ce6e57945d5a63befb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc17321e7df56242cbd1486844193c422f5aa5a078f100d1418b4ef24065df062858b29671c465ee116b846d30027a7f38c3599d40afac1d531661164362436fe38b36212ed1585dcf3dd3c0cf595;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123241d1b5cc7409e650b670aa696c26f8ddfe21950eda1f802f37b83fd232580e9b6bf9fd45a534f535c0692cda193a4af88e90cead55df1c5b2bce891f2a5145714e007378a1e8705d9b673fe4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb352f1e81b176fcc966337a18b5b755c82ba854dd1222620da03054a22a3c236d3de8c0914eb4b4c13e019332212ab2e419cc9aea7ed2802f204e5874486c472da65fbfb448cb7719dfdd5c01ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0776a24e7843b1009ea514b7104d749aef1055feceffb1763d7691d001a451fc13d2dc9be374ec203d6caa7a55a653b3e419560ef8068eae24081a9f3121a16d047a051eaee78df1ccb0c4148;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78a9acc8ef60636e4cb2c04672d2fcbe12fc90fd8e88c9edf6c556da26f5a36215225089bb6d73021d4c5a3225732c4c80c36a20cf0efd2b49c292129efd24ddc7dd53ec401911223be189c970c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131ae0ee883b42e891fd8db2fc5a223f459be99ab2d282e2edb8efd2fbf13b1fcd42bc1953de77913064350775199df1d1b3930b00fe961bc1afc846711abbcdb7d921f7a306b65894b3262d494a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfad759e0d3f552b9218a51e101389c8abeb6bb6307c0fd597eb4a77b2f70e94cb7c3dcf242593108cddfc303b76aaede017a3ea74f6392b75ef70eb327df1e2496ab53e6053293dea8226c30fb3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e790ea706bcdebe3172877c3a9a196e6fa60ed22b021b486adee3b07bc1f47fe470d18ec704d21e42e4dd7930b1e7e31f39eef8397e8590a0001a5e17684a1306ab6a4c22db35e9821588a7306b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd218b9fcbe19477cdd79eecf52659a68862e30bd89020fcff148588405a82a8099f52e92dcf17e18cec50580bb96f03298a994b4584742774a02b2f9d055019c245a871b9ad0d17df6096a2919f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18db8f74814ddb59e9cedb9e2c839f8473b4eb9792852eefd50ea1dcb251c7fd886fb30f1c192342724eabe4a6ae3938d81ddf7ce5836750f01a897b47c52ebb20635a3160744720255516bb36661;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf13038c451942dacb242774311e8b9fb5f98050725dd286d28f83027b58875586a308397fc12c708574ea172cf6a9fa43d83e01d7b15998de5be62e3dae252e857057e67f9ce4daddd7c189097a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb882f403b17b7ea04484de921b3a657a4b1d9280049d2d7289588c60ebb885c1e01536420053019fd5e470b2c0a159dd9794aa50ec13b5e1ae2031f2e5be529c8f46c2643166c76bfc950825dda9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58c0a757898ddf177464c5d949e7488858c1036a0b4e5448d92519ff14c12a37d7b2d869d0512f68ccf94552b7330cea2df2627cef3c2793086aaba6b4e8b2adc64d73ed56617efde476855e33cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0bad3ab770f835184db067b03026672bca8781e0224b0272ffcd587c08bb0df70b2115b573c9f04bef5c2eca45f97c46570e67e8d32f16894e01b3c36d33873faefdc8588f511bcc19408192cde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a88963d02e49e56878ff5b581ea61bdcc6ede15c421ed32b933745ecf6eb31aaac0d39770743f7f2f6f6fd3a6bf18ad41722e7161019e80dcae8ff07c25c111c14bb819817a254574f846fc4eca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d1c66fba67ebead9fd619457b07e75b4936085f5fd71c764ee17e51655067c5ebc7d4d5d589718dfda7b7bf941ad337ea8b65eb4159e839a05fe923362ef31042a1472905efd28c007f6db5f25d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128dc1f847b204c0faefbeee292394d7e3c6b232e32fa210d90d4f8932b3095085e0673d14f22a163040bfc88d272f65f387bb4d892a83abda08c5a862f201ec61297d6abb915f624c4651293420a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h428501fc5b3649d01f05233071e75b67ce5aee3bafbd8b2cef38b1b475ee16d61556b8d52cebb327817b6f9eb3e0eb6ac36abc010441cd02f293a3d7d5f5dffe82a69f429c7fab43ba3ecca00ee0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3c526652baa4536cd4971ef14556e0cfdbdda15ec64a3a7d382f6a528015a92eb2e7a7ad4ee67286e7350156604189dd373832b3ffbc266088e807c42bb51b7f56b3ca6b49083d63bb8c29f831b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5e82b48e526ec33be1d104c12594bc47afaa4faeac0f651378e4643f1f47523e07a13df660acbf3488c29b13a5067cc88345c176e16d0dff82dbc5c8ac70498876e20bade4874977a4ff732290e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58f95e1fcc7bf7e20dc837493467e1f32b5efd181681eb13211515a0bab7c5ed430167d463b6ee0d6a0a749e551f50a786a96fd3537c1004b9f9703cecf70c11f89c7a9de18f64a7b4c234a07199;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9193feeaa7a918d433ee76c1826354324a57a27ecd5fc48e18410049993f091366971ce35175c738d8b21cc7a99a1cbfbc7eb9a91db68927f53b6642410b5c98eefa1315c18deb2991c5db23aca6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e686aa08387807d0beb026dc12e204c671fe191c439515616ffc3aed7620a7cc1f0c1700468f2fefb6245ec5f7ef09c6c4a967fb5cac45c20534468ff5d2976bc1a25ebb42ee309344e0cd7945b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed8c1595ff7e78bbddbad7c8483b77294bce9813f943d718deeaf9d5fb84ddfc26d7323592fecbeb40fdf37192c95e431a00ba73e9674d7922dd135398cef4b34892e1b1f13fbd7727ef16f78b04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1966e849a8d51e5fb5ac5969c9a5a344cb7573a13e62f2a5e6c759b7a4a436bedd50a69473eb3164dd595e9e151994b2b58470ef650344adcf4900bb714d4f0da0be20b7c02c1138d21839b9baf14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfd7cb56d606e915b0af7774f2e6c21c99a2cf053bf4aed40487b5c84b69f801219fffa9f4da5f5c767bebd41d7ae49efccdfc257934fe68698b7dd619a2e34603ba55108b04eb1bdd3afafd81a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha06dd6039fa8aa650f2c72f33f1378408723f63499f5582fefae5d5427311c527e9026c3418f123b7bc18b5ae808f1829aa197afed9ad8a35cd089531b5e4163f6ad7d13dac3d6050c82478daa26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he66cdababa85067ee25154ec62d514cd0f473e43379e52fde486baf3f29fd21206ece2c83343e7ec1aebf786a2e04c42e63e0f2bba144c109c7c398693f5b71239bc934fa5984dca40942c08a910;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f357fa031534fa9e4570e406f6a1f645a50559b7fc6643f6101f8aae8a9e849bb6bf360a8be553369b3153629c0607dd49aa517b6a2e8a68a58bb8e0771610194035e418794098bc3f1d66a4474d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ded4089febe7079f207c7d9eb038a3d32ddcd8e129e6add5e8a8ae1862f791069889793d9aadc9bcd701a583bfc9e7921cac7f3f2ada4914a61e5aa5a0ef3fe8db2d6fd7d96928bc839c4cd7e271;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f17484cdd991db450fd7be4c5f1b623845544f1d1da081dda15adf4cc8343b601bbe171af4067bb18e9821ea26a05dda499697fd09588b319fa8a5e8172937b29e99d4a5d027cb384020abf398;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191ab959f267f0851642c548f6eb04a90c326ce32d36f60122aed3c1ccdfdc10f6701571a603615642ac24e7598b9509edb06f5f5b6e7bf37ff0754c86cae530ee6e38b455753afcafd65c10ed765;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bbb06c4efe628491bffbdc040c3d410b3f9db05af05e21a24c95f34bf5c0062de5ac5623778a3b5f77f80cf55de9189deb1425987d7e76de5a78785876bb17c7dd40b49af42cfc0255c8458a8eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be083eb81db936d91da19c8ed14d90c8aa4ac061080c71300d69a735ae690e2b6bd8dc16a47cd2643159cdf8a4b53318942326aacc87370aaf71c46a8ff948343e9f2d613bb135d321430357265f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ebcc06a13047bca67952a656914579610b1b48a3208d62221922153150cfcb6f1c652f509beb7bf076ec329f618aafb18b2f7c078014853e811f70cb2dfc74b8177f664291321701459ee60a2cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142c880fab5c05b669608d4e5b6d62fe9af18d2bb27297667cf4b0ebe12509202839d3adfb8bda30ced460ae89439c8f55c4647f612873d5db902015057652ef561896ae06c7d01535f450bb659b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19df3bbfa55e63f7cba2886614114d3550543fbc9b3578764eb462b2d378345d43d98a6b5a80fdb02936610e12923d9fdd61b4a6de4bfd5e54dc6f561a77add61d6ccfd56bd73955accdfd9df281f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb873559ee96f51fe3d72877ef8acf79f766bbdff1a055e8c8e25c28694e3259acdca1daf3e38311a20177b8e1ec3e09c29c4efd1766448150a961e965ec2fc0fe2d3e1a9f4e8b24d2f721c932fad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bb49738b3003eaa6625bc0a8114157ab201ab6682a89430d7e19d5056a68b15ce47b73e13851988aba98653158e3e3cce41cc100677ba288cc19d48ad1ec840a408da087a7d2dfc55824d3258f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6fd7accd4a9f612abce510dc73040cfbab809b4884a0d6e4cb2745329ec94cb7eedf4285088969dd93a70dc286746dd097f0a6c5466297c6b9ab35f11937b7e821d654868e8d20e0bd38a2863e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55813d8f027cc93d1a260e242fd33189f110c03b3ea1109af4a594690b8c194876601cf55a88749a0197f5186f1fd6f1a4682c842dd38fdc90801b180231a49881b7cf9630678665de0762e90202;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf274c9fe643c2946eb5277a144d695fbe4e1a43551e2cb18046380594d6d6228ab81f1c3f822a8dc36c6d1c726d92e1de31e5d1b4f97b79b1b5fd8b9f27ff18a052a8c137a08517eb0fd428b65b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he69e2b961baf9f868c0662e22e6ae6b2a57b0c8290a6ad31862aa5f256b8e1b13e818f8ca349dc21b69799dbe49f082628a843f953df93ec7eb85dc326ad77dedd8913b76cf92af0ad5f640c4a39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113107e05e0eab18653e2471cb6606e6dc33b140c5078e861c1b7c35c7fb18f0b425ad048df0f29f396d455c6c4800fa9c5de670b0563af4a3a5400d7754fe4fe15e04ff9d71dd961387b73814703;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d44e8620f0d8d4aba23a76a4eb7b11f327ab8cccfdbbfa65773ba9afd1f6fe5c3295285853324e88044a10cc558606ab89f54a58aa481a2679cfdb7fa6a9f344c4633956031e2d756da760862b05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171502502a78f8b1e01792e8e97e535e8ed51c9c0a233275503be14a2aa8ad4aa8dc85337cb2f3039a5cc3af1b8903043917d1c5e307249602795fff2aa325558e2ab4647d292e78e2272ffe830e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50ed6776d3772c6e02c0f7d9a900d4d921d42b8231837dce85e8a098dde62fe3f524ef2456a193e6447bd0b55ae89e176ce4903c62c61e9e800e9c337284508a1460abf0746c3d13a369f48d7e2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138d879d889abb0bd30924e1636946d95076aaeefb498d7724358ef8c635d89c2f1045df46dbf6bd84e98cf2e86d298badeef06993458caf0e7b807017777ddaf7d52877fe96b84b9822523e4a08b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8308bc0e10a5c3d1660b502db7441acd5203046ab88fadade993ded6ad7a089e41a251f3044316e57aba27e0f4e5d68c48cc0dd390e8c748740d41dc0bfa9863bc7d1d7d397cacb4c7a10819c1b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4462c165d3bd56ff575689eb9540ed82d98eaffc700747045775a241b2fae5c758d0b5c7a1ea53dfa9b683c216c417164c9faa021add30a9ed4882733188e4f37f1b62339bd6b96d83ca9fbd52e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6defd7b5fc54ed653a5c8ac46cfd286a6510d87163282aa4151fb0c673e11bd5c9e14cedd7d040740169b134ad4ed4a39b0033981727cdc4e9350ae291416dbc01cbf11b1d46aa70bac03ec9aaa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d578f78f07f93f8871fe88fb6fff34162161b7ccf88d783db0af078da422e07c65871fa4579a51a95d7bb3e0dd15030d16becc4d8986090e6a49499a4adfdbc8d477f4df7932c0ee5b775910c935;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10201c7b0be4523c32dbe7193fe79dd8c22a9912ee39dcfee6a47026ea99786526eb351a4bbfa89b53903d0855bf8f36582536f4b7d77f89b37346f3991c8be8843d863910c4fa268b8b4d03d0e1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c64fb67c29ea62138842a7eff3d4a007d65508c269b9d9ca6e178ed8697fb32e3383da8e0e80d99a8492e746167d28f9fc8bdfa124e93a22705d2df20bcc8d5961f4403c16dd0f97a389a411528;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd68fa333becc935a583a29e80acd1e7d5cfee61ebcc7dcadf2f6fd8654f95021d4e488a0d1607ae9c3eeb1ac740c6535155fda0e05cfeba95b88ae086f33b73673bf667a93365dcb8125bb257be4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd06a724eb16a60e5eed6e2c16148442fc103fdd273938e3177fd7c59b56e5289dcfdbf5c1d76f82cce95ecdbcb56d26324d4e0db8a2f7dc6b86676c2561b08aa8a6a97d8ad03f87ae6065d448e0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71e46983e275ea79439809a19b062c71323172de6f93f7c6df9eda0bd9dcfb1c6f615b67d2dc6b0550c58342373d40db0e936e302947c48445291c526c9d531e616fdcc974ea00a72987a537528;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e7e19ed12765ac470dd740ae6df456eaebe1da986ea5af10229cabdc7565af539a5353e8305816d59bfe27ea6cf8e4ae89858c35e0515affe472109e178095443d13e8593ddc00018bc8b606dd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5734ffb5ce068e986036627387718481d325ea00033a47009a96e74ddf41905f8fe2a7b6af1a5f308b1f20757c3f83ef55d20a62a0a46481464b24f797cc77b4b8ddb3c6f1bb1ae4b374153a2e80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162f743b588d4f238b7274c8ea6cb8427463fd8ba5ecd5b5fb2eac0eff538d0ce77dded330781dbc4deaba4c52189eb05548b2b27bbb7c2a271a01fa1b6833356d54a6417a822f522ea74dc5460d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1666a34156f45e75ab6a85adccb7b585e2ed884dbc00df8ef193d7fcd7cc817c789c29ae9c0c2ac24004f1d9dd5a443f6af7b67d6fc8b67dbd56101a70fc3a213c2a3e7654b081d27b34159960663;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141707e819abbd0a5565b6b88837ec14509960ae46902fdf96421f63db0576ce3a301ef298f2029f7db6dff915cd1aa414cc5c4cb9bdd402b718506c0b352b0916f86314ba7a630431e76d0b89c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9ffbfb7c555b5e387e09f713e09bfb395274863ff6c16f004305de08528de11b4d01b97afa0ccfabc259e2cd842ac672511762aae3400faf371a966d122eb8ce7783a2f742b4d76752a91f6885;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a90bc4df8722c4121de7e8c62b023283d44829e3d2a529811c31fc8bbe3a11cec0f019de0c357495cdc91b945bb2133c070e4d7b5a1f94fe365b4af1ef15648d5e05697877dfded2f8072f6d6704;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136b9e5754aff74864e9bfcfeb43e870d5a21659f79298834f246dd249d1027f698ac87bba4fc468b8bcef7080994725c14c924844172695deb31530c389621ef937ff38b80524487d4662295d618;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f93b994ae8267262fc503b8828b0bbe84dc9732d9b1456051ff1d464ea08d87ea8e856a816af1d348841308eb74b759a85ab8c5044ac8240969fa66fb457ff5ca6442f4b3e42ade1592d3d9837e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b7090fc2778f69e24e6350b8ababf1786d25602acbe4ac990862feda45e928b8f6257fcfb63757c45b5a0e9bcbc911bd254277fc2ecb21ead25f49b895673d4914408b0057571791c8a5abed0e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111c90880346fc2c1a06b4f4d906f3fc82feaf6b21936f569e856fed71a8e33a28c41ffcab5b9ed2c247fa500e0e2a50c0685fd57c51d486bd8184e336343316dc80b1d5dab0a691bc48086d15898;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1929050d1e9cc53fe69c7e29bbae7eb3f9a5c272b842a3645628fc9d870a6861aca57180d790e8f3d597a02cec85933e76b26040400b23a04202f2b0a2e898e84ad6bcf912d868c62d5fad6a88e87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49708414328110bcf4efca0ec23a6c1be2357b01dd60ee4b3a8c0b4634a900682cf9ba9ed658cfe4fd8367d3f3028af7d4e97ccedb84e59613fdca0d0935d1f453db6d9c4573b2ae87e569a5181d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h734bb79eabfc7d99e0a4fee67acee442560eb770d19616b57d090469dba3a5aa028d54baf47bca2cc2c5e6e886a316bc11d7a3575699be0e2ab30ea923b5ae2e3efe29f72249aa5847a20d8f5f5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124a1ee5f5362a4c1dc5a962314dc40f7e66b8e72d330c57ae4a5c5a0bd20c67d3b603307a91133ebd4dd16ccb8a00b605da47ebef7e2c1c913d8dbab8a875ff5f50bab0bd450ce7f79785cfe4ac3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe6f9ce93db0c13b742803946e643eb9cb4a555ce068e3a7d9dd45c5f140ec1b909a81e18d1c97d29c903f43e0d8ed8311c6fdd73a994754ac3edeb073c273a924769cc8804efa107fe13cb2f9c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1557a2a57cd2878942b190d17080d82948f926723b11a0f357bdae77357799dc9886f21857d2101c5fca2343e6532b8f4664c6ad3db6a829b8bdc19723a4a2a64a8f80ec2bbb7b5b9fe9e95a65527;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b59a8665c6b7c73dd5fed4332a6063a6cb457de3e659ae3937edc3a5d41254a0757645ffa5c846778450db1915a868e473f4c4264aa3dea1fef37803885de123ce33d4fc6f08d36c770246db031;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e757ff72c9e6af4444b161eae99743b882423fdecd1d81c40b6fce8095d8f26d196bf22df95d6fc97e256f0cac50736b4a69d8b6f983dc055ce414872fe5e10cc17965dc8975bf53ddbe3dca1e90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cfd7b278aa9fbd698418bc2da795105aacca397f392867f0d79800bc1fb49ad248e3bafd93b83b73aa48e0adbfccd906d280fce344d3d2f4a721c0c3bdd3a9fcf051a517a0c4b0891b8a95d5ebb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b72b361fdc75956ca0832dbe398d1e0e793670d0010a635341a50bb586d1dd6ccd5945e9e46074380228c1498b437c7b22e2c4cae2fd644b0db72c0057939ddd8487f891f5010db8ccfe5cbba27b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1999bee2a59ceff4519ff8631da5fc172f815f3e86ca00278f2c9482e49cea637f185edb801973bb1fc4ed86afe15bfa6a8c8229ae6d6a9107a4397a693919f1e26180000d82256106928cf4ef497;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1185f93befa643b69522451a8a66ccd250ad6aac8c206ec9bc6cac91515d06e26fc8fa94399069cabd811411edf5b459cfa0fe0b0333b85e7d7a8fbcba969ed521dee8569558e006c7a01016674f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fc78ab78aa65a7290275a974c914306b0a8758cfd1323a61f0e50ee0b06de9c919292fe4ce86603f3659071d3d82890a8072d74c9e44e0c892ec1f4833dfee939b9a4569d0773a8120c0e0e0d80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hefcf5b8bcc86aa8501976b0fe0abc822b32db95899309dea39eff111ed22af7a033e63facdcc3208b89dab06095b0d5d9df245187ab8d7eeccc7d133530958ae0a2bad1d9fc89dbe4d0d580723e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15027e57d2cd23cb339124b9312edc223200d6f733bd30c554b9aa8d60737bbb108a196d12413bd61ebeb0f3e40c696184226caea92974faf2c8d1858f1eb0768d49fc26886e6d81f14409a0b700b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13306a8d75e382f4fa28d5ab6eae3d9d5c0f3377299012e2ab9b9ec324626a65b6a4d4bdea613510c81b3d2d08fb58ca8dc584d9c72b2ac4be446b63d9b9978452f2194c875fee0a0c94972277e98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab23fc47be8b337e509b0fc2ff81846f0940b6801707bff51e4215e940cb746dd9235496d35e3e5cfd82110ca9a3db7cecd21f771863619d17fe7d880eb02fcc625ac47863ad2ebbeb6a19f6409;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e16b8d1a99a04de12b10a69018075f77b91f347c77d03a8b053a664ad1c0c29d4176ce62512919f04efdd48493097bc973b2439efc6eea96f351fcdddf9164486db5ed584c58971c48324c3221a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3838a11b13011bdb1068952244a106f644f1722a69621f4a74b1884da16519c256b2f928fbd945803761aa7f008ebc5333e624224f439a2184cf469869f1e0b93531498f07e014b0ae3895a2756e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125ae91ca540a3b835cc7e2176a122051ebb6fd236838b2a5b972cc7f5639ba2983b8ae2edc9aab9693cb04dd88d5c1b3576b7a4b9c554c48086feeb0ef4e2dcd83da327b00607785cae59f992207;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c1f45b887963e777abcb51d35599dfc95c7018f771629294da551fa4441dfa1540498d32ed28ec26e188ae42ce9aaeb870bb50b55a5e2731005ee6bc99a599266240c9b2f6c17d08074d1f291ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ad7fe17938b96a3710891bd62a86cb2b363b4822064689df40e628aa22a3bae91623b1ef7de978fe7891927a52e57680650e960c213a3cb65275f7d66e6e532f15cee8ff2c8538ed38f80ccdc31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8d0a9bd53196e5455f29d0fa54357cd055066bcaaecee500f2730d4df1a3872eb8112ec8fbd9528130643f3f6f431d18894d3d464c3d224cf0e6414de4a5eef339982f42c7c2ff7c8ce5de212b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162ae8ad6f7161f7984bd9590805a081d5dce3ad7380494a506ec3f55a133dee4a4f7563d1086c9a2fcd9e575b19a84a572658db9f3087fb7c3841b2adefa8b43e452c0d7242626022527a4eaeb7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a2452bf7c0c77ff856273992bf46975b8b1d91419c6f9c70c37e83aaff3870e67359bdebdd8638942f7c154ae40c883bc1d08db843b4fb7c96bbdf4364a358c3c46aa9c0539869d0914d0156f46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171c7d5688b21f29e3795fc49e84ca74e568e5629a34a212034ad2afeada2e1b5b3caf5f5bfdfe7810addb09406e2bff748022af560f48ed3399edda54180c76a536706bb4903b1bc892a595f2fe2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d925333a379a0e64d3f7c3cf85509004caf31682f16f51aa9a0be375a9c2d7f01fbe380b8b0ed2c51cde88708a3992b63b1b7d9f6933cb57bde114ea95c22237e11a2d47236e345c40f4bf90d140;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108d44aee2f98947c3ec670a2b91dac3fb06db0d34b8f043df6271adcdd56f089800593ab84bcfee25331d507ce27eb1ec6df9e1ce80e8d220894eb694f68444bfa7a6f514ff0e9d4c40ffab04347;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf96f692a04ee77290d37d0d6bab4ab142049a95600927505317fcccc7a7e8b34c37aa3c61e78d2e343a22fd810100db3b852299983442ed198a107c9bd92f47869a69ea10019cefa498fd54e352b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ca5c9853986d46ef0e2f8637f7c210edf528b9636be4d418870851978f7d24908116f06957b9452b8984296a14c42cc48585a92321a333c2cdfb1d050a15b22c68c3ddf0936e5589ad69ca2393;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c9ddd6582212370190b1027e981759481d768987519b508e49fa55a9ff7c7710d2db9aea7da18626a7a88fe67ae6282face0991eb1a5d98a9d9a4af6e4ea213e744cc24c5a3e43594fa72edbe51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha323304b5db9a7c6298f3054aec6805b7000ac723378ca17e7e581500ae0476bc928eb5d61e054a4d9cdbb81f391082a352f6244edcc1ab31074f0d3a59de4c2647d93ba0dfd6d35dfb36f1209f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183e95983680c8d3413f49161a351efced07ee91540d3ef981dca29d22b99a391b7a35e2baaa9b0815b5759ec1d71859fd16273523b05abd22c7aa7928167f71b49b00b526acfbfe0a20907a8a4fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171f9e9dd339a7ca8c7020ce82c1b7f73564edb2224107ca6fafcd0d3395417874738d5d2d5eba9605ffb52d857ded351186ffc8e6228a1c2e9c0f69e254d79de6fd49e2a50f38fbcd0591667715d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d3634764b613eea20803cb5315e8f154521c6ccd621b4ace450e56de8f61ddaab959a79f839ff266d083ecb948269bd2881bac9d90705fb110cf857f3da3e401db5c560b5833e3e33fbcd666d6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfb1350d48a6c92b110b3ec1843eb0a0b7fa82f721cc9d552bf5cf0526536ff2ca9596b8dfd2fee029b49e60a9db8d17f1f4bc6383e1a2803ff206bed73065a30317fe4dbf616d66781dfb161df2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6407360eef7c6577fc450dad9392dff69caf73b3b3481ca445a302697488f10590948d89d5f24831c1abde07c2508c49ac88fab48a851f40619ae7e3fbf84282ef4d536b14e15bcd4721d7c669b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0818de69c3b1f73bdd70f82e7a59a1b77d581c6758d1c5d33cc98f80a9d3064bc5843ea6af04044ef18fc2826444132d22e77d07c5ea0dbc0d9fadce2bcea5b3230f9b696319400bc7503442a38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae6129054926394b299b1bc77b8493f87ca8bca2e09fa236d7e10a5be1ef6d100095feaccc33123f7bfacc48149ce83cd1045b58cdc1b80498dd1e2fab4a2075eb9e4b415d2ca67edca8f73ba2cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a53b14ff7f89156474358824d8534f662a7b262f33ffe0a282d568372898fe481cd266d75fed3cfec53f0f2daac2a8826cd69c675df13e6dbea684a10e8146f01d71060d7839bb4151e8b9af7a30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93cf3b62c39cd22c1e7c0b29277e16778263fd56207753e424bdf486a80fba81f7242f164514be1aee8061355126240ed5fbc88cb8eefa1d2c8477b9fad6b7f7651f5aecd2567a72d5d05a366168;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1691a0ea6e4332af553123d3a38dc77999131a4be169bcf4d82b545b793d1e2153e28a1d56b8a8a46648d2b19881a444d9f30eafa1ac94347fc58359260660ab0889b8183d55335e01411cf198164;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67f3419e0766f96322ef6abbacddeed3788b8a62ece4c79b68eeaa5fe101e04806b5eb2eb1180e02842b766a0766e29b8b4c28da252554d37d78ff2b822a68e71a5cc01582a01fd525080f51a9b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40ce4d3c421cd8355475cd780fe2f116afcce5a2ba04f439d33408de29da5690dcac9ff98440059b24be6fd7d8c86c909f3c0b5302e4cea553735cf2b0745dfc3638061169b0cce823f0076071d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180806b7a417765aec0a7aa11e6653f341df3df032b1896683b261fcf872bfac8e30974db51f0ddc28a41d250a14dfee376e3f6bff604c0c8f92bece7e28fa8377d34575b88ec814be84ded81ab45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11359bef928b832974e5eb1aca8bd38d72793844d5afef9bb8acb445f8a6e02a98e39d4597c8dcd3c13add814e5f7a969b831c48066361a799a61ad2fc8931173b05c535605fcdd905bcb832e860b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdeb7cc929f9731bc6d10f85d64c60d83515c5e25e706b1dcab35e9a608b3e16575af16c641ad16d6269578adc8be5f5771853d1436b9a05acb4d7e6e499aaeb4f1f97985db02a07aebc56b350700;
        #1
        $finish();
    end
endmodule
