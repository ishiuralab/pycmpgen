module testbench();
    reg [14:0] src0;
    reg [14:0] src1;
    reg [14:0] src2;
    reg [14:0] src3;
    reg [14:0] src4;
    reg [14:0] src5;
    reg [14:0] src6;
    reg [14:0] src7;
    reg [14:0] src8;
    reg [14:0] src9;
    reg [14:0] src10;
    reg [14:0] src11;
    reg [14:0] src12;
    reg [14:0] src13;
    reg [14:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hadd56d140ab977102b033baf68758399b2030718eaa53517a7edaffa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6e2b0a4cb6449e43c7c7ea42dfc38ecd1f622df7f940dd0b4654699;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f5210fdcf16234d731db6e7dd210a445e955438d3bce9e059652d00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h379b7997b4614e756e8e4261d0bcb227514deeb6d7ace4654f4a5b3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4666653f4a5375a9ae84a5399d8c7bbe1f31eb527477fc6656e3191;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1253c70a35b2daca9b043852d6225e9265c92a5a7a8853b3bf066b7b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a86c3d80a3cc25fe52121f8b7176f989a01dcca6f14238ccf8bd9af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2fcca9f0018ddd5fec27fa86bde42a7218a4bb5951f6807a2a5f179;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heafbe91834ea8d0f2f9fdcb48a648bfd2c793427d614bddb4cd69015;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cec7726200a2631f79d3abd19b2e40443994b917ae471708f8c785e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13349f10252eda04972b7e2830b8f801d31a688a8193d61c05cb29781;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h913431a0c8e81d1540ed61da55a3c6605dedc63174b33459f27c1afb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5779332e5a5ec136f2ffa6d0f223c9a6b771ce43dd0f5353b95ce8d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3885bd2a0c7de8aedafc7364aed57db223dbd83f7997202a09443704;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1992a7375115425816acb44464812d5008204ef3279263e19755c5529;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e728ae5b8cfc4a20834e581dbfd0a4765ae37d476c89f8f6920bea6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117d5d7cb21eefde7fbeb39b08f154466e43dc4d42188698efc552aad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hab6f1c5bc8f0d80bc232ac28fa72d396674eb1e238f6e1c9363abd5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5fd2899158be65844a7700953c5de878d39da575daad27e79f6a886b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d9a591e46d47bab37f3e1d995f49c03d1f614c0275e104dbe4cf9ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c7939d639d6d65c586edcdf40c0932b3a6a7fd7e9a59c3b66745aa7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdab843883430a808bfead6c1e76d2d93aceb93b653f7f2bced64054b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef6ac63a99325c7b12eccb8a83152d26125fefb82dff627c3869f5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87a36d2cc36b206637b2b1133773b539764986dcd50b6e2e9c10d4f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e95200762bc6fa159504c069a6762ace62fa7efbd95973e912e2958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1c1967866bfe37e62a6e9af7bfc55dc9ee68569b6329ac8b0277aef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a3ca73019100ff8560307609adf05cc2c8b79214c7f1b56def5128a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f06e3c9505fd7dad349d67fdb2bcfef105df10d56297a7573dfe3ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f168f1f30808c2626f202b0d675a07af36e59e773f92e7b7d45191b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9887fa01979eb7eb896829d4f9493683572839c4fc0a826f07bcdc58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aeefa0d77b0e8f952d120181a5dd6dceca59d77d291747b66223445f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f9271223f239df5d13b7776257a10d47460209c113a44cac34ad2fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d7d55f1378b8be042f03646e455afa760b95824c5415978325f9265;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6f950cc6fcb79c49a281fc23f951851808fd7a2296b395d177236cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h843113e2c193b775917780facfa66ca5612c54baa234a22a92132971;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d633ee0886dc557c037b526e42978373dfe81194ca45dd8ebdc82b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b81e494d9dea37a2c002903d4c0d86b6f1fa9ea5c11dcf668cb93054;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1819b41126dd06e238a02bfe6cf07841045f6a52c474a6e442e5f55b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1965627a389e00ee35e7efa3fb9ae74e778a11045827e7f5ba69a3928;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63a795c5b4f627527c239733ae7fcf4abee5c3e0c01c4a0a56044076;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11433fee801867c42565e7c42ddda1cda7e66c3d7bb34832ed3410bdd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf21e205f47fc84d2cbdacf33a522909fe602fa79fb4a68d662274105;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7456deaff87893b9026a10c798e1ed591b22d2b2232309e229e46a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135a034b9c0bef245d985ac6393207256b994de3ceee4846cc3c27877;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb1284109369dc6a415521312c6bea52c9ca61623c81dca4e5fc84114;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c44a846cfacdabba3f23a967be411edc1206442cb4ef4136d626075d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb9d2d097bdc2a346270a5e70b3fcf2e0d187007510f8b7a4b52bc01f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ade66c8ca5a843617bd5a38de079c65b43e3f0244071b27822cd9a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1067ab158689fd4782449b2f8293e40a8db50e26bbb9860b9e6de85a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb4cdcdfcf7a532b427d22a9339fd5490940db8bc2edbcfa2be2b32aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc27ab7c4bf98a8b86ec5baec6e6f76d49af087908d9fed6876d8291;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ae3024ad76d76fae03cb4db4a1766cc7fb3378d0c2c607bfefba52d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168fd040df6cb8df0871c35bc3cd4935ca4223675954d85124feeb773;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133e0ab6bac02233e35783cad9200027998c041c8fddc5ba266e4f97e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7abd3e33bacda2581cda91ed352a4a6c11f15bebb03d8c48bfbf53a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185b8066c611d449f28860584fe3f677f50ffd036059b1f0f2b50f1e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e215ee274e94d22a049ea13cff6871313d20a674e892197bb4fd075a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174131778b9f7204be028f0ccb10570bc3bdf7c4e4cd3d90c5db116ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf473f44c50b02fcc6de4e385baae12a7e2e379b6c32cf7cdd69464d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a7a977402e59aa02f5b6e5c9023736c86bfd3a5b8de950fed6c01f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f84d17c5e5104420ac50656e3959703a3250be29d961bcafecc056ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2110cd51ec0bf2a2472f364a6bf0c2d1b93fd8cf0f8a2f2cdc87e97a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hecb7a678eca305dac6fa904574012d7fd429add65abfcd2d5f6be6f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac31ac988b0cf5bd6dda3a75705e674636e2035b5d705d443cef4d2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hebdd3c8bafc902b987bf95099b353489818261584e6b51eaa96ef327;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5df2f0f9d567818e9e4659ca4b4e492b6f94cf5236cceeba8d139441;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41549386ac6ad191fce6d134b48d4c5f167adf187ac8fbe7ba61db30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf50bbd8fc0ea59219b6f7319bde522224edfde4cc7618561066865d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13479dd73914e7d9624d4a1abc70665e1f6fc51228c25b28e2b7d63e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had377b73d9472ca2fbd5e5ebfe6b7d99b4286d9b77773ddd1e591e51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hadb69ecccf15982a0a1e101a5698348120d1873af997b253d7f001bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fe7e6e195b98602f021ccd7ccda746118c0aba358a73610aba8da44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef189df02be68d99bfd738d0483e6db5abd007e4ed24db0e143ffb04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbed3ae113d0595a90d882c7a48c56ee302b9f938626f844c2b032ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1665b031018d6d7557bf420ac829036899270415e7ede25622931f452;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2b258d13fbb9da2c018e3c986297901ba8650caa0ef60708c8cdbae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8da9f2fff649d9898456cf9a1ea9dd05d84b5bb289853b3a53fd154c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h202e53a5b5e7ae5a6744c07c9a266707d538d92b8edf50a84d81f7eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1978a90bc831367a3c26fac7b2a56e7f5531c3dbfeb8b44424612aff9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75c9e561bf86f236b855477daeffb4340a46d8ec1b98b7eee9531cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h77982e5d1946faa297990f483dc837e5223ef8966172e231961443db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd2cbbd47b08fd0c9d06f44cf65e8bfdde7aecc4b570356fbbb3e515;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h750166ce56e03eac4bb14296ffce231472aac1bd7c8d225f671b3765;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf33078353133c3789f00030b08e70a1a7ab6743b11b22dd44804d69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13704574f8291d73df9ed37f5834594f4732ddfab1a82c4431fe7b70a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fbbf7df1ee1cf255f611f8b3eaee286b5dd22ca3e5c17dec6fdad979;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6fa234a6f6aa24898176e7ec43054b07125073678d6813d2b322892;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd491e99d8854d02023e8e0f0e09834ec78d87d4ec4503b50173af5a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1083e37981e335f00f333f1fe577a2299c21f4b8aea5bd9e460fcd126;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h97e3bc5d31195d4a027f844ae78ae3227db41152b5ea509fc34bb971;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10684571ef64d94462989d6b5a5b7fff10d4deb8bc14f0cf6516809f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14867f58b162f268a93e79b84c1212a98bce4019bc8ab28362a579e7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf0613e379a4a10d317fe52c51f66b2d8d04f5179afa14ab2b6cc6fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4c7bcb426c19c141566de6390f4fcffd67bbcba20fdd301f707d58f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a9dca77e6bac50d4a91917d6a2af4933a2f26218c6ae1142fe5cdba5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157cfdecbc8bd02ff098533ea55c24afb67c5cc946fad11ff1fc42871;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120f931124494822b5943e1b97c5b31baaaeba8fd88438e20021b7249;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h261a208950b2a1f7dcb12b6068bc4e532b55ae3efe96c95f35e387b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he03af1e9951a24e6f7612dc783a1cf86b7a8e164eaf90693dc30357a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c635e53a0cae2c839c5620a71052639efb0596407768a1ca1ad8fdb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae5c99b6a1bb8a6368a9314ae0dc9c74ed2fe82677337482d70baacb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha906bc0aedcdcf3a45c58153340ffffdb764dd7ffd54b8ae5bc28493;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd02e2699c5654bd24c17af65defe504bce1f99028860b35338babd05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15aa4beb63073f5aae35bbb391a10f36b0cc9b3a4beb87755ebcf8add;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b93c75449b1f556c330441224b068b905c42fc0efd6b66518d0d13be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1f8a641514bfda6e0035f07f3316bcb5e7bb42ddf13f0c8c9a1bd76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3bedba3061f16d4e4ca2657500e792c5a2fd5299b38a2ccda8587cf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f66b3915bfee06a039aad0c9f2cafce34b192d9db3fc7eaa534e7d44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f9d5505e304d80c839193c2112b7c1d5dc82b60b3d5f4c654f1fa96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11904841858191126eee6740e0cce6b95ecafbd0aae2eff17e77493df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c195096b06e2298aa32633a264f287ecab3887aa17c53518ab7bf2f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152fd3c115702c91cd88f54ea68618a05701baf183d2196f8d1d1900e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59585d16c722a64fefc86308d09ae8fad25a755b5c9a7849ebc821ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174e36efc694668e7e1145c73978de6cb63ad5ab528b3c43eb4306d00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb835bf8e7e34500df1d8915ba3d1b03279e479ca2715e2443ddba6b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15af8630c633c3684316ca68964eccf807bc0e5fa39485173e5fb8182;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1661dafb5dad1c2d95032e8fa837de2f538046c8396377d0694428746;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0e7ee43299987a43973498247183080d6876dd925db89a1a28ee57e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f87e82b1a9b94b484d9de79c1eadf2dc8dc2d64cb69b961491422b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ca8da3fabc51ddf66f7cc923ef47e3bae8c5ada89910fceff5b48a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137210d77db685fd5eda081e2074e52ae61a279d5d301bfb2fde9f39d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d57547cc5ce1707ecba6f489ee8ca9894494c6d32d06d36faa6d807b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h817377a6795e463a102deb778c8d4bd2ae2b85c6b3050a3da9c40bf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h453768e70d568e27fa93337c80e9572720ce48abf8e22d7cfb919c9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdbb104fc4c1bc1e3fea3b5a745399800249a958f31a4d0e4680cbc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h166b1d6c621f59c302173b87d988b368cdb5e83f30a86bfc6b9c3d4c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195aabf244d18f76cda62040780aeee0cb4bf008535b7a6122c8ca2c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e567e7a8f75efa7932f2668cb1f6f9491ccf8d4db733f4641ff1cf32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181e6efb6625ea0b0b1cef98312faf7991411dbf1cce02b3159fc1c21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a5e7bc40161c351ffb45f1811e230c64213885fac880e47a0cd3377;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dc451f79aab72eb8c1fb83b32eea1df940c53ae19899aa93e836ab5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181fcd0f17b9aff8febd10a55ccdf7571d2180ad449e724fef874cc3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ba2e189c4f306651304ebcd32ae636a00fbd5f18ee7ce23bf316eb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf1eafb83ee5ccc1582aa11d92280c55eb997ade988712781cfaf36ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17aff8b790a3c9a5e7810366da45138f9296c46a280a839b63fdcdae1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15486300a7ab3170ca080087404765aecf37a1e8e7ca2f23696c807d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d6915c755fa2a098928fdbe7421a097636ee100cc0128e373fa26cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16078bc988fd597de532a97bf5a47ac8ba03f5a3beb6a0d6adbad13d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb9dd5039b94a8ce37493cb2770a1fca7709cb1c2de5c28d49870dda7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haccabe65c089972187074d51d446f836657f20f4da6c60285dcc1516;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c76b7bee3fae3c7a89348c4650a0e20e9abda6c9f39600f07c8ba23e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fade108763e0bd92a33dfccf47bae91616cb2f9e99abdbcc4ae9ac5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14849b1a47fb20464f840491330d6e35bc8202acc8b405022e8b87d74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1485efcce6db864d9a30b6c18f2965633576d8d901b3ce2386efaf87c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1630545d2b4808e157fd47259d9b5b4b7fd7494038ce3abe91a6e21f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h160f059b78772084b6528314ee648d6470dbf17e19d4e6ccdd4d8d7bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hce8a3f4eaa433c35e9d7006818004b73deef47252e1f2adbc2087d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6e1bbe475f2a7f49b077260ff0312095d7ebdb403f00cd5ffaf34bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b7619cee02f847674ec7f047625777a657cbd3444f5ab0d161a837a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4d65aa1e577af82b5d73491203ebe3ed329af500271effd2e0bdf6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1105f8661fb1ec7092b2b338c162101bee5d4e4ae15daf76df9bd3154;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a451d17847c42dd49b825e2b7a18368c5207110276920316144fb0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9b873f47053fe61d309d6f7e4691244d939547295d6ffd463ccf435;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d49967f7ab70f980cb6a5b9e3b9a5c35ffcc0e2503f2de276c8a66e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eacfd29eb1ef241cacae50fe82c377339180aed697db1af1858ee6a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d130d4f4549e7262dc781bdf7f28b60667ead2ae0a42c22a39cb8b60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4e6d094476ce35425646b7b576c809c0d5b61cf3b6ace133f802b61f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10824e1de25274ca7f75fe117a5222ffb792267030a105c8d7539644f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28679d5f605338d2b82e6fe1454f11b0f462d19a9afdd86731ff5017;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfdeb4222467ddf8d29f8c96ccc8d6441d660f6f32e20b18bcdca6f75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee2c6b89cd9212fb33d0cd61e0507f0a2d9907d0e3a312b9dfce3188;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f242e9e623affbd36d8f049378c390109a82660ed4f03355437b6da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55f9c38ac9858a8475232fc92b6c4c10a64ec04740817ff7f64f097f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c8d5e89e5d7b8915860f92628c9021a5b38b9ee6d4dc2f2bd4f51c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a62ee1f5a6936b73b9b97d8515fd268ee0819e5c6d5c4573c00f95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7ec375d3ae7bdbb028558c9639c693c5afb1b12813716a50b9ba32c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he83313d9371df0d8598a2b26a71b03e43c7bb2d2b0c6a89b1614f1d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59911ea5da893c049861143c7c0b6fcef7aff8b94fff7304d257d97d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2e5beccfc8174d6e820625ad3186b3368f2ee9848f8b37b4c24108;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ddef2fe624bec5529b3a640087834352461ce0a2da60c4c5f1d2a1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h112d2c2fda1cc4946dfca75694c136b5fbd72a8ff833a9240c032c07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa9cfd95da258ec162e1421a571677cb693ab3bf56beaa039e8879db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a564c651dac2cbc31f0967e25ca884c002d0058a963348b67b44f102;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed6edff2c9fe945c239665bcc26627d9721561d7e5d15b5e7f17745c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h812663042ba09c065193dc604843a52f99eddec32fa08cc5e2f6c553;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1939c5e7f21e1ec39f1bf8d9ea8c8238df32ec2c2a038486cc053348c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ae2b83c0d451fecb1ac1d3c68bd1e6b05718bbc0fcc4f189de6df706;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76630e6785db028cfaa2e9221e11479cf8e1079a05081477f9cda39b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148b194cbf42bc2e6f452978b7c7de2c991aea4f522c805a1046c3341;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd4a63c010a73dbc01c760a60170984acb882e3758a481eb778558d36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b82bf5652c6884b8e082b9fa2208bbb295667e2840c717541053aa6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c864b342ece6b9140d88873ae7e1204623864ce0ae669125e7e6fd23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a95e1d099034863330497e80537585705e29fbb4b60119f521b7d3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h704859aeb038c293a437c93fca54d4f821d9279580ccfce75854ee63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c57b80fcb69ffdb8bda4dd82f5c9b52b6768a2de59ebed77b05b186;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aee2a5d800e41eeedbc4e34b5037d332df844b093297e7912738b259;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f8ba1cffe6a0c3c84999039dbe909aca3d5e887efe9c639c2d14d42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9092667c97068e33589fbe0df995d6296c5937449a1aabfe4cf99749;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f3edec191a35fe0faecf9b6c60643fb82a1dd3f3102bcbff8a74f21b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64d9ea62a63b221e87c04040f2c2d9de01f3108c9a569480c6b403a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a2278b6a326483527ca02479bcb053ad79141c3210cb26c8c0b82d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ce1f5a8151388e6f0a0ca634df6924a14048aad0ce5c186ec0d21c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f0480e43ad6e7c0c463dfbe262e17abbeefebc416e72d6e1940fa17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1c9f54eb441bbb95d4fedbccd858a4caba709a599a7a06fa67b2e4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58a671b67f778440da0db3e788bae304f4d2743c1b1235c18f7aa74f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd2dde6c9207dd071459fd751fdb5f96e84e4860f9cc75aabaa6f05f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1424a7a591d5839b519f124a2c72070d3df6844a8c75df3116e9537e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9960a8ebc7710082f39381a3542c7ea342b5172f394645f4fa46ec4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffb53b5c74c922759e28a6f39b59e794e760d0f117f891b17aab086f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2ef41146ca3fc354c63bf1121b22ee0574cff88a759f858b55ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b967d0e62fe036d90efdda84985e346e5ce798b264b1db2913e6156a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c1a3d9ca39146d7deec2172b469118ef038364b7f6ef041e1e8d2a20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h102eb3e608853d3e10d0f99b91b1626803514698b8a125f4631e949bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7239fa8aadd332de1656eb8d59a1118a5e9148675eb9e36df359984c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1471e955e61ba409b87409ccdb1e0a22af71516814b4d26bd962c9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a97c5fb54b7962bd8d8848ac7a1e8641932f32f26b62b10342af276;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac340485adf23d17cbdfa2d69e230e8e4f4ff8eb183f1cc2e5745973;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61f99861b6d1c6e9279dab4c53d057f48af048a93dacdc8f244799c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d857cdad191e7271d4e9bbcd8eca5808637c0ab3aa5fab057d8b15fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h25e1eeee7faf178a6325871fe5dcf8bd06c5bbbe72638a475cd0ff5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd18ed7729d8f7c42fd1ab6b1fd36122f8ba7dd72028afa7b551f954;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1795387b46d435ffd700b56261c9c8885fd37e6c639e8ce64051090;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1111c35d8e0320fb3b98748e9f25c5e17be7ff4d120efe96267af6afc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1af7055d9f1f172538ec6675deedbfd5e24df552e5893ab3499a8498a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87db6aab44bc0ff2245a891f9d90fa93df401338dda4f07531dda74e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b24e2b1834468047910baeec81a098d7456d44b208c13858dab4cef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74129e45766fdaa9739583ab49a762fad4e528c9e5314b668d047c62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf636751418a9679e3a643634c81f898a74a83833b5b0a782d2b1ae5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd8f50680e50b6dfb745785a941440d4b8b0b6d2d776786e956883c40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he53f4d387802e11806b9ce9312e921d10e1f83446ec1b22da03160fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e364b42d26043d711ea0b36b268f81d5e58182a25fe7e950a0a8608;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcbc8dadc1228273ff964ce607b371e80da0494ebcdc391178c5e5db0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1926d07fcd04099b736fa2b4525d7a1f3fbf7992576c017b1ac5a40d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc6482bf031a55f2db354820fcce9cd5d3fb8b98fd3b87f931ebae137;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8db47d1da0d44c4d2b4f8fbc9b89fb20f15a7d7840b2c2c71bc896ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaf4e3f694b18781424410009c6b08d529e4ea635fafd5b511fd052e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h335bac94360dbb7915cc0c6f2a9f2bb43f3ad3d15c0260057bc75d99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f14f98d41eff5f723d7cfe08ace46ac43f8b6bb9241b0328928bd3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18778867c54b595384659410b867b625b8f3a0af61c0fd2f19c128718;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2cfef39cb8d6b0942f1ffd57ed5512ed6a1b38ee169efb55f84efcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef4da900691dfe001b39a65c16d11499d0fb50f9ad951a9c916eadb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b4141cf24fb8bf842ff611ab07e1fb2fe4e3a37355994839a965578;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b832522109ccc157de74969e3e77dc59debe509e83329df4566f837;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109e10a082e2c6b69a24b9387b2ffe15550425a5135b863c15bf0e2a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92db2027d20b3dbb8d507992844eab9aadcbf7584ba84774e6518bbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d373a14b562ddc856e18311c1a5218a2087a34f7619e84f32abef6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h845aa603d8957246df344dacda27a31c886572c1c0b53cf4c837ca49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf09dc7225487e4eaa5a8b093a430c2b617cd98fa0ea78af131594e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18bad7105441024bbacba517a1b6f4af8cfbd774bd1ea9409d47c5522;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23f419d7386238750e719a15acc4f4a41e5c7eeb00f81736758f5e9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea49d7e2901a8fdd572b513a0998a15e29851c81a2ed486c7b92f526;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h140700c6a26117eb0c6b3bfaa48ff26292af14ac283bb45af7d456c10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3562b860509e52943337784f872935e5f209eda9d81fede151cc1d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d5f7f6ba61285c736e1f96fad97c06b8363ace1d366ffed27968a92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92890251ad0bec3cf65c2d68bdb6d785a2e82a8f3857e7fdaa66f9c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fddbb6d7b580ec96a56107e064a22f68155058c00dbf94cb57fad268;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb624663238173e6b5651692de5d1c27af82a4be6a4f62f80158e724;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd2c5331944172a6a7b65e940a07e07c04173ebe6a164ad8f817d65e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c4d66fc586bb83392f675b442f6bdb166d57d41e0780f905479fcf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a9667a6f33ccadaf9ef60f3c663c27440767905dc2f5d26fa6a6806c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e08a13252a6056195681f23a284dc620b2c278df3ca26d94cda9378a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd3ae9b831f682f6fb81a4fc4885d6e8516a3a0aa8df09339e1b8e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9e978d67b7e9d3e503ceb6fc147245fd11f539fc97679d9083d6506;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf1f7b731f2886ef8054239448a5e60e5bb4b04ddc574f66a1cc92a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb21f586ae49b04100995761d5fdd64de920a4a892494ece4a1aadd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf47a76284317c63cf5372f5d130adc78ca7b270bacc28651807a42f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1656bdc9599bed230462f7ab10f259a1a071de61cbcfc87687e4dc370;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc3835f11d168a8260f5a97d04c5f00e50c79382680cac207a398eea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c10c239c73094ad426594fad8fdf1d1108b18a7f22412b7732d78d43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19eb04b41d0a2b77d3d6128b990b594438aa9d708e6b709d3784073da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb6369243809a0742e29ec6890ce1de241f6a4f61fee7568387402a43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119e4331f8d476e7fca90eb594b5d9cf80b6893b5afc9d58a3c7ce243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70b27c057b086735c59ecca6c4a0421944bb1a69124e501939d6f037;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd62b94924a001865e0004a36ba1b942e5ce5a6377ff205d023c61b49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a499b62d0ea442779b69bcc42dc2b93427d81ff5cbe439d95bbe208d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h881c2c6682f77c49587935a0f7b063a4ea1a42d686a544b76057fdbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9339f33c3f3360400906a224b95545c3730e0c1d4abe4973658f1d47;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he03f4977ccc9e6bb6ad8000c41ac705e830804f2d9687f53117f735d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53fc1c9d6224641aa65299250d1d7105067c9da8727aeb66a19eda54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he127fb6cb297d3fe67a1fd7cddddc6566b1005d43b739b90e6737b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h450555a4ac14a4a463a8ae7a2085ec7737d5353e5405ae41987b8fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc2ce1746e5a7f0ae6fde71b242f5aa1d8b00efc7c0d71dc0d80e95e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55d5ff64f63400bd1e361939021740768dff8353aa9c8ace80433d05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b4ce1696fce4a8afd18757c703734a2d2dedbbc456699beb0e17a51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85b577a8db2da7ebc63173fe02a3b979ba20aaa62e72bb9048a753;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5853821a0b8fa2069e84a32793fa91efb655b4933f8f0bf8c65a792;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7f1127cdd6ddc57f5fb88ac193e591fe115c4e82bc34d942cc4abf6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82ea0108ff16e448485b3688b518ef712dfc93932d0a76a56ca2d792;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19583af0242a7a5ab5c5cd2ab48e4054a7e6c8768c7d714b659615e68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38bc177b9d1db20e3fd1f229976d91beebeea628fee4a07e9f82ceb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had87fd49c75adb6f9c77815f729382f5ed84fc0bd8516362514da16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha939ed709540159982716404e4260a1b59cc71c38a3d1ffb4feb5e7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11e64b6ca2de3e39ac0623ae97aa1e3c8c0ce4b74b72d23adda4a46a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e922163968239f8a8316596fc0b5b88de6d6d2beef482ff75b678f75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17560739ea181928fd1447be43bdd003db3f498d13c64386eeb286ec3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19608b40718fbd6aa0ddf2d269b04b104fbc463d2e5cccff98ebd2d27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf91874548d0af23d99befcbd9b9509bb6935ac67c99aa32e03ec7f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d1537e8d6df1a2243ec0ead0d97de86c67944ebff45cdf43f6432f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1de3275844db970f5097c428a90f81c42257eece9d4c541a3fde575d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha61ce0fb1d79b4ace60bc2bb4472a19b864d377cfd5ab63b404e9862;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6d614ec7e05296659f13099f7fc10c95315d3f077a0622f5912cff6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129aebe8ad272c83edcbe401fc34e6c7a91dbee1ebb569bcf6959ae9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164893f9c0f80c6436db350c8d67fb818ecfa3eaae1547834e103f938;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1012bea4d41581181153948297f5a73d5a8097cb3e94a526ca0ccb33d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5af3180e3662e1372b0859259631ab32dc5b6c4ecff146b5b5af8aef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf355cbed3e996b7cff28acbde9537059e75efeadfe04e7880f1cfe0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19300b9c9158eab06bde95be48636f0f9d33334b1bc69604a35ff98de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eda2be002ab80e70365fa9cacd7971f4d32216c5a75223c6d54e1fd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13454fcd0a353b24775919c35db2bbc2e2cb630111036d9f04a0cd9f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1065758d3c6e48aa4ac821f1eb5e52f381c5012d80b435efa446e2e15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2a45ae0403e3a165515b8f5fa040d0861693bde6336db62d05eb184;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14eb20f1359be1392b2fb1220821858049ec7e2e9758391f2c8e9b113;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he98cddf6e52f40cc006325d2d79c69c246ac54fdf757f7a0a0738195;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c0eafceacbd70b3ed130fa437705ebd3f54ab96abf3ce2ef6d19e8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59f502d5d84b2330365f56058bef13a513f0172b2a641b3582a796d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1030fc6da5c9a3e7c1494598b6b0ca83fda2e73f1d0bf7467810e802e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he0c1b95148802b43cb65d488fb77b9aa6ccf3b8b435de977a9690d6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad5c66d2b911c27eb7fcbd25cb3558b050069716fb57df340fd4481a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1920692134cf5b918bde3061316405bfc4126de7aece7fe991ccbe0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbdd7b761cfd02a4f4bc32ba2cae74e04163ee0f136b814cc5a02ef6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa7a3b48cf27728f00269b1df121b114ac141fa9dd1ae5e1dbb861b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23dda0e40dead49c874ebedae236d4d1714c6142928443c97ed3a426;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9c1fbca13a9c25bcab947719ecbf9a33e38aa119c88a433e5af0683;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c6dca879d0200cdd7cd07ceed36716c7eb40feb807413e7a6092aa0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1684f9fff2592aa8dae930f39f8001463f6f4b80a02b5f4999e90a9d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36b95a49c2473b8d471e3bedc9f2f28ed57a8e55c5413d4113d8646;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hecf4daaf04fa3fdc97c7006df8d712f4e79d37ffcffaf1acd6d169;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194078c6181371d1224fb0ec1684d8329a95f952230a487882e8ee933;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d36e35b8e4dd7a96e7d4c0286e609419d41e57ea2501a01852fd05a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h132fbe18003ee6a77691b502457f9a5db600865b7e04d38f9f4612152;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a822fc2bb01e4915ae144316a880ac7909a22acecf14414809a31a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haebb9fe37d6ac7fb19b30d5ee4327e4b9085d3fa059111b5bed39dc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aed5236e97c040675863169270c446591c63badf8e2ece31b6f873fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58cbf3d057d0533ce9dc2ccfed16a98191161174ef27b5592f1e6fcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163d96ee0a4da917985339c463047f0e1ff6c3a6934ec1e13c9cc29cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63d3ed06f06542dc72ae63f5aeca2f7f33c49e49a7b847eb4b64e147;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h145012ebba7ff9a47917527d2ee735c8e08752bf06dfb3ea839d2c842;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6b8e51e4f4b17cdcaa10b58dccd88dd576da10ca23a6e297467909e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d2a0bdf9eddc96057a6cc2c7f339dc5a13c00c03583d823f809d05f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18eb460e95d736adc36cc80ee71d7b89455184df48ec2672507810866;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cfbd95cfd8eadb215a1d511b202d3b420ec1ea76f90cd7b97ab9534a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37854b2463b84ef33ca1eae2c60dd569b8b68a8de321530bb46d6ced;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dad593caf2e71c41d51e700f4f52841d181e39fdd362cac14c34aa41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b155765ffa2baba8b108660c877735b70a2d72c7bdb91c8bfac1751;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b7d045e63572750ee21b8faa7a2423addda43bd19693f78d1950b1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4da99cbc432b8c87640123c0eba14449658dd50288426cb884abf30b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc596a2c1490868d2fc09b089cea9c09a7cde38b3383598d28f2f715;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfff47a87241cfed406bbb9e0c5179f2cec6d2263771a9cbdd8e00596;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c050d83d6673f232be4b153eb70970c7ff6895b1a689778d9ec7dc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df5bf5000d3e3057b9694cbc055343d77cefb99909ff0d13da1658d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c54e4eda9f4cdcc1b12c352a46547a430288cee402093a5c30c2b406;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d096a99c28d58eaa27437c09d115871bc299b0af082d7b987a969bc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133fe7fd66589b02c552ddbe3ea2c42c633ad2cfd9af65494f34e4302;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4397117d18f18a966db084f7a5c3336e62b09517c9a992893f82a36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7cd14ccb58996de69adbdbe0468b811463f84134b13a004ff2f06fdc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a17257d663df974f81a4af2e148728fcc8b3129cb3a381c34b59da0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1799a151b99827df488f63b9c8251fa0c6b4089199a7c9a3d0f0efb68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1836d0dbbe2fbbe9e37e3f50ade2e2d01a4dd3b319cfabab647cae43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0b12f79a886fc0d3905b4c2a2a28526fb35ce5d00bc1d0c0a379a43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1447e89b59a45979b1600ba0b5e8018423bf4a62fc4a71b97831debbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a63d1441d38fe409f2c4501c5a37a39d34c1a556f4c4dd57d397f2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164be7e01e1baaa1b44ab338e5add325233316e0a4d26a63a0479326;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haaf77f8d62f4eb0902e89e8865dfa41ac149df740055b6f015ab71fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f3caf4ab541cd75fed7625fa9e5f0777036e107e5d5efee1fce6be5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h140d5c816768fa687eb958b91f9b2913271c2fb58bff33778d359f0d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h42f47fa67e403ea8813faef97c2cdf20e090dcd795a7430317d909c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d8bdb1709e5a2516d19305706913b7e76f2c44dfcc40db9c5605f0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19b2c9885ae8cbe4c4cc2c9b1692c4a138552d007d3bacae91a9cb896;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h122762637037e354330d93c4d77eb13885b38bcf2c1043df105d3cf28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6e13ac88249651f52cd1b29cdb524f40a3c58b79068a044315b4d9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1615666eb7adadda63cae9d3b15f98549b30d8dbeac7b56123a674c68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14cb30b569cfe8c04ace449c56438792b8590cb0cd7e9801ec5b5a6b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h392d33f403e535d2e7a87ee3de7f7fe583e80d436f4e1c0460455ac6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a4ae4a37970e77ae35925b81f7476b4fdcdeb28b89361f63310d5e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e9be930eb19d2b1e9974892bb4f8aa475d539b5b566e2a17944e9f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1b8c8f81ac020aa5bd1076b287a758f2fa857b62ddb3e9385134f34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d298f2e33b350b1e4fd9eaadf4df51897246e3dff63e281e5d4cce0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he73f7d0761871bc9bc39b4216622be7ed9eddf2e7d25ccf6fe377757;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b34585c46e628e3ce605ff4929615382a2aa492d2f4ebb9837fb8b29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1efc278565524c5ae731b28cc2898b633afc2029b85ca7e8265f980df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h500c9389dbe74a2f0e5342c385a830864da9cd89cbda33386f90336e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf7d93e11eae46b8e832c4249dd0a0db7bb1024e5dd8dcedecb96080;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30526b4feebcdd2c5d622073b9cd5965cd3c47da3177837e651f7801;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h54deb7b6697d0ce33c290e927c58bdfb2a7bf3290518af2300fc4aaf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h89bace713088f570835d7a8cac90e100097aa4357f1cfc6c25827ced;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2416ebc1b250f95189c740aa5ead5e9cdd6733dc4d7d329c37cbb7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h154a88453eb1b5008922d4ae6399eff7c4abff1004b2851f4222bbcfd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a984d02c4dd61ac063cc7b15b234130c3f5c76d1c0879d1f3b90efd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d91e1e6cae9a9327131d871615ab82e40185ec4b9db21e833648409b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c2b9649c1affd2c13877fb505ae808fe2cfc5bf4c00a1a694ffb5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aaa037b8e711d369fc538de77d82f878d9850e6ee391a07fef7bd71a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a54bbc0e47e2cd36d0a760a5f64f035c2b33b8523e1441a3860a13b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1daea7b33556b205b99228fc514e6565fb575a4347c9de868db29b3bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1257c48270a41c9fabcd4d18ed42de5e80dcc9572ee4e2e0d650ae08e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21a5a6cfb48480c76a1f68b3a916753c2a76a2264dbba14301bde6b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be83bf3f9a542b381fd83146b9b06623f3046daabd51c7eb398c1e36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5b947a030dedf412ef9d011e599c60d63a67768343a1772c96ecde8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f8228e0591faee8cf9b2f0150c547f6977e275fc97f5b94e12e2cd00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f8105289b350af203f90ad6a86c92ac77cb230dd05c304f33eff929;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7daf1dfc92011664300d708470039eeffb6878c0a723f75efd7b91a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b7be41b4b066269ddbf17575e237167cd4ec838bcc4cd7836721a21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0f1445d9275c91fcb27114db280d00d8b06bdb3cfee02784ca6a125;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4333682423a1bc0d1d582ab04d70967b8a905e1ebc0b684ac084a00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h600c49eeef2bf97810f4030bc0db56edfc25a796e21f0a50b7a42905;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1164375915c1f46900d00e61fbcf19bf88a53a81a5bc623cfefc5f176;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdeb0a45eceac2bc057847fc9a5a14cf7bb927e2a198b961d86c2e9a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1e1b3e665ed77fbd9db13fbbd732c5bb24b5a838505acefc2ce15b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111c34d724bb70c097ecdbebfbf1e505fc91effdd19a6813038e73d30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c1f4500b89e4f6171adb0ab50d151d8bc525da438f0490ed00db24a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1005416f4b4e23e45ee18779ef97155876854bae2da773a5b6d26781a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56ecf5ce89d31d4898e9ccc8feac1a7cf2f223a536084cd24b2366d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45e07cb7c52a1eaa7fc06c2072c7d0db12c522f792b6a489ffecf3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1875e136e1c61ff80eb1a9fc620feeb49efc0ba6295fe8944edc629bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f22669943417f18b1220bb67ab4a3c706390c7a005efb168af5a4f71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117b27e8093de4cf116d177c9f3a8d5398c7f8758f3843bbfca97fd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6f6fc1b53238ac0547ed70ebf0e3310eb542775eafb945959c288b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e004233327fce63106429333e6583928387794bb1bce13e86a3cd8c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bdc8a2da783a8a3fe668af9d11154890edc84aad1505a1078cbb30c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82e330710384ab8d81b2510feabfc1c867045028885995f0478e3a46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd7e2350a675b983c9e56ce0ffd1e531051c0a1b2ebe4b0ef3a73fcd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee8620cf9e58a642534bbc24976e80ed3d970b62da4390a15b211eab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c43f81dd02b72c11cc595ed3db7e3ca646e0999aec13d524a0ccf53a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1919abd26d2217194d96e260fb0e5a9b474cbdfc70c84c9fac0b53f25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125592ba7f24fcefe404496560e11c53ccee923e9488ad03f5e569fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b85963c26eecd1d38a2c59f788eac23dfca99861f0ab4efb64ecb396;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb96eebeb163765aa6298307a31db90ce5d9731b089d09cbf2e93d945;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf62ba4b54a2cf702128cc828261db31dd18cfc05d63b03556229d3c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40f22d5b88220a3de507ce18807c64a183da071979fefd6870827cfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he81ed6510d1054bb4f88b8ea7f50ee8d227f7ebc4e8a6cf4c3f016d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14544989ea0951686a8022a9dd1ae80b87929e74ad6df0703143a111a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1896869649869eceb1c7a832c8f4136df1702e6aeca04c49a3827e427;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e587df39ab21d09e93929c314047358f61e6951b3f99a888eae1bbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b62e353e6c7eca383c6f53df774f3038452bc837f0f713d936378e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12938b62f886467b4461ab030e714d39475494c73564a6df59d8a1fb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1583a6a0ede0bc1596280a868d8ef4caa189c1ac413b23ac9e338e4ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113fedc12ed1a496b507a6781ae442871c5595845c5771090ed4f69e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7b9dfb04cef204ff6732bbf2c9b260745ece652fd04f5ced3bd6d98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec4099111d4bc15cbaa0fa4b09a755f7116a29ef698d0f3f21f746df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f98ea43b0071fe280a3f060387917856a3b2dd1be2fd2a33c3da44a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c20c32d45a14cddeb30054bc92a2c35f0a3476e26db91d1949b0c7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7aa766aec34e4dc8223d6776f80548800e9ba6154a53aea328d23f8d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h102b11b3de33854d2d54e1006d8de0fbfb0b4527e148690280277b295;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe0e9b143b680117ea3844cdb6d36a7bf74cf1a36149d3809d2f6ade;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63a558fbb82e07dbe5b2cd13b37512049469cf7a2ed0e0a85c73d3e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c41a02fdb35b01537ce0554b4ebce115598e0d08be7c62ae07c575d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11bce95705d1a0b1de82490f03c2f2b6014613ceafbe632b56ac1aa62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1037f0cafd2061e0c51db9de5b14e5fa4ce1763269d2a6850ac29d426;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136de35f570c5b5772dde27bf326a4cadb33bf47089867a28759d4428;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a60b75b1fc0f34df789885580f23f62646b86aaa665e91bec2a7b3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he45941a9f2ed511528cc1f7b9071ae1528ad3bb6aa702fdcf6d7ba7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169cc4e01a64e489e1220a0265e1344821e4c08e8bacee54a96e309b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14febca39f265af86fa0057bdd5392ae2555124e219c3ec174a33dab6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd818268cd74cdfd5ea0fd57f418daf09e061d28833836a079b8408e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc3dc458f38f93da62beb5ed0206c3f0573804959e94e13044df24f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48a9643daef8e6c4db20781c4c80c879f981c6e4820132afcf5b9407;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h776737ea0ef25d92cc6d3c3dcb976d9fa38cea76372e75880a429c86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d899f3683aeed4080b7d41bdf2d85ccf27bda55b982883914c61985e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13bea018b10ddf6472cc28a1b2526ffda690666409003a47769c8deca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df713b99c014b87b1f58ffa92b00af78c59e917f4001fed603c91730;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9b95af41400ef43b6b77e94352a4a69a7b3e59b2ded2fc0bfa9dca6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h966c340bc8e1773f22cda0de655e7b494ec416d39d93516a6d1db036;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b5a03bccd38eddbc279b21095f3dc806ad19bdc80e62d042d605827d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db7b5f67158b5362676e2bf522b7427611eb902f3c7deab0a7f3988f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13b80b1f1d808e064e3c32c2314ee7d1ab8769127be19a5dc14a46001;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f799b6ebb89100da96bd85c18a9f5d2dc7724b878f48e85883404e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18138a16dd4ce0161eefd8a58b0e1246e4826fa77d0af0bc61c49034b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h25d7db8dac1af2438a954724f155a6f8e874ead1aad98adb69135bac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdbfe90a49852bdadfe67f6541e04ab9c3f4d8812b97422b4d50d50b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb59bf0cd3b94fc54d6fc45e94eed5b3f098bb005de88ed9e864f5921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h673054637a6c9d17504dc72ef283ae3fcb997163d7e350645969c915;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d2645834430ae0f7a6e4cfce8b1aaf9e423f72861dc88358c047490;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h22fdd0faff096149d72d113f37cf967b8a9a31d1abadfd3b05eec168;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb7c6d9daf382dacb5bb0541aa646e1ecc6cb68deaffc7d330a86786;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5b6634416168550e68098f9438ab020ecda27b3bfbc653a63f8eddf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92dbe3a5747f7d752f2138fe3f1b19b4150149a056a0f18d8d882b97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ac96f8098076a47ea9c675d1b11b5159218b07a7db8940732e58a57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e4eb81025d6a01f2ccb85167d424230d2736dc4b50044d41bc5aec94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7cb46cd6f5a2776d5807b02e3d82ddc20046b046497ad39331c3ba1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habf972271dffce0e56bf20ed7aa48ee2d049bea6ca70f1e1a6787816;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7da29d5abe175058c1326042e002f8b0c108b56fbe27840f56f0f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14bb5cf288a7b80099bee9ead60df69d7072c06afebda387cc5164e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7af1971af7ac2e5046f27321b3b9bb0dc96fe94e55defe6d2a3cb1ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a9d300811eb1fa0060c3bb9e161d6e2d7ccf017d0cadfa0de13ce7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d819976ae130420ae7e7ea74af054fbe8be4a14667721df5c13aa2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11991e3ddbe8357589b0a77f82d1f12c46ba82ac578e10db530e435db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdbb9383aca3d059d91f90eb669e2ce8b423a672ed12c1288cc0bec8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c11d1800b4a1a1429f3521f5ddc1f16934f856dc9953502601c22ceb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a82bdfa2229387a8c002135ab87eb33db5ba9792e6d5cbfeb6431642;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3157818caaa6f8b45960bd9250f670701a0fa6b594ca72b536238d03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h812b22646e54f92a9bb1e0ec168400c7d1917262a370c85649d06cc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbfdbc045cd0bd820650ec69afaad7c908b0d05334665d9bb666b3b2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d084727f5ec793f2ee93d009011b098ee021323d0d187f44f87f657f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h399275b7fc0770bf5a338e8335714ed77a517c13e5a44c6f7e2fb34f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90de00d49d009281f2619a3f41504e4e883878b9949a2f107c472752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c2974f0c06a9e401c718e1cf085a3733f88e3e4d8118fe7e703d8df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1781849f77d99e2b4c3f7bb9fb1b433d9d3d16e87c9491379b9ab9217;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf6e71717428bb6edc8eadd3cace4bec4ef5832e81192d42f25535d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e70e703354c11f861d506a04a6e61a35bb77a818a4e50365ebe0094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1322ae1fb0e2eff1f9eac70bf4a7cd11171136a8ef8dcdd03378ce373;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h281d4d358203289ffd0b2598bbf69942af5a0e2094503bf74bdb7c03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a9ad42c3b722944f5b5855774c1f68c178f2fc8b2bd176d6a4f217;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d75219e91c6651b945da9317e4bd31674d20f8f12df4f7b9dcc2091;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c32a84eb17067b84dc72ed11d034dbc6bfa13dba4de58b815c409f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18155f316de9a61dabd2b41452cc34a70ce9dd9c8a9cd1e8a7d45bae0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eea832ca3c21e24504811617196f59f9c579c836ec62290e67f40a44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4e76722c6167ad64fcc18a7c1b17140315772625a477e5fd1f27f26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d2171f6569d42013bc744a14bfbc35566c72a7c11e73cf515c70e89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf509ff1c04b8f2ac1db7c81351d7fcb646c9bab2f44848dc4acd5c90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h461ba74e853156c6e49cd00806de951e1338358bde0e70bb2e84603a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fbf069bb713321163a3d0525feefb25e758928734bdae55fc902b96e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde80f961b8adce069266257435a835c9f66ae85f3bd4958d943e5c9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b3e7439d22644390ba9f9802961679babeb70dce69934c2a33a2b39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19940c01e496d9486be68dfbec6532cfb39c923fe93070b01748420a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13586ca613a9da5ab8a77b45c588b7b0d31edc815f4862808a5f0419c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193d684e6751463ac1cbca610333391e17820a393089b4a8f5054c8a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105f2488a4489bfbc33cd6b075af6f5c654ae96aa4da9cb1b63948d98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h161cc3a6b28f14fd78b5bac96af79387b62912183c54600e4372aba18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha398d0d8fe335775f68f0e66ace4f60efaab90cc00e7ef044ad31b6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1536c3d6f41574216b30b558ab7d24264180dae1e299e8036f96d6941;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e89fc1a0537742c8061684420070a63b6b765d869d32f926798c2be7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18200e5b00235eaae940ef8db4114e876219796e00329396a40fd4831;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14351e7c2a67dfa853bfa3e2d0896ad4154b6515ae1ae1356d18452ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heafcc31faea69c2f1346df5cbdd5608f74603e4890fc8905ee05880b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7cf651553b67fb4223b138aec6f2692fecbe4d409feadb098cea4a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45219ea124419f507376303fd1f7842b3f20c2fe2765076a277d47e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74b072ded3385543de23295dee6edc67ef0a11db02c966c4f987ca4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df15f29b7b26161ca20a32e032cc1f948c137f091a5eb35479ccae1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17068f94ea261863d3f03a708d852dc1ec08999201bea87c881a96bd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdd4c28ed75d162de2fe2417bbf6051b1d05fc0f6e69f53f18f143312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4b312f9718369554c54218396a320ece9e78352785e83e3b7b83e14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135558699024396aa5924fb57b6715c86f0da4b16d572261d66e00d00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ecb65b7efb1ee2411e2d5c712b02ba3f3e07b5c7293528ff2500ab9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb07b5bfd1e6bfee256e99a5f169d8916fe82d6730777efde6d7bdf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109fb7f73f4aa0813f2a96d7b9388458543aaa05ba672f7b69aad05d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc2f7bb5902afbc876d5c7dfd7df6f51ad0b7d8e958ee37149dea669;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169fab0c0e7c8d13c0b6c3a4952f629f9b035e5a5acd22a58527ae2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7851149bf69af8134389d48680f31d2cbfa2fd46e2b9855caaf6076;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f63809d5478c480406ee49e2085e43edb2f4b4f618546151da4e939;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h104393a325d16ff2964f4b2e6b34d3872eb5cb106969f063a90f458d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2c2aa9897c8b00eeea9f1b3a2fb78fcfe060fdfb70a7498b3526128;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h746025608ad19db05cffe75e93aa9985d022209242cc0c3b2a5bd301;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1284d41c4426cf3fc385e9031310308b51f65495b4444373281bf0075;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed4345a60cdda2d2520d200c1592b7783cea5045e4ca472acd4925ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he07a199c798500637d87a7ffe52bb2afc5b08764dc0a0b39895bedce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c34c64044e28d8d293519cc7f2b6ca80d52689de3b59fc8e1d0eb90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ca0288d6214ec2097b7121481223d0c8f455a60fbf7904079b636e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d569ffe99d912e7d2734b02d1a6e019b92aa5a36a84e4464e0bbb62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c5b77f3989b795c065fc114fc9fdf9c26e9587ccef767f3ad380097;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f23357ee68ab01b2396830553c09c6926aad5f2d8215e923f3a4f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfae6a72f93f007588cbf61077d095b50ec96eee89c404f5777d4386e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7cf60f67e2cf3dd4efa603accf6c809f076834a685c624e4fca790;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf6107ad901bced404bac06072c1d2977a4ab7a1b14084aff504500b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7ba8fdf3f6cddb6d9f73e0bb16b62f993d3e716f53e348ffa84f774;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52b373f36858bf16262b7f2d5ff795ed9651bd254514ab1076eed3c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d5e5ad60607816e0f54957dab2c84082a18003c7ec9c5da153e5257;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1965953164b9261fbed4696ba887afc3d4649a9f34e17a4d74012755d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1522f9d1e6b0390a619dbff32186458b5dd9fc9350d128d01fe655254;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12971e9b2fd43c04893b0f50cca48a66c6d430db815aa516b2e18a345;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1c39dff51ab8cc23cdfe170c490264973ed941b3b158d6dec3a7e8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc47cac065a4382da78a75850a62fc68445b2a87b7c40ec5be5e373;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c75265e7370cbbbf642756524d46e9d561f102c9544bd3ef3080d4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b0c869ab31cc05908242286c732ea3e48f6aa02528d8eaf1edddcd93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6abb927d765bc8b4109c337bee3e2ae61276a3880d051742dc93daf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda16d6a0bd94175f77251ed72c4dba5780990c4fdbbbd8fa77f6fad5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he2aefbee0e95bf22f076da104d1e25ffd03a0d66392f7ca64f7238ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1b1cedfc1cc8037ed20963adb98f11b0a15fdfc1636f0da290925af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f65eec10ba16a42635d5f224f345201848066b4e3f1ab3490f23691;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16439398c0a5a7518d3fdab7785315f9c633245b79f7cd709b1324c7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8b1f7a06044ea8d7880a71b45cc8f92d61bcfe24d26a09a11d30f02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e245969cc1eb20375a24fbf821c81e62592e884415d398899c166ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b372f37ad43cb956775a18052f2ce6a7efdea971086aa187656d9bda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7236f4b44c685a6714b14f0a1a3dabbad1db6fe60c718f859791c038;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f125f678fd5c7fe8f99a9f5210344e7db80d4fee796f138ea8d6995;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106e8f785c2a30f5e43009174aa394a8b2aecf028f66c69f0d7dabb94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1409e26d69ddea76fe4af38da9c47ff88e5def76c1417ec338593671a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb78b3846e8fe585eecbde4aff074dcc0891646199d6da50a82c66a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8006622d0a95a30b51ecd3417e379e54f9c2b1849f731c8abc49343c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e56db570233a250555b518b32cc99d162db6fcba6beb4aa559572781;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf9ddf3bc64cd3c30482f33304a7118b90e4492c5dd12ca3f8760df7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h144ccc9fd26e7a4e54fdd60eed7e547d3d1c152d7a3479cec6a5f4538;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34add4a8d5539e9cd5452141a5ed9580ad1bfca29360f8fe09a052fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h73298b29376d2954be5524d8df614dd961af5291250df6039a18367b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee16c763876421233527ac9337e97c941491f635875e17ecd420338d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h187dbea909ace3b7bf1e989a70169cab08f039870fc33df8fa8f3732;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1513a9bcabc11b107329b56db729d5ae7d3b8d3f7523599a36d4eacdb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e54ae1ace023fa21181d40266fe67e484ce16195facd4108f389b61;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he26f67eb79c7d7668df353e62ea12a47a8c858dbbe93c7d678dc80fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fed4eedec0a6033f0236959bd4f870c2548b7ba0f0fbafa5e6df69da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1641159e6c7f0132ce1818f04476d527f5f8720dd1e1ef98bd2500776;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164d5054079c9edfd117f197d56293b6cb9ebdef7806d7022b9babea6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4237522594f2820b8d89b004588237e1991984462b04f22f46946f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdcc690f6fa177221b5fb785e58c9489112f5ea71e458869facd9eccd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd77f669157176521f8b8395d42d7049f5c28850c2d30d6dacb66e75f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19cd74e3401ee438eb369221ee3e3ab56cbe594ba974196910ba4cb4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157f0501434ccd94847feeb591d6982f9d8d8072cad72681cc830d18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18ad03f7b59050d8dafe8f8b0c1d8c393e24317e4c85ad5b7fbe37266;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f736a2cefd1d684887df63095a845b1f0d01b2d74d1a081a579efa67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c386aaeb36d777f5e29aacde25497b27e00730fd2930b2908842700;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64779c15955bd0334b29093214b9a61f65a905f818b918f4390a593d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb41522090e4d0ebd9e81de58e092ab129193021d96ea4ebc5c9f4700;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc028b8cad33930f4c77f0dabee7d81f10dfc867e212091f21813104;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3bf9c04fa353c08810bc0b34f5d094cd467b6d00d2184ef83fde827c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7572d2ecec572ad8a108d7ea6b87f48a8bcee40bb243c7210e4697e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1922caff129142def8dbaab41f9a41908848fc5827549710890b7a907;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf649664432b5ae0770e1cb57ab6cc64c309c5460d90f5e72308bcb93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d190423ba0e8ff8b79d0fe38657348b525b8baea9ae4b7e2d2d3242;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b359c07e4852b91b802313fea21e0d14b26317320932a83b31cf22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f664c082994a27a5e0568c42f67d0bbff76c75774bb210ce1d47142;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1348ed1e57b4c7aac965a81c3a8b99c96faa087e1a7309bc3951ad2fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1519f633ddb500e2c0639c1e9c432ec8c761e653ae827205f56963f87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a119c9082d39c290dc6f5059c2df05743d215e6ca6993c80edcf5a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7585ef385c83ee9c1378c03fcba52e236bc1985c99360d55fb836e97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafbc8d74049c79534487f80fa4ea2c68cba7882a1c7b1bd13ec0d539;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9fd3312386e618c438ad1d8016b123f682e7f92b47f586c98f76470;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h960a8bfca13d3933ea4d54fa6b04219557ea0a23837e4fec9760a648;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2543339cd0df0370d2bd32220d17afaef1c0adb5b14c50eb3b228876;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd2e159b5b89d481ac3ba895557d080b1239f13d5d38d530ba2335ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f37032bfd60a351875b923f643b2e0e577277c1541c1821ec9e21b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb9cfbc57a17f08cf7404b5482200f706cc9cd249d567e2a0f233a7df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7140b20d1f8bba27abcb003681c9b882b3a750a2fdd7e51a277f754e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd4209d2ce9cf12a36d466f21ee662761e5d7e7e9f71abb25808b9936;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ac6f866eb24ac78b9f1846d6793b1b693358f8f6a7f6a1b4144f695;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b5076bfd64d1e10d3cd2fb16bd059a87182d4a78c57d2ee56251fbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a4314c1608321ffe6fbb3af069855177b2bed05eb8405a737e72d6eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h151d1ee6e53c6f4bf5c3ac5b2845a8238e2189d92f8d9b0f01096f029;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f3873b6835a917a428dd492d4302467466a206db15111dedd662827;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cfce7658bb99f91c778d2a4aaa5f50288b65fb3435695309df161ae4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd42cd1421ac0c08ab515ee592ec4201d8b0182438d5296e0dab2515c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h439239c920a299c4c49f675d47c7b5deba8af6796ac65be63528ed19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcce7d3ea75d8a83edc0408a800ccd862e9c7ca91090c7874f44c06f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78f0656d4ecee7910609223c98d597ddbf2dade67d40bf108e3e814c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8550d3b5e2ca832ae697075bb5f386d45c5ac1024d31c01e9150e190;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdb4de84636b2371a671621a6b3690edb61dfa5c965e1967f76bdc1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2a050173215b2e0f44a5ba281e381ec9b7c5f7539a392f282d79ccb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13287de95ccaf85061b28bc7770ab0f70a1a05b6ec400a6ec98aad356;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188a39b3c7f376f1f06de936351c2afc13dab98c66987392f226602b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb9cc8db343e372f5f78b4f8f5303321fe4abb17977e9e96482e5d710;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8684b4df4ad5e5801cc1c5025e1bca96077c0718ba70907cf75ad400;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80807aa54b1cf912632f6f133ce5e1e14db872c5583d0edbfabbd52f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1910236805a4a8d7710a4127fde4fcbcb102fee112ac3c7c36fefae95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17992771dade3d8bd684c22049cb0cfb0461763e36e355eafdf0d96d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h151cc05b7084776e54ed92cad0616337b9d394d4ad0fea8f4b4f0f466;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5b9a73a0e985f09070e31463e72b400c0b4a0b354314d6da63a327b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb188aed4063b8d58314f5937cf1f6931921d6d8f179446f774b62a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ae437d9b0601fdbf9d09e0d9828a514628607661369ae15dd0c048f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14aa349c8da6bd099e8604f317aef511a76521057f1329bdfeb54aea4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde95a5b41c0b10c8f3b8a4b6e7d1c2837dfc1c78f14539eff4a30266;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c371f67dc0d3cd1c900361575f83e151555b48b1398402762a26241;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65428c648c51204897cee6d0c862bae44a445c1583e8338f658df3e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4bea40c69f48047858fb6c8ee07f132bd5c0361f571bd02cf71e044;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcfc98ea019f2f0348a40f1682a24a063318d5a3b067ee6833e1e2e15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2fefacf44c54ceab3243c1bea07b2c6b684715a39b2d3437358af37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4735c9e705a0b67d0de0783f4628f3c21cc3b56c501f72f78f14f098;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd63add97058a4b9931808f8bf33824d393d73377a3bcf93a1652ede8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b419a5389600d24af250c34aa4c27ee46429ce9db69b9ab750fa5f54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4646ee32579f84dbec891399db6ec559b73e1e2de5550bf8a991c52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ee6320eadfc9f5f719c43329862687d7c74a26b8207d84f2b7513d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h679fe676a77c23e335060e989ffb791616936abf83276084b39d9be2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc90e156038bd76a835197e20c7c03dfbaa508b6c1c126d292ec100b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11484a95610b200d6973c11ca89c26ddc69f8c2a76a539838f690cde9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a259b3613d35627cb355c48194cd2c8f62dc032455fc4e4680c9d19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169f5f5ace6791fcb89563c5b1344cb57c15d92c35af816e854f65e7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb44ef563724ccbcb0fd71f7d2a9b1b64cfe5fbf7d255a3f56781b84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f23e07f483689c1a771d0666e5261abb7d718224a3e85d21bb3ee0e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2bfd2e257fb96422144b14ce2ab692af04a1f78579d13e7d8047b01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f69bd8b206e9623293970e47c7650720b31d5b1a205cdb495bf0713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1868163533bf0ad0706d03ce432e6463ae993abc8b1616922967729c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7d0d40f7ccd9dc1c879e22108d82b38bbe68d96a3687fee3084b1eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129c0e42894c30cd843649181ee101a28b0d5af19e5775e6057688afd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1668be02f86e9ec714ddf0cdb8b6de2df23ff176ac68558bab29da409;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2421674806edf70d357887a3c2ec13f04dbf80f786e36e071c46344;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3995d8c78d6cb11a9fca759ca57b24169ff54ad853f8bef617eedd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f256afe80d7efd3a41c3d714213d819af63c93ccf570901d78433c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he2367cf8a83275adeaa113a407aea6f13cfd7e73d630761453612794;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c020f096a3c29d8e202b45eae80e4ffd35e72803a7b58737cdb1ae4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf8b9eb4ab8cb86b19114aa491b512128d31ecbd0a1e37803bcd61a37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6a087625978a6799bd6ae94273ce75a894e13334b1cb6ccb673721f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e19a0e669cb4d4203bf448fca19d6002a9dc2d5c3c356d4f92d86b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1161bae17eb0fa1ad2e02729839e13ed7ac2b89380f262179232f446f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h246fb41ba845d09be272d345de4cf27386ae42804cfee9c9d9f12302;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h73065960a3ebe134b8989f362eb95f992aabe4e46911984a1226efa1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f795019fc39e9ecbaab13fd911fe9fa6d59311c8c9bf8cecb308171;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcbb915b5376383764d183bc694be7638c1209a23d4f8a82e6abc855b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17dfd7324004f7b35cd5afe03b4a4649274374bff9eab973875f08b9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h132753c2a64c93dbd2f842fb1e68674c26987af438048b1dc99f7dafa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h552bc2dfd5227d86553f7d952c0147578eff0e0499c058438bce209;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf50c39ad02b629f861b5aba79ee2f23fdfc71462db6d24e356c6cc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b215e379e266edb849aeb534691087ff07008427d60896279805a9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15aef46fdc63f40811ab894a05819ab08b3fc2977a3740dd9a5a66263;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62421c83e3523961f8dd7a0b4f4747cda0bc79b7461634428af90c98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0482379d8221c683c6faaf225ee1f351df8ea7b5244a0caab03b017;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb34198f8f5cc75223709dca9622f5aae51639cba9ebc8e7be57b7f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e63a4c305d2637bcd7eb132cbfd34200a057e06874a0af6854b6d1a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h303bf8a3a5f49383c97c6156866d73d0cf1b12ce85bc07a765506dd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a374a23205ff37af480cd1edc985f5575e06f0c296290ccfcc370f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b1336a264d73cd88f322ebec57b98d57867b5c7f1cf955f28133095;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2410b7603fe6a38b6eebc1ed27db7c81a861958aa06372603a6c5025;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16fcff276b05c6c07e4c571fb954f0bd2e907c89261a9237e86d08d2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5c04bf93d955335e75083c70e3f92936073fc61c5cc1eb66545bab9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a83b0b578e307b960fc37267347da9904756491747c5fecd2566f852;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd85f0e051853c93e485a79d5d8d9b7146620e7f40a0ead1f9fbdcbd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93c53dec8a65a35caade2460b3f75ca838a865137e054488f7c634f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf362c64781fd19287b388d2cb13a31f74b74ef99a7b9b0a5acd9e66d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fa904e30f5f46751943dfcdc763b21ad72c1d5855b654f57eb0138e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3478556ad87e85ca6f9f9ad41c56be074eaf3b5feb7592b8232f49c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6276f88e05e3ad8d410c28523dc339521cb7f66df103009fbc77e8c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc209daa2365d0fadc6224e866b82979728da27c0772e00f846f8281;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6aa2172f27ac9020935537e78ffea2577ab21d5f8dc56798a87f31a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18624bf415431402bd88ef140e649db127a104a9947f43a0c6e2c30ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101ce11b733369a875fe8fe3870a4544f77aaf099e6fd325da6661feb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9bc64f48621e4f48166bfede927b1439c4ba7f8e78a7ede76f69cf37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195f4be896925d654da71809c431fd716c33dded69f8a23304a060fc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4c91d9a6db6edfcb773ad0a4352c77e4188fa264f8686494be6d8dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2c27221745654a31f4ec7b5fb5b6bbd17b131b63b0be234902b3d2f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101a6a5be68b3453d59d0b265c2255b3e8e9eb0481cedc684f2025c8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cce14fa91b52a4d27a2d13fa43fc54dbe363e877775d024269415bc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e1aa405386b1b9295d1d3b661166b1625f65c7c838dcd76f04c0d1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fb3dc7ad006031751a64b5fd183dd29cc2eedc5ea506a4644cf6f4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h162f59f23d1dc164c51931fd19f413bd8fc9407629c7a3a7f68a64a8d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d9c88ee0fc16cf98f6c991b839f48e89b0b32a92afec7d2f4f2e7dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h96796d2fe33a7276a7b348fb0589bbd2cdb19b0cde55165d26414c5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9f74137da4dc89ec4e0962594a98098320e0d1bc05f7afd0713594e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1200a06f7c0d2ac4a39c630323549c413c3501af4b581646ffcc3b422;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172188d86ee8cdd4ae70c8543e2e4ee56bc53d008a4e6772916f2dcff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1389c114cb263bd577ad3acfe142195c9892831d3b585b776fc9b81eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea3366f1664f0549018a50a4333e46abf46cc15ff1488b99e2a0a5b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h220fb39fda8314eaa3612211635484bfc109bd8e7e086c82611a08c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a5168efc387c490339b2af98322347f463963efc6de3e29addbbf49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103d43358630ee95b3c725eec40cb2b4b1732c3c34eb44ad2507bb6ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ff04aed2ef91a4723dbc473dd02f1a5afbafe19cb3417e43d1d1d0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc27cf5a6268fe03a4c0a4d6063c335b668bbf4c4ec9d2e35235963;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ae2f342c82f21a9899de48c7bef3f76bd5aeb71521f8131d29efcf5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c6a26394906c0970a9ebe8d117940c886d61bea47570f5cecd63df4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ccd43362b977bedc8d5ff8f92d9b018a26581d5fa42f09906fc2c7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc894a169d01751593e299fd9fb7b36564a26c4199a11a15977c319da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a70f6efc3697694eee832cb565c6083a61bbc33cf48b60e38711c583;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d9d2a9f32eead24bebb2f7bec7cf734df795f696f84f047049c1115;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h47bf1d014a248d2b5624adc72d5cc1e962dd369d28a090cbbb09dd0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86d92e915474547a50eacb6aa6ae5eb6e316928ad196f5ee8417fbd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1451753b9a477948c242b5017520865d62888155c7ead2faba19d16bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2da237c10363b193e8a40dc2389a0c0cde00e364cc6136b9ee47ea8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174d5fd7062c849042f858a08b5ff955f342fad7fbfe5736565a4ee91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecfc1d8c4bb1bf38fdd2742d39154c956b1df60c744a2a1d30614c41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f0bcd68b3f927bca8ce0646eb6e7635a73ea30e066558a747c19fdfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7bf120830ec2c8c0aff42a1a458630c74e57f3b67d1e37ae9efe8f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h786cac55644804e674dd1c08a3c257d86ae08809f41f2cd0c754c2b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e17a2b3e430813af581de385a033b0ee8a31ccb486534785b51f23f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51b280a48385b00fd1696ad6fc0ecf1989bb491fb529fa2ff0dfc4b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha756c7ec763500102ac81b68cee8db2432183d7f3b98d2ddc146a9e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3ee1dc49152a33ad5fe1b0ebeba953e40ff192715034aa89844ec231;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8363fb402b3308275ce496327b2538bd721d90c043b7e0ce9014714;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h31b38b4933528db77fac72255687a32b5c1dbcc1406e4157c170fde2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha556b6822e50e0aaf2337e830a58f7c1852c5686bf9e0f742b2a4a31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a64a43e9341abf83dc191473a8a890def8195725e99cfa3603ebc0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h727d74325f2ac093a96f028f2fe99242ebdba35bdb1cbdef9d4c6228;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h22e041470b8b552afbdbffb0992004ae9550383ebfdc6969ba219453;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113b79df9934bf601cc6088b46e996dd85037c76064481aacae21e904;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109618be3b405c1159fceafb364a01dd8a9db5e828172277dfeb017d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e79f7e0218e59c43d9842009e7d4b81649038865f0b8fcf732d9087;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e98952e1d4bd7f0c3c1c0e567b7278887b573b187a28d51e41be523;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h593e034e8393a017be0d0dfd130d4c4c507af002095a6025224c8cd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2d8072b21bae63c1bd07fd1e0b11135228bf72cdd875b1218f7cd2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c11142a24e8ba866454ccfdc9e472dfbe79dd60ddb843b2c14bf980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19233c17e456d6653554fe332b03561661407287b240e766d4ecadacd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5aa6a96fe820b7b36c43da18e8fc228ac46ca92beaf64557d6b232b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1416a3a321c00784d8cc0689744be2f940e0a903287251c6261b7b206;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f76f8733feceb1a7fd92165e489a64574eb928760c7804913c590623;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c9d88d417e4060b94eb085147a93ff5ac645747b590acd7ac56542a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ae6fc61dade00cef74ca16ac18146fd29adafa760b42210afcf337d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c3a505ca5a0a3d62266d4d7b3179f612779ddd53cc3a2a24bb7ae92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b0cf14a85519db7943f477b6aed76ce13fec5ac877a7f0c25d6fb94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1725e0b78106e91c44a5ef7462cc543faa5359d1b23ad874e2ec8e300;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28c54eeba92b1179a07405a98ca4d53ba6ea42b09f466b5bf99ce259;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3feac451d73aca578afdb47ce2ed69d1992ff90c98d437a15196e57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7a493c341ae75e432683bbeeb4dbdf7a66ef264bcd56b80aa3c4a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha11559358fd21598bdb5fab6e381ca1cb51db454fda564278d80bb35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c65dc5499cc0f16573162bc37edf77e40d435b73a6f875d758ec7d60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa3dcdcd124b925b1f3548b69a7b9d8b4205e2681849c0dbf9dede78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h161d29e9a0dbb856b3bad74e57d5e2981c402ba791e107762bb97e2e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aead159a98322dd54a3e44f308a56f54c27bf04daaf9166dc049a1df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h730e11686b3bedd6eae8b95fab36f336844d6b35bd481eab8608dc58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac1bfc40baa4cf19501c3307606d8a7b2c3c15aaa6c70db5e7af413e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c1f0be92e6f004ac5d5a0fcf74db906b0fe0ddb017ced569e54b6f4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f2177b013db54048ec1239d3066ff6eec374136f95ffada137ba5ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20a2e3fd7e9191806c94671fd216b5ed108f97b96ba33e31af4a2cc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1046880890b7981e682fa43efdbcffb28ae63e7b179dd3a333631f35d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7892397ee2eaa3d511b75264d95d9b9bac7e632bd99b43ada8a54b90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h425b23e6ac4f957cd5f629bd6662fdbc1c3545e834308db63e0de71b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1554bb03744d1b4340012931a53f2cafbab2856bc9f8032618b5b1ac0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee80a682e11674c188033dcd9579449eaa375e3a1ea17e13330fa725;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e57bd45da10a41b1a5afec25db31e681a2c2603e0aa26cfa74c2da9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51961279225778bd1beb0a184e51a31c7baffe6c4290a65fb2d91afb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b809312a7c87484e4a0b4351dff780d97680b3b99fca4eac44c7767;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18abca67afa9117a04000ae74f1a8e39bf44915086158b0d1c4b5bbf8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153c5ac31bc0e79fb5315ad3da1f415334b855bf080ed799a8163fd58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h821fde715c50b9942a62983279ef8f4325576c05ba0b9facaf0aba21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff20acb2ed409e2599bab0efe438d41bcd00c0b14974dcd5a24e1001;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc17899eddfbd8576d6f37ec24970aed11666056469e38cb1cb2e70ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6a5f636d7f5c70fc831edaf7691428857ad6d0b48100c82e6aecd60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b375c6761e54c68801de6ad5832ab208dc695e01a9ac312ffaf6b3c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7801e8c14157a83bd045537c352464abc2a630d99d72fe5696b83a4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1172788aee2f2cb78ec41afc42e070b59fd8bcc1479f2b17ff1556c23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c930c3d7a3ffa2b32054deca46e8d43634fe5c32226ca46d75e56cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f96861e9d39333b16d9d47b17af0232fbb01686821cbe53453e2efa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1103e507b11f51cbacee52b8d04dfd86e050c07057bdcb32ada5469c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha59bd2e39f3d6d7026918acb806b1260eda0e8d55b675f556ee6748a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66ab26cb0d13ce0775bc7e44b8b2efb9b8fdbf1de9dd8da6a74a798;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bfa6444078401955cae53a347fd67317d58266d5bd6e27032a82d94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h933a65d8e9af7746b8f84b7bb506627d36d3237c41b988e25b11f897;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf59b3802db73b6b7d0e77bb0f6b00f01e6ab7aef960b7f5483c70c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32a0108bffba36e26748c186fec697f1f66e6c74a5594074a110fa78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ca8c1ad0fd0cc8b52af8adbff32621ee2dcff2cb217391a88e6e5e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a88711deec2f9115cd81c0fbae76c09a0632e1d3d25cd06a289896f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142fd6d4094348fb2b846c155bd48e4b29900607e2e31e2d41fe7923c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1301fb01f61cb303e14697c7474dad884d27b128196b43c6ff8f2acd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h69bebf1a505252555ed01ae8c86b59f9102c882059caeb7a423fdbf7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f05836e9de1312be48dcaea3512f503bca5636049c701c48b95f7c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94cacb65e0f8a30c8a3438bc78bc17a4586150c1bfe50d0068257404;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4dc3315f77fe80e5f1f52e2c7db68dc490d994bac9e31b101c2e828b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11e4e303fbc7e34308f93c1fca5f83e64fa18bc1d986d9f2659a1b47b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h908b6511f1ad37df8f83570d739df586d0235b4b44e96c2eeeab869b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f18a6c2c0a3889ea955e94b7a4f9c41d1f1cc357d9f4dd67efcc962;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd45f4d03b0adc0a9da9e3f0a33971bbd551ca7694ab9aa4d78acf7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h182e0c49edad0930212cd77f61cf88139c06322ae20ea40d1d88e772a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba0e755a03de76dafe4b4bdba47e6c9d1fce72c062c9ed7f09f1b6b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbe7598f2868520b25f201faebb2be50251984b152e76dab521264fc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c22fcf2e48328a7ed8d5624a140e8949d3050c6beffe8a0cb3806014;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c76611c651c448ff3fd6d2cdc0172c2bedaeea724124d79fa16afce0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd7312b4eff5405a4efc8ad93aef1a700196d31dbbaa784a5ac639731;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c322721c20b631d83fc60d8dc8b8a04310d9bd3bbb66114f7034a14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b5b76c12a007bf590ed223a2f38af927cf95ccad55352be5754b37d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8e214860acd19cdad3445ec39ca87fda31e68edee9e23029910f7f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2067925110d42c7705bd04648ec3fee86c25ed8c532d817f2847b25f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4b629d883c8f7525ec226f88a3a5f64a8ff62cfc9b709f0d949d045;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7dc9a04eaf7658a028ddb8d733fef55adf5f6cd20f6a20c0b8f752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd2b7a4fece350ed30b2e65193d592b80b4fd79ff85701bdc96c7583;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h495caaf7ca8146ce762350c84d723a27c29229fd228db813c3a17ce1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfdc169e0a965a404d72bd4bc09bd2ac7d92ecc547bc596abd8dc6eaa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181a7652780aa20a5d59c0cf9d7ec46f11bda0cb236ede5db8dee60a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e7b36ffb7ad9acb305b214773a89eedd6ae8833adf7f6eb2c91cc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ed0565266f17e4c9854ab07a7531a85fd71e6bc241cc502cc6e9fd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb379502d9d26afef0fc6f3f26f6b678b563f9ba49f433b1f840874be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ba326a2579b56e7c1222d7a5cda3af6e60ac5b1fedf2a9eb44be794;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1621d10f9c535c5dc62c6fb312c2cf01b491b8dcaabaeb9d260268d6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2398e802b53e597f6a18b9033918c0171cf48d6546f42ba1ddd31d8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a58440cee5a4fc5d41f63dfb0d6104b6630930e488609b92050f65a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h668c01e422404858b38cadc52039d1c0dcbca8c99cb0e6003ebc9561;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5a5647ae34891c3eb14461f3c3be8923b91cd4c1e7d439760393580;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1002fd0de8a9f597d3795726398c76c49d581b1820286b7e0850d8599;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb0f8e07d28a69ebe4a30d2b3a39ea8603d557858df4399fb6ed5c7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd846877707db0988f9b01d072b938c1fb7b1eb10b78cb669dfa7460f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d3e98de71f37f8afd1e91d6b251307c978fa3bfc5c797a99d5affdc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1644139c1c550561002796986e0b318b406d794383e098aca742132b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd0bf2a83fc27b68fbe23157156f034964d28a1a8f7d24828e179dcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h89aa96c6ff1068d2d28d56aa365c45cc709dadd9b2954a6f57f65d54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6fba622314b165e3e0d4d1e2224f2dfe4ce7432836ce4a6c5748fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc1b3df20cd90861102524b513433e06ca4ebf643facf70692ee9841;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha22fc4d23404519dced316cade50b2198b50124b3ca73bac751f62fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6bc40090ebfd9d37836b13550d4e22d32556256584a351444a675be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha6b1d55526269a1bc667c2db662044f00a2b10548604f95f4ca4cd28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1611ea68466c0db3a040fd84f61ec21d34c9b4b15fe822a1d8f54171e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e6782cb3c5b4371cf26b2ced4c184dd43e472da71c2f33421dd89fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd352dc6bcd921a86a42f5f7a17a5eef81e0ecd83ccb1e6c3277731d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a5f52a78d4306488ee6786237448c43785a2b634b0fecf5e537bba6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf46f06555f4823d3d07a9005107689108932f969276a01f714271b3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a67e9a3f7d30d69fd03223c8524c5a6c36870480ec9e24f08780dbd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b4dcaf13ad3ada785527615f9e35b4ce18242f14bd380c3ab38f439;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129d99315e1b55e2895b64b7896d26c4d085ad2704c4085a483a4cb21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d7bea78b908a719f4106d77571cf20dbf827f0173c539a6775c1a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h655a75cfdcc8c94406a37bd1eb754361dd839a714c7b53bec43bf89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a9706999c072716d2721bc9cd356d22143711fd8eb66becc54eba7b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c71c72c03ca63cfe79db97a1acd3b163f8a32f3119992796dbbf3285;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70a9e963267872d0168e566d2334ab34c7225ffb8868cab05487c0b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h47879837e46b64095d5b36101f79f1c75402635b1eb477a89f3cc7c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157bb72bd90022d8a608ee5c47d3992528bc26ec980fb6f418c65a101;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b04434acc7b2332b12f7497c6ad4687a5a9f737be42ce649a232a607;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10d7d3fefd19a3726fddee53271182a84bad575bb6b83057de0fc75b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee6186247efdb86ffeac4ec5ff76e65b675ddc5a700e105d3ecedb19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3bc0b8a0b2ec251698298f769dec33ba22241d526f7ac2da91a194f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb244153dce1ca609fa05995c93245b4f52b7dc2d484eaaab5a483da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1235a78c133d97a7a04e888d97bb10dc593f199b11a97ace94c3c8d01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h960a8b12714347bb2ec96a2120453135a84aac91c7a868308c72c2b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8be0698270e162c301dfda311907a7f8a71d618025a7c6db95fbb162;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h67bf31e402dfff28256f47dcc97d20f11f888321966bacfa653ffd56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1649accfe14821ba7145e951b1424defc85569b381700356fd4d67f6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hebaced39ee2216bacc564c011da16c8a5fdffb8c79197f723065add0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5129e37bcf27289a5dd9772e26c89b3318af1aff8dc37b2ca4934855;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h22cf6759c43a8eb70029362cb5f3daff6c4fde7d6a248da1733f9082;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h825f4e6fecd910ebbdd2288b43baeb369e734c4b3557016517248c4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d4739198129b95d961e0e9dfe65f751175f40305bf1f8f3cdae5628;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h568fb516f065cb31e4b282f0b600509eb67e0eed577e7d3d855e7069;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf934b854f48cfde912b122e617073fc1b04a3d17415ef844577ab7f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ccb9bcea7591435bd0a195dc96fd86f5616311a6ae79513eeac417e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1d91bed08ba85f6a645607c108f3632df00717dd86c882ec2fa53de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he98bb80a68770dbbe15f49b4117ab2e964908737ad90e161a1cfc912;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f12d60c82e8e3c93398087d97e9379449db1da7636d392d8b90c7a3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f5d76741916d7b030c416354fbe5a94c29173f348ab6aafcfd08c3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17eacab6f548316c655ca3b9b6b04428985e16d12615d4e262e8921f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb73625484f8c59cd3e01fd121f6bd416e833cd1beaa7af257be71e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ce8df3809e19cbef1ffdbba118b3ec0cc94ee84d845e17c0e947fbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h539f0f373c1cdfceac80704d59774b3ee0feba1cfcaed005bfe58e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a2b60823faef6151c2641832bd977790dc289398c75552619689f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde5a7c85394a6cb87e04711ad902008e5b20d34be51eb134c8bab6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155ece30dafc54313f6ac081aab65550fdf824cfd6ffed9aa0b002a01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h834ae1de23a4095f4f2fcdaeb9a2b37b182d128ffad454ed039824f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129c2d2a0dae4ae97ba783936fd29e7678219ff68f9ddee9f4399fc97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb784e6ebc82e198ddf010e4d3c0e88468c59145fb89197dad6ef2af3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he51b5dc77435e5eef7a10b744d13f3b6f5250330b0f758fdf9cb001a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffb9263b37e165e81d65d41ea82eef595b9e47efcca3e3bc494ed3fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h629e3cb3f39faafd15c64f29b1455c3c3e6d6595fffe519ffe47f07c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18e6c18d7e912f5c560b6ab05229786c787739841f483b2bdd4d5dea1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1f998fe365fe56709e1cafa4b89e236441419e4ebff9e0f63de4081;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafe84a3ae592069677b1fa537b64c34955054a0ea2af98f88b26450d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b2f0da2ad50deeb69be2061e007cc91a781e4fe2d8934670c2100ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18af3d5ccd63c439c09dc2ddb4212daef8fc26caa7c8036aafaca9334;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a071aa792bc87fa816f289b7115c6ab95d274aa703c6277d14fa4d66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a87d38282122c832f4b1cf33a6c66bfced7f5e12b41067ae452aeb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h835158b40b895a3e57ce026c05c7931d592d0af217a2e373d20019fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1529fac3ab1d5092adbb7432184dd17486c272f07ac26ff1aac5884d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c691381d58d71938dc815ba50e6d1606e358ed995f1a747382c85ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15cdc06843f44c1c56ac831e05cac2273771c481c15f9d76c6e98f615;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd02f583210fea5d8e2342bc2504831102edaeb9aaa30d81dc2952c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49eddfa703428277e6c9c991ca08568d16e13cdf4156d101b0dfd226;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55e5ba5869c961d9a7a62de1b378789f3b32edb9b59a9f44c3371ce5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4c8a416bf0b0d50c533ad8be991811619cfc3bfa827dc546bd9a524;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf73508048ffbdea1b61981a0b2da0295c0af868167936f4ffb864ede;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc4265caa6a46b6be62ba9a598059cff019cb8727dfb2ac742fc3c04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10a0f23ddbe75d6421815e82e3ad56f533133b34904fb860fe1440203;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h84a857ed08e9c1fcd16468e465332ec344fcdebd3166c9e66911a411;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc896593ea43dc37d8ecfdf8d1aac6a41842100e2c2a7c948c5db659c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17126ece7c08f4bf18d2c6108f00979fbb3af4fd27675ab1b6fc11f40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fbbe2b9709757b2896c851d3025973aaacd64074df1dab9e0a4af9ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e3584597992aec7fea45fff48be6d6f177de22c4dc206cd4ca6e190;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haeb8a95151b31134188c2930bdfc09d87b37b63b378ed809455967ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2c0967e06feedcf4c2df6514524522ef33923e85d24ee61a94c3a29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h986dd2f34dbe5b73fc9926ca610e51a9171d2854f9288839b6144db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1508c8af0980320e68cb0af6c7e0896c97448db103e884f591b97c4d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6fdd655df25fda550f2cb4342506084c34ac83e024cf68a9d2b41281;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152cbae2ea1ca5af8c3ef2425a10b42fcf99736a47c7c522669177c67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0c7ed47937a12858e48444333cc2779cc49b3c20123c86696214c04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e51a62d1cbaadd2a94fd71c75f16cbdd217302df5096eb12a07efa5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd989e3948980ee06b65c4b458101760a687c0290948b325eb3737506;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fa1faccc39e87f730ed5145e346b96a30a0f8e17ea7f86ca65683a08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147637fb16df1ef91236948c7a7d781bd1a6000f3a363c9a3be4477bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd4cc2758e120b72a3451abd2fb9c3ead9a21f27f1fc6f8c85249d4ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbaf570af0a2cd49511cd1fc442508db08500c6789b882663773620c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cc5f9d8aefd3a77fcb84328bc8b800d180eb57965a1015ee60fa7b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c54d9bdced52246b6488dc0310afba26888b9d67fd23777893f5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f00c7b52f7d4cc1e412d43709c32fbeff887b87b5232c6169bc52d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2ebb519b1ca8832d236739bbe7b8540822bb8495caf683de0bda2d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h953599bc52fc32e83aea6ab97eee18d7d05bb6d69d4563f214c0c755;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ddccca442ec7fb4a2af16070a741826eb8ece902bcea8cf79c0ee9c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113d5704a92547af91f6ed577c61a76b3a5836338ed97eecfd5b647b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d67f428ef584ce196ab30e110a067ec4ddbf0ac52f1b32b7fc703ee9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a90df493949c2813a49e02e9668ab3cccb901a54b80e5010885471e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da5a5ed91e30d5cfb4a2a082d4ed5e29a63142e4e61f1f451298bc8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b06417dc85393ed5f95a3dc6529673a083193ac60176e0a32a1434a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef419eb1f45b953f300eb5b5929bbf1ed09116c534c1a41bb209e4dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188c2547ddadc335cc4dfa9c48168427d3ca81eb0a0ec5caa7be4d087;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a18570f67adfcd4bbce9dce8deb724d2eb156b182ed19a67be869281;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7821be1b4d6b6baf71d0b361abb6d842a4faa4a8f5be2530a3da961;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36fe511ebd0e6f8fda944a044348982e17540c4f3eabaddbc869a3f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80cc028335cdf0eb780f2e9f9b1b27237d0d4b7b10c0b3eaf9d49b09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h357b3e90e64fd1396266789874f32ad2b4ae1df666a298259b09b287;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha94a483711bc7db1be2469998effb75258cee29f3aed7635f41d588c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176da57a5d9fd72426605a0518df681f854314b71c2319bb62e2898f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5920cb8ea6d352573a75819bba4a3a6d06f04f9a791781cd36ae3de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2786746066412ed5b2c5d5066810eff440c561354cd4e42d20abafa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd33610878a39dd7a2359e7ea6a84e0a259fe4722e16177d6f8747f76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda66025d52693214292b0b7e4705ee412b72da194b0dc2f4af3c41ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f21ee8a7a68315a5a27d41d371ea5c425c3b53853cbf35c3fb9e0de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8f2ff3df4442a0d6efd94e8125f260405781ed30bf6be2ad2507e25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36ed6b60bb0c98ec31f0a03c12f233a57a981858455fbe1ca60063eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153a0a2975d66fb807a2ca0fd293129a8e6e89e215fc76976df1137b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff0700526f92f7c43d6cb334909f7293cb35a6dbcb15721822a71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf41e4df2ff4e889681082f8f40e68d34b3eb322d625b18aefb77c18a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f5d59eea8ca0a13889323fd01426400b863028c2929c243e22f5952;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2892f6ea1f795be23f431aa1db55b66cfee9eea7e63fdee9126b2f42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f65f3bc2aff0ad22075eb367ac406e69452094c3699e9e01c824a07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a3beb91c60f6ea56289ae608505b2db70252434005079f10f993228;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad1f742a5a013c8b080f8b2b2a52584226353a8c140634aa3e5bb134;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f9de2ab0d245b12a15d3919d010a80c7f56146a278e03a81794a95a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e357f1b97eb968e1bb5501395100b45526ae753bc66dab7eb5de9fe9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b098e58976378c9a5195670218b44ecefb2a34904aa7284d4ebceb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1614badce67f53204885a9498c90ac7c671d520d3d20cb8eb93ebac73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1041b36287c1ebfc5a66003169eb730758b256b58dd848457f19b0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1770294ae663a600c2b68fcd99fa18664b682a4d5b459db3f3bdd6b55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h178148466707e3dff1207a10d2867e3265663546fd199891bb30a0c2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c134ef0bc85d2f76084c0062bc56ac2f712cd0753a231f6bd5579636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ea1a50ba7cd5367715c95bebae2c57bbd408acd84e9489f73263ce8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18202dc473b5d220b25adcef6a1da9fd0daa64dc471c8ef54791df0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d2648b562e6f657104f7c74f1d4c08bef34573d3b14dcdb0bfc975d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1cf70463717b7cb092c48e8007e2b88361a4f2a663f2bd1296937aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdb7ce4ea3021d780459b0ae98139214132e38d08873caebec104b60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58694708003e247fe82d2d4be9e6961a6c0fc610e6eeed48f2d07ef7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f3dc3af0bf749853d80697dd11d02d9fb916516174d5562996ad9be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d17599a95801644a54bce0e5dbfd0578b586a01931b03b811f32088d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c052a9c5e7a5eac8f74a3376aad21ed28dbbcbc3ea23859e30bd412c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c2eca8f704d8a45ce0496f4b733941e3c7d9a05156908f04dee2776;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d448cc1b66b1ff5e744241ebd50711cda3e57daf6f431255228d432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1776edbc667146194fa475b49e24c1788e12c546d4f45d208f96e2e72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12356ebe4a810dadcb0cd5f4af7027c9fb092bb45e28582df1767e1fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he35c6993a509e06a6774a4f2c1a85b17413f6abf13f52222e651c1df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1199ca3593ed6c7a82aebd07323b72a7ca244d17b763c0f71f7da34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d22e08a849018e213a11c270198562b914290353bb643c371b6c9ecb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0bc37afb8a17afad0e41d68044bd318e3db2b52f3871a102f57e383;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h77a9a45f2b08b2b215e7583988e01f7290e72f36359d9da570d21c8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he14754546ecd9d0fe0adefcaa6f012e984a6a57e4e00fb44756ca6e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a6c85aef8fe99644655c8aee842d41c07abf723d13e579f4c2dfb16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1101fce0a7c5c859acff72b5c49a703a8357c0c2a5abae39bfcf0decc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20a49f43070b7e8cb576fc04f4c1396cbe9a85e0f2e612b433da1f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ea0bdf9ab3f5b8c73500575102418026966f05d0c16b0ba4ced4947;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2668a1c2e38928949c80bd06790544e22f5fb26205a5af5d2b3bb70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd8edbdaa58c6d0cfce21942961866d1158833dcde3c44a0e873f51f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1592c807efef6f8fa250a5c66956fc6d48f7c6aa885a6c1d4b48aeb0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d85e878fef302bf12e7089b2ec820bae691325d9c13edfa681d2fe0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b9d668c93b511fa985ea3d647641f6a2579c3523f07613eaef67156;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1e65cd895c4bcd1d273ced3ec52a88849b96c2cf57419bc5b53f984;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heca959562ec5104ed43d2487ee7cc37e65abca76ff6f1dc3c7ca01d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b9f7649e6773c84d653283ea26433eccf61ba5da7c3118177df5a57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb024eb80ad7c7e716dd9683746dac90f0efc84c90b33486bfeae38e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5c707ee4bf01ecc144a1ab8342992ee1670c49c9326b97cb6c10ad6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c73e6ce7324626e004df4667062a4dae8c32f74222cf025f8b4b38d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150d519558710836d2e4183bf22a2047edb2ee3365ac1ea0cd8e399d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a752dbf5386de94496776674cac02fca038e846d4f38741c5fa2592;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d01294d2ec6f3389b7992d26ec086dcbaa943bc8d228536d9f86309;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a29790e24bd9f0cc9ac60efad4b570c1476492320d318c151737240;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7cf5ef46250b15d638310228aa555b1a1f7f973f47cbc4695bd74479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108eb82d23f200161097750800b79660217a78cdd5b9adb995a78c892;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14960ea567ed4308542b8389ad7285eca83b4c82b39d1db65ed152cf1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb75281c429332de12e9eb44513115f152d804d905397420aa6276fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93d62bece1fe706d1c53df0a0a5c52c0075aa8343d0c0ff6cc6ad125;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79d3730dad5ca458d5901eb27db1d797f3ae4e20122e22a08de38743;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12122c2d94cde1aeb769b63e58efe5474b89c0fd6ee043097f23ed8c;
        #1
        $finish();
    end
endmodule
