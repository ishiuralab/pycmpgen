module compressor2_1_128_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, output [18:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    compressor2_1_128_12 compressor2_1_128_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
        src32 <= {src32[10:0], in_data32};
        src33 <= {src33[10:0], in_data33};
        src34 <= {src34[10:0], in_data34};
        src35 <= {src35[10:0], in_data35};
        src36 <= {src36[10:0], in_data36};
        src37 <= {src37[10:0], in_data37};
        src38 <= {src38[10:0], in_data38};
        src39 <= {src39[10:0], in_data39};
        src40 <= {src40[10:0], in_data40};
        src41 <= {src41[10:0], in_data41};
        src42 <= {src42[10:0], in_data42};
        src43 <= {src43[10:0], in_data43};
        src44 <= {src44[10:0], in_data44};
        src45 <= {src45[10:0], in_data45};
        src46 <= {src46[10:0], in_data46};
        src47 <= {src47[10:0], in_data47};
        src48 <= {src48[10:0], in_data48};
        src49 <= {src49[10:0], in_data49};
        src50 <= {src50[10:0], in_data50};
        src51 <= {src51[10:0], in_data51};
        src52 <= {src52[10:0], in_data52};
        src53 <= {src53[10:0], in_data53};
        src54 <= {src54[10:0], in_data54};
        src55 <= {src55[10:0], in_data55};
        src56 <= {src56[10:0], in_data56};
        src57 <= {src57[10:0], in_data57};
        src58 <= {src58[10:0], in_data58};
        src59 <= {src59[10:0], in_data59};
        src60 <= {src60[10:0], in_data60};
        src61 <= {src61[10:0], in_data61};
        src62 <= {src62[10:0], in_data62};
        src63 <= {src63[10:0], in_data63};
        src64 <= {src64[10:0], in_data64};
        src65 <= {src65[10:0], in_data65};
        src66 <= {src66[10:0], in_data66};
        src67 <= {src67[10:0], in_data67};
        src68 <= {src68[10:0], in_data68};
        src69 <= {src69[10:0], in_data69};
        src70 <= {src70[10:0], in_data70};
        src71 <= {src71[10:0], in_data71};
        src72 <= {src72[10:0], in_data72};
        src73 <= {src73[10:0], in_data73};
        src74 <= {src74[10:0], in_data74};
        src75 <= {src75[10:0], in_data75};
        src76 <= {src76[10:0], in_data76};
        src77 <= {src77[10:0], in_data77};
        src78 <= {src78[10:0], in_data78};
        src79 <= {src79[10:0], in_data79};
        src80 <= {src80[10:0], in_data80};
        src81 <= {src81[10:0], in_data81};
        src82 <= {src82[10:0], in_data82};
        src83 <= {src83[10:0], in_data83};
        src84 <= {src84[10:0], in_data84};
        src85 <= {src85[10:0], in_data85};
        src86 <= {src86[10:0], in_data86};
        src87 <= {src87[10:0], in_data87};
        src88 <= {src88[10:0], in_data88};
        src89 <= {src89[10:0], in_data89};
        src90 <= {src90[10:0], in_data90};
        src91 <= {src91[10:0], in_data91};
        src92 <= {src92[10:0], in_data92};
        src93 <= {src93[10:0], in_data93};
        src94 <= {src94[10:0], in_data94};
        src95 <= {src95[10:0], in_data95};
        src96 <= {src96[10:0], in_data96};
        src97 <= {src97[10:0], in_data97};
        src98 <= {src98[10:0], in_data98};
        src99 <= {src99[10:0], in_data99};
        src100 <= {src100[10:0], in_data100};
        src101 <= {src101[10:0], in_data101};
        src102 <= {src102[10:0], in_data102};
        src103 <= {src103[10:0], in_data103};
        src104 <= {src104[10:0], in_data104};
        src105 <= {src105[10:0], in_data105};
        src106 <= {src106[10:0], in_data106};
        src107 <= {src107[10:0], in_data107};
        src108 <= {src108[10:0], in_data108};
        src109 <= {src109[10:0], in_data109};
        src110 <= {src110[10:0], in_data110};
        src111 <= {src111[10:0], in_data111};
        src112 <= {src112[10:0], in_data112};
        src113 <= {src113[10:0], in_data113};
        src114 <= {src114[10:0], in_data114};
        src115 <= {src115[10:0], in_data115};
        src116 <= {src116[10:0], in_data116};
        src117 <= {src117[10:0], in_data117};
        src118 <= {src118[10:0], in_data118};
        src119 <= {src119[10:0], in_data119};
        src120 <= {src120[10:0], in_data120};
        src121 <= {src121[10:0], in_data121};
        src122 <= {src122[10:0], in_data122};
        src123 <= {src123[10:0], in_data123};
        src124 <= {src124[10:0], in_data124};
        src125 <= {src125[10:0], in_data125};
        src126 <= {src126[10:0], in_data126};
        src127 <= {src127[10:0], in_data127};
    end
endmodule

module compressor2_1_128_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    input [11:0]src32,
    input [11:0]src33,
    input [11:0]src34,
    input [11:0]src35,
    input [11:0]src36,
    input [11:0]src37,
    input [11:0]src38,
    input [11:0]src39,
    input [11:0]src40,
    input [11:0]src41,
    input [11:0]src42,
    input [11:0]src43,
    input [11:0]src44,
    input [11:0]src45,
    input [11:0]src46,
    input [11:0]src47,
    input [11:0]src48,
    input [11:0]src49,
    input [11:0]src50,
    input [11:0]src51,
    input [11:0]src52,
    input [11:0]src53,
    input [11:0]src54,
    input [11:0]src55,
    input [11:0]src56,
    input [11:0]src57,
    input [11:0]src58,
    input [11:0]src59,
    input [11:0]src60,
    input [11:0]src61,
    input [11:0]src62,
    input [11:0]src63,
    input [11:0]src64,
    input [11:0]src65,
    input [11:0]src66,
    input [11:0]src67,
    input [11:0]src68,
    input [11:0]src69,
    input [11:0]src70,
    input [11:0]src71,
    input [11:0]src72,
    input [11:0]src73,
    input [11:0]src74,
    input [11:0]src75,
    input [11:0]src76,
    input [11:0]src77,
    input [11:0]src78,
    input [11:0]src79,
    input [11:0]src80,
    input [11:0]src81,
    input [11:0]src82,
    input [11:0]src83,
    input [11:0]src84,
    input [11:0]src85,
    input [11:0]src86,
    input [11:0]src87,
    input [11:0]src88,
    input [11:0]src89,
    input [11:0]src90,
    input [11:0]src91,
    input [11:0]src92,
    input [11:0]src93,
    input [11:0]src94,
    input [11:0]src95,
    input [11:0]src96,
    input [11:0]src97,
    input [11:0]src98,
    input [11:0]src99,
    input [11:0]src100,
    input [11:0]src101,
    input [11:0]src102,
    input [11:0]src103,
    input [11:0]src104,
    input [11:0]src105,
    input [11:0]src106,
    input [11:0]src107,
    input [11:0]src108,
    input [11:0]src109,
    input [11:0]src110,
    input [11:0]src111,
    input [11:0]src112,
    input [11:0]src113,
    input [11:0]src114,
    input [11:0]src115,
    input [11:0]src116,
    input [11:0]src117,
    input [11:0]src118,
    input [11:0]src119,
    input [11:0]src120,
    input [11:0]src121,
    input [11:0]src122,
    input [11:0]src123,
    input [11:0]src124,
    input [11:0]src125,
    input [11:0]src126,
    input [11:0]src127,
    output [18:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    wire [1:0] comp_out18;
    wire [19:0] out;
    compressor compressor_inst(
        .src0({src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    rowadder2_1_19 rowadder2_1inst(
        .src0({comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out18[1], 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[18:0];
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17,
      output wire [1:0] dst18);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [23:0] stage1_0;
   wire [40:0] stage1_1;
   wire [41:0] stage1_2;
   wire [57:0] stage1_3;
   wire [63:0] stage1_4;
   wire [61:0] stage1_5;
   wire [44:0] stage1_6;
   wire [43:0] stage1_7;
   wire [62:0] stage1_8;
   wire [63:0] stage1_9;
   wire [42:0] stage1_10;
   wire [43:0] stage1_11;
   wire [41:0] stage1_12;
   wire [20:0] stage1_13;
   wire [11:0] stage2_0;
   wire [8:0] stage2_1;
   wire [13:0] stage2_2;
   wire [20:0] stage2_3;
   wire [25:0] stage2_4;
   wire [22:0] stage2_5;
   wire [27:0] stage2_6;
   wire [21:0] stage2_7;
   wire [26:0] stage2_8;
   wire [24:0] stage2_9;
   wire [23:0] stage2_10;
   wire [19:0] stage2_11;
   wire [16:0] stage2_12;
   wire [15:0] stage2_13;
   wire [8:0] stage2_14;
   wire [3:0] stage2_15;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [5:0] stage3_2;
   wire [5:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [8:0] stage3_6;
   wire [11:0] stage3_7;
   wire [10:0] stage3_8;
   wire [7:0] stage3_9;
   wire [11:0] stage3_10;
   wire [10:0] stage3_11;
   wire [7:0] stage3_12;
   wire [5:0] stage3_13;
   wire [8:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [0:0] stage4_1;
   wire [6:0] stage4_2;
   wire [0:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [2:0] stage4_7;
   wire [5:0] stage4_8;
   wire [4:0] stage4_9;
   wire [2:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;
   wire [0:0] stage4_18;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [1:0] stage5_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[18]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[19]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_3[111]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[18],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc606_5 gpc42 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[19],stage1_4[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[20],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[21],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[22],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[5],stage1_5[23],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[6],stage1_5[24],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[7],stage1_5[25],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[8],stage1_5[26],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[9],stage1_5[27],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[10],stage1_5[28],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[11],stage1_5[29],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[12],stage1_5[30],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[13],stage1_5[31],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[14],stage1_5[32],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[15],stage1_5[33],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[16],stage1_5[34],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[17],stage1_5[35],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[18],stage1_5[36],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[19],stage1_5[37],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[20],stage1_5[38],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[20],stage1_7[20],stage1_6[21],stage1_5[39]}
   );
   gpc606_5 gpc63 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[21],stage1_7[21],stage1_6[22],stage1_5[40]}
   );
   gpc606_5 gpc64 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[22],stage1_7[22],stage1_6[23],stage1_5[41]}
   );
   gpc606_5 gpc65 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[23],stage1_7[23],stage1_6[24],stage1_5[42]}
   );
   gpc606_5 gpc66 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[24],stage1_7[24],stage1_6[25],stage1_5[43]}
   );
   gpc606_5 gpc67 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[25],stage1_7[25],stage1_6[26],stage1_5[44]}
   );
   gpc606_5 gpc68 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[26],stage1_7[26],stage1_6[27],stage1_5[45]}
   );
   gpc606_5 gpc69 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[27],stage1_7[27],stage1_6[28],stage1_5[46]}
   );
   gpc606_5 gpc70 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[28],stage1_7[28],stage1_6[29],stage1_5[47]}
   );
   gpc606_5 gpc71 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[29],stage1_7[29],stage1_6[30],stage1_5[48]}
   );
   gpc606_5 gpc72 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[30],stage1_7[30],stage1_6[31],stage1_5[49]}
   );
   gpc606_5 gpc73 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[31],stage1_7[31],stage1_6[32],stage1_5[50]}
   );
   gpc606_5 gpc74 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[32],stage1_7[32],stage1_6[33],stage1_5[51]}
   );
   gpc606_5 gpc75 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[33],stage1_7[33],stage1_6[34],stage1_5[52]}
   );
   gpc606_5 gpc76 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[34],stage1_7[34],stage1_6[35],stage1_5[53]}
   );
   gpc606_5 gpc77 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[35],stage1_7[35],stage1_6[36],stage1_5[54]}
   );
   gpc606_5 gpc78 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[36],stage1_7[36],stage1_6[37],stage1_5[55]}
   );
   gpc606_5 gpc79 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[37],stage1_7[37],stage1_6[38],stage1_5[56]}
   );
   gpc606_5 gpc80 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[38],stage1_7[38],stage1_6[39],stage1_5[57]}
   );
   gpc606_5 gpc81 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[39],stage1_7[39],stage1_6[40],stage1_5[58]}
   );
   gpc606_5 gpc82 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[40],stage1_7[40],stage1_6[41],stage1_5[59]}
   );
   gpc606_5 gpc83 (
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[21],stage1_8[41],stage1_7[41],stage1_6[42]}
   );
   gpc606_5 gpc84 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[22],stage1_8[42]}
   );
   gpc606_5 gpc85 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[23],stage1_8[43]}
   );
   gpc606_5 gpc86 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[24],stage1_8[44]}
   );
   gpc606_5 gpc87 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[25],stage1_8[45]}
   );
   gpc606_5 gpc88 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[5],stage1_9[26],stage1_8[46]}
   );
   gpc606_5 gpc89 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[6],stage1_9[27],stage1_8[47]}
   );
   gpc606_5 gpc90 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[7],stage1_9[28],stage1_8[48]}
   );
   gpc606_5 gpc91 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[8],stage1_9[29],stage1_8[49]}
   );
   gpc606_5 gpc92 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[9],stage1_9[30],stage1_8[50]}
   );
   gpc606_5 gpc93 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[10],stage1_9[31],stage1_8[51]}
   );
   gpc606_5 gpc94 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[11],stage1_9[32],stage1_8[52]}
   );
   gpc606_5 gpc95 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[12],stage1_9[33],stage1_8[53]}
   );
   gpc606_5 gpc96 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[13],stage1_9[34],stage1_8[54]}
   );
   gpc606_5 gpc97 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[14],stage1_9[35],stage1_8[55]}
   );
   gpc606_5 gpc98 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[15],stage1_9[36],stage1_8[56]}
   );
   gpc606_5 gpc99 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[16],stage1_9[37],stage1_8[57]}
   );
   gpc606_5 gpc100 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[17],stage1_9[38],stage1_8[58]}
   );
   gpc615_5 gpc101 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_9[0]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[18],stage1_9[39],stage1_8[59]}
   );
   gpc615_5 gpc102 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_9[1]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[19],stage1_9[40],stage1_8[60]}
   );
   gpc615_5 gpc103 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[2]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[20],stage1_9[41],stage1_8[61]}
   );
   gpc615_5 gpc104 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[3]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[21],stage1_9[42],stage1_8[62]}
   );
   gpc606_5 gpc105 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[22],stage1_9[43]}
   );
   gpc606_5 gpc106 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[23],stage1_9[44]}
   );
   gpc606_5 gpc107 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[24],stage1_9[45]}
   );
   gpc606_5 gpc108 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[25],stage1_9[46]}
   );
   gpc606_5 gpc109 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[26],stage1_9[47]}
   );
   gpc606_5 gpc110 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[27],stage1_9[48]}
   );
   gpc606_5 gpc111 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[28],stage1_9[49]}
   );
   gpc606_5 gpc112 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[29],stage1_9[50]}
   );
   gpc606_5 gpc113 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[30],stage1_9[51]}
   );
   gpc606_5 gpc114 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[31],stage1_9[52]}
   );
   gpc606_5 gpc115 (
      {stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[32],stage1_9[53]}
   );
   gpc606_5 gpc116 (
      {stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[33],stage1_9[54]}
   );
   gpc606_5 gpc117 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[34],stage1_9[55]}
   );
   gpc606_5 gpc118 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[35],stage1_9[56]}
   );
   gpc606_5 gpc119 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[36],stage1_9[57]}
   );
   gpc606_5 gpc120 (
      {stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[37],stage1_9[58]}
   );
   gpc606_5 gpc121 (
      {stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[38],stage1_9[59]}
   );
   gpc606_5 gpc122 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[39],stage1_9[60]}
   );
   gpc606_5 gpc123 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[40],stage1_9[61]}
   );
   gpc615_5 gpc124 (
      {stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_10[126]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[41],stage1_9[62]}
   );
   gpc615_5 gpc125 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_10[127]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[42],stage1_9[63]}
   );
   gpc1_1 gpc126 (
      {stage0_0[127]},
      {stage1_0[23]}
   );
   gpc1_1 gpc127 (
      {stage0_3[112]},
      {stage1_3[42]}
   );
   gpc1_1 gpc128 (
      {stage0_3[113]},
      {stage1_3[43]}
   );
   gpc1_1 gpc129 (
      {stage0_3[114]},
      {stage1_3[44]}
   );
   gpc1_1 gpc130 (
      {stage0_3[115]},
      {stage1_3[45]}
   );
   gpc1_1 gpc131 (
      {stage0_3[116]},
      {stage1_3[46]}
   );
   gpc1_1 gpc132 (
      {stage0_3[117]},
      {stage1_3[47]}
   );
   gpc1_1 gpc133 (
      {stage0_3[118]},
      {stage1_3[48]}
   );
   gpc1_1 gpc134 (
      {stage0_3[119]},
      {stage1_3[49]}
   );
   gpc1_1 gpc135 (
      {stage0_3[120]},
      {stage1_3[50]}
   );
   gpc1_1 gpc136 (
      {stage0_3[121]},
      {stage1_3[51]}
   );
   gpc1_1 gpc137 (
      {stage0_3[122]},
      {stage1_3[52]}
   );
   gpc1_1 gpc138 (
      {stage0_3[123]},
      {stage1_3[53]}
   );
   gpc1_1 gpc139 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc140 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc141 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc142 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc143 (
      {stage0_4[126]},
      {stage1_4[62]}
   );
   gpc1_1 gpc144 (
      {stage0_4[127]},
      {stage1_4[63]}
   );
   gpc1_1 gpc145 (
      {stage0_5[126]},
      {stage1_5[60]}
   );
   gpc1_1 gpc146 (
      {stage0_5[127]},
      {stage1_5[61]}
   );
   gpc1_1 gpc147 (
      {stage0_6[126]},
      {stage1_6[43]}
   );
   gpc1_1 gpc148 (
      {stage0_6[127]},
      {stage1_6[44]}
   );
   gpc1_1 gpc149 (
      {stage0_7[126]},
      {stage1_7[42]}
   );
   gpc1_1 gpc150 (
      {stage0_7[127]},
      {stage1_7[43]}
   );
   gpc1_1 gpc151 (
      {stage0_11[126]},
      {stage1_11[42]}
   );
   gpc1_1 gpc152 (
      {stage0_11[127]},
      {stage1_11[43]}
   );
   gpc2135_5 gpc153 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc154 (
      {stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[1]},
      {stage1_3[2]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc155 (
      {stage1_0[8], stage1_0[9], stage1_0[10]},
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_2[2]},
      {stage1_3[3]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc156 (
      {stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_2[3]},
      {stage1_3[4]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc157 (
      {stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_2[4]},
      {stage1_3[5]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc158 (
      {stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31], stage1_1[32]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc159 (
      {stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37], stage1_1[38]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc160 (
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc161 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc162 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage1_3[18]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc163 (
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage1_3[19]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc164 (
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage1_3[20]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc165 (
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage1_3[21]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc166 (
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_3[22]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc167 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[9],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc168 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[10],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc169 (
      {stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc170 (
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc171 (
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc172 (
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc173 (
      {stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc606_5 gpc174 (
      {stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[7],stage2_6[14],stage2_5[16],stage2_4[21]}
   );
   gpc606_5 gpc175 (
      {stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[8],stage2_6[15],stage2_5[17],stage2_4[22]}
   );
   gpc606_5 gpc176 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[9],stage2_6[16],stage2_5[18]}
   );
   gpc606_5 gpc177 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[3],stage2_7[10],stage2_6[17],stage2_5[19]}
   );
   gpc606_5 gpc178 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[4],stage2_7[11],stage2_6[18],stage2_5[20]}
   );
   gpc615_5 gpc179 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[5],stage2_7[12],stage2_6[19]}
   );
   gpc615_5 gpc180 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[6],stage2_7[13],stage2_6[20]}
   );
   gpc615_5 gpc181 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[7],stage2_7[14],stage2_6[21]}
   );
   gpc615_5 gpc182 (
      {stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[8],stage2_7[15],stage2_6[22]}
   );
   gpc615_5 gpc183 (
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage1_7[22]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[7],stage2_8[9],stage2_7[16],stage2_6[23]}
   );
   gpc615_5 gpc184 (
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_7[23]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[8],stage2_8[10],stage2_7[17],stage2_6[24]}
   );
   gpc615_5 gpc185 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[9],stage2_8[11],stage2_7[18]}
   );
   gpc615_5 gpc186 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[10],stage2_8[12],stage2_7[19]}
   );
   gpc615_5 gpc187 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[11],stage2_8[13],stage2_7[20]}
   );
   gpc615_5 gpc188 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[12],stage2_8[14],stage2_7[21]}
   );
   gpc1163_5 gpc189 (
      {stage1_8[40], stage1_8[41], stage1_8[42]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[4],stage2_10[10],stage2_9[13],stage2_8[15]}
   );
   gpc606_5 gpc190 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[5],stage2_10[11],stage2_9[14],stage2_8[16]}
   );
   gpc615_5 gpc191 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_9[30]},
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage2_12[2],stage2_11[6],stage2_10[12],stage2_9[15],stage2_8[17]}
   );
   gpc2135_5 gpc192 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[1]},
      {stage1_12[0], stage1_12[1]},
      {stage2_13[0],stage2_12[3],stage2_11[7],stage2_10[13],stage2_9[16]}
   );
   gpc606_5 gpc193 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7]},
      {stage2_13[1],stage2_12[4],stage2_11[8],stage2_10[14],stage2_9[17]}
   );
   gpc606_5 gpc194 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage2_13[2],stage2_12[5],stage2_11[9],stage2_10[15],stage2_9[18]}
   );
   gpc606_5 gpc195 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage2_13[3],stage2_12[6],stage2_11[10],stage2_10[16],stage2_9[19]}
   );
   gpc606_5 gpc196 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25]},
      {stage2_13[4],stage2_12[7],stage2_11[11],stage2_10[17],stage2_9[20]}
   );
   gpc606_5 gpc197 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21]},
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage2_14[0],stage2_13[5],stage2_12[8],stage2_11[12],stage2_10[18]}
   );
   gpc615_5 gpc198 (
      {stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26]},
      {stage1_11[26]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage2_14[1],stage2_13[6],stage2_12[9],stage2_11[13],stage2_10[19]}
   );
   gpc615_5 gpc199 (
      {stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage1_11[27]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage2_14[2],stage2_13[7],stage2_12[10],stage2_11[14],stage2_10[20]}
   );
   gpc615_5 gpc200 (
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[28]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[3],stage2_13[8],stage2_12[11],stage2_11[15],stage2_10[21]}
   );
   gpc615_5 gpc201 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_11[29]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[4],stage2_13[9],stage2_12[12],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc202 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[32]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[10],stage2_12[13],stage2_11[17]}
   );
   gpc615_5 gpc203 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[33]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[11],stage2_12[14],stage2_11[18]}
   );
   gpc615_5 gpc204 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], 1'b0},
      {stage1_12[34]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[12],stage2_12[15],stage2_11[19]}
   );
   gpc117_4 gpc205 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[18]},
      {1'b0},
      {stage2_15[3],stage2_14[8],stage2_13[13],stage2_12[16]}
   );
   gpc1_1 gpc206 (
      {stage1_0[17]},
      {stage2_0[5]}
   );
   gpc1_1 gpc207 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc208 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc209 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc210 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc211 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc212 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc213 (
      {stage1_1[39]},
      {stage2_1[7]}
   );
   gpc1_1 gpc214 (
      {stage1_1[40]},
      {stage2_1[8]}
   );
   gpc1_1 gpc215 (
      {stage1_4[61]},
      {stage2_4[23]}
   );
   gpc1_1 gpc216 (
      {stage1_4[62]},
      {stage2_4[24]}
   );
   gpc1_1 gpc217 (
      {stage1_4[63]},
      {stage2_4[25]}
   );
   gpc1_1 gpc218 (
      {stage1_5[60]},
      {stage2_5[21]}
   );
   gpc1_1 gpc219 (
      {stage1_5[61]},
      {stage2_5[22]}
   );
   gpc1_1 gpc220 (
      {stage1_6[42]},
      {stage2_6[25]}
   );
   gpc1_1 gpc221 (
      {stage1_6[43]},
      {stage2_6[26]}
   );
   gpc1_1 gpc222 (
      {stage1_6[44]},
      {stage2_6[27]}
   );
   gpc1_1 gpc223 (
      {stage1_8[54]},
      {stage2_8[18]}
   );
   gpc1_1 gpc224 (
      {stage1_8[55]},
      {stage2_8[19]}
   );
   gpc1_1 gpc225 (
      {stage1_8[56]},
      {stage2_8[20]}
   );
   gpc1_1 gpc226 (
      {stage1_8[57]},
      {stage2_8[21]}
   );
   gpc1_1 gpc227 (
      {stage1_8[58]},
      {stage2_8[22]}
   );
   gpc1_1 gpc228 (
      {stage1_8[59]},
      {stage2_8[23]}
   );
   gpc1_1 gpc229 (
      {stage1_8[60]},
      {stage2_8[24]}
   );
   gpc1_1 gpc230 (
      {stage1_8[61]},
      {stage2_8[25]}
   );
   gpc1_1 gpc231 (
      {stage1_8[62]},
      {stage2_8[26]}
   );
   gpc1_1 gpc232 (
      {stage1_9[60]},
      {stage2_9[21]}
   );
   gpc1_1 gpc233 (
      {stage1_9[61]},
      {stage2_9[22]}
   );
   gpc1_1 gpc234 (
      {stage1_9[62]},
      {stage2_9[23]}
   );
   gpc1_1 gpc235 (
      {stage1_9[63]},
      {stage2_9[24]}
   );
   gpc1_1 gpc236 (
      {stage1_10[42]},
      {stage2_10[23]}
   );
   gpc1_1 gpc237 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc606_5 gpc239 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc240 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc241 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc242 (
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3],stage3_3[3]}
   );
   gpc615_5 gpc243 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc244 (
      {stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], 1'b0},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[5],stage3_3[5]}
   );
   gpc606_5 gpc245 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[6]}
   );
   gpc606_5 gpc246 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[7]}
   );
   gpc615_5 gpc247 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[18]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[8]}
   );
   gpc615_5 gpc248 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[7]}
   );
   gpc615_5 gpc249 (
      {stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27]},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[8]}
   );
   gpc615_5 gpc250 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[5],stage3_7[8]}
   );
   gpc615_5 gpc251 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[6],stage3_7[9]}
   );
   gpc615_5 gpc252 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[14]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[7],stage3_7[10]}
   );
   gpc615_5 gpc253 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[15]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[8],stage3_7[11]}
   );
   gpc606_5 gpc254 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[9]}
   );
   gpc615_5 gpc255 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_9[24]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc256 (
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[6],stage3_10[8]}
   );
   gpc615_5 gpc257 (
      {stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21]},
      {stage2_11[1]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[7],stage3_10[9]}
   );
   gpc606_5 gpc258 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[8]}
   );
   gpc606_5 gpc259 (
      {stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[9]}
   );
   gpc606_5 gpc260 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], 1'b0, 1'b0},
      {stage3_15[2],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[10]}
   );
   gpc606_5 gpc261 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[5],stage3_13[5],stage3_12[7]}
   );
   gpc1_1 gpc262 (
      {stage2_0[6]},
      {stage3_0[1]}
   );
   gpc1_1 gpc263 (
      {stage2_0[7]},
      {stage3_0[2]}
   );
   gpc1_1 gpc264 (
      {stage2_0[8]},
      {stage3_0[3]}
   );
   gpc1_1 gpc265 (
      {stage2_0[9]},
      {stage3_0[4]}
   );
   gpc1_1 gpc266 (
      {stage2_0[10]},
      {stage3_0[5]}
   );
   gpc1_1 gpc267 (
      {stage2_0[11]},
      {stage3_0[6]}
   );
   gpc1_1 gpc268 (
      {stage2_1[6]},
      {stage3_1[2]}
   );
   gpc1_1 gpc269 (
      {stage2_1[7]},
      {stage3_1[3]}
   );
   gpc1_1 gpc270 (
      {stage2_1[8]},
      {stage3_1[4]}
   );
   gpc1_1 gpc271 (
      {stage2_2[11]},
      {stage3_2[3]}
   );
   gpc1_1 gpc272 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc273 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc274 (
      {stage2_5[19]},
      {stage3_5[8]}
   );
   gpc1_1 gpc275 (
      {stage2_5[20]},
      {stage3_5[9]}
   );
   gpc1_1 gpc276 (
      {stage2_5[21]},
      {stage3_5[10]}
   );
   gpc1_1 gpc277 (
      {stage2_5[22]},
      {stage3_5[11]}
   );
   gpc1_1 gpc278 (
      {stage2_10[22]},
      {stage3_10[10]}
   );
   gpc1_1 gpc279 (
      {stage2_10[23]},
      {stage3_10[11]}
   );
   gpc1_1 gpc280 (
      {stage2_14[6]},
      {stage3_14[6]}
   );
   gpc1_1 gpc281 (
      {stage2_14[7]},
      {stage3_14[7]}
   );
   gpc1_1 gpc282 (
      {stage2_14[8]},
      {stage3_14[8]}
   );
   gpc1_1 gpc283 (
      {stage2_15[0]},
      {stage3_15[4]}
   );
   gpc1_1 gpc284 (
      {stage2_15[1]},
      {stage3_15[5]}
   );
   gpc1_1 gpc285 (
      {stage2_15[2]},
      {stage3_15[6]}
   );
   gpc1_1 gpc286 (
      {stage2_15[3]},
      {stage3_15[7]}
   );
   gpc606_5 gpc287 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], 1'b0},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc288 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc289 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2]}
   );
   gpc606_5 gpc290 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc291 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[2],stage4_8[3]}
   );
   gpc615_5 gpc292 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[3],stage4_8[4]}
   );
   gpc606_5 gpc293 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[4]}
   );
   gpc615_5 gpc294 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc295 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[4]}
   );
   gpc1163_5 gpc296 (
      {stage3_14[6], stage3_14[7], stage3_14[8]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage3_16[0]},
      {1'b0},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc1_1 gpc297 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc298 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc299 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc300 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc301 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc302 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc303 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc304 (
      {stage3_2[0]},
      {stage4_2[1]}
   );
   gpc1_1 gpc305 (
      {stage3_2[1]},
      {stage4_2[2]}
   );
   gpc1_1 gpc306 (
      {stage3_2[2]},
      {stage4_2[3]}
   );
   gpc1_1 gpc307 (
      {stage3_2[3]},
      {stage4_2[4]}
   );
   gpc1_1 gpc308 (
      {stage3_2[4]},
      {stage4_2[5]}
   );
   gpc1_1 gpc309 (
      {stage3_2[5]},
      {stage4_2[6]}
   );
   gpc1_1 gpc310 (
      {stage3_4[6]},
      {stage4_4[2]}
   );
   gpc1_1 gpc311 (
      {stage3_4[7]},
      {stage4_4[3]}
   );
   gpc1_1 gpc312 (
      {stage3_4[8]},
      {stage4_4[4]}
   );
   gpc1_1 gpc313 (
      {stage3_6[6]},
      {stage4_6[3]}
   );
   gpc1_1 gpc314 (
      {stage3_6[7]},
      {stage4_6[4]}
   );
   gpc1_1 gpc315 (
      {stage3_6[8]},
      {stage4_6[5]}
   );
   gpc1_1 gpc316 (
      {stage3_8[10]},
      {stage4_8[5]}
   );
   gpc1_1 gpc317 (
      {stage3_12[7]},
      {stage4_12[5]}
   );
   gpc1_1 gpc318 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc319 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc606_5 gpc320 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc321 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc615_5 gpc322 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc2135_5 gpc323 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1343_5 gpc324 (
      {stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1163_5 gpc325 (
      {stage4_14[1], stage4_14[2], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], 1'b0},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1_1 gpc326 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc327 (
      {stage4_1[0]},
      {stage5_1[1]}
   );
   gpc1_1 gpc328 (
      {stage4_2[6]},
      {stage5_2[1]}
   );
   gpc1_1 gpc329 (
      {stage4_3[0]},
      {stage5_3[1]}
   );
   gpc1_1 gpc330 (
      {stage4_5[3]},
      {stage5_5[1]}
   );
   gpc1_1 gpc331 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc332 (
      {stage4_18[0]},
      {stage5_18[1]}
   );
endmodule
module rowadder2_1_19(input [18:0] src0, input [18:0] src1, output [19:0] dst0);
    wire [18:0] gene;
    wire [18:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[18:16]}),
        .S({1'h0, prop[18:16]})
    );
    assign dst0 = {carryout[18], out[18:0]};
endmodule


module comp2_1test_128_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    reg [18:0] exp;
    wire [18:0] dst;
    assign test = dst == exp;
    compressor2_1_128_12 compressor2_1_128_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, dst, exp, test);
        src0 <= 12'hfa4;
        src1 <= 12'hd51;
        src2 <= 12'hf98;
        src3 <= 12'hb6e;
        src4 <= 12'hd54;
        src5 <= 12'h731;
        src6 <= 12'h95f;
        src7 <= 12'h354;
        src8 <= 12'h2e0;
        src9 <= 12'h711;
        src10 <= 12'hf85;
        src11 <= 12'h9d1;
        src12 <= 12'h1d2;
        src13 <= 12'h169;
        src14 <= 12'h735;
        src15 <= 12'h987;
        src16 <= 12'h1bb;
        src17 <= 12'ha69;
        src18 <= 12'h5b5;
        src19 <= 12'hc9a;
        src20 <= 12'hc40;
        src21 <= 12'h27a;
        src22 <= 12'hdd4;
        src23 <= 12'h44a;
        src24 <= 12'hf4a;
        src25 <= 12'hecc;
        src26 <= 12'h467;
        src27 <= 12'h40b;
        src28 <= 12'h1f8;
        src29 <= 12'haee;
        src30 <= 12'h7b0;
        src31 <= 12'hede;
        src32 <= 12'h71;
        src33 <= 12'hb83;
        src34 <= 12'hd9a;
        src35 <= 12'h905;
        src36 <= 12'h954;
        src37 <= 12'hdb6;
        src38 <= 12'h9a;
        src39 <= 12'h2aa;
        src40 <= 12'haa5;
        src41 <= 12'h217;
        src42 <= 12'heb8;
        src43 <= 12'hf51;
        src44 <= 12'h28c;
        src45 <= 12'h28;
        src46 <= 12'hc55;
        src47 <= 12'head;
        src48 <= 12'h573;
        src49 <= 12'hf53;
        src50 <= 12'h52e;
        src51 <= 12'h7f2;
        src52 <= 12'haa1;
        src53 <= 12'hb47;
        src54 <= 12'hccc;
        src55 <= 12'h245;
        src56 <= 12'h8a1;
        src57 <= 12'h8d6;
        src58 <= 12'h6da;
        src59 <= 12'ha2b;
        src60 <= 12'h386;
        src61 <= 12'h6be;
        src62 <= 12'hebd;
        src63 <= 12'hf6a;
        src64 <= 12'h52d;
        src65 <= 12'ha3f;
        src66 <= 12'he43;
        src67 <= 12'he88;
        src68 <= 12'haf7;
        src69 <= 12'h95a;
        src70 <= 12'h7d;
        src71 <= 12'hd08;
        src72 <= 12'hfe3;
        src73 <= 12'ha27;
        src74 <= 12'ha30;
        src75 <= 12'hb29;
        src76 <= 12'hb51;
        src77 <= 12'heba;
        src78 <= 12'h5e0;
        src79 <= 12'hc8d;
        src80 <= 12'hc2a;
        src81 <= 12'h3c4;
        src82 <= 12'had1;
        src83 <= 12'h2e9;
        src84 <= 12'hb6c;
        src85 <= 12'h2ba;
        src86 <= 12'h149;
        src87 <= 12'h949;
        src88 <= 12'h76f;
        src89 <= 12'h471;
        src90 <= 12'h438;
        src91 <= 12'hb93;
        src92 <= 12'hb08;
        src93 <= 12'h36e;
        src94 <= 12'hedb;
        src95 <= 12'hdae;
        src96 <= 12'h2ec;
        src97 <= 12'h405;
        src98 <= 12'h2ac;
        src99 <= 12'hca0;
        src100 <= 12'h74d;
        src101 <= 12'hb0a;
        src102 <= 12'h9f6;
        src103 <= 12'ha30;
        src104 <= 12'h46e;
        src105 <= 12'h70e;
        src106 <= 12'h6ed;
        src107 <= 12'hcfa;
        src108 <= 12'hd56;
        src109 <= 12'h9c;
        src110 <= 12'hdf8;
        src111 <= 12'h16c;
        src112 <= 12'h656;
        src113 <= 12'he87;
        src114 <= 12'hb73;
        src115 <= 12'hcc6;
        src116 <= 12'ha94;
        src117 <= 12'hbac;
        src118 <= 12'ha34;
        src119 <= 12'h476;
        src120 <= 12'h66a;
        src121 <= 12'h16f;
        src122 <= 12'h503;
        src123 <= 12'hdd0;
        src124 <= 12'h1c7;
        src125 <= 12'h763;
        src126 <= 12'h1db;
        src127 <= 12'hbce;
        exp <= 19'h454be;
        #1
        src0 <= 12'h95b;
        src1 <= 12'h9b0;
        src2 <= 12'h572;
        src3 <= 12'hb63;
        src4 <= 12'hbe8;
        src5 <= 12'hc66;
        src6 <= 12'hc6b;
        src7 <= 12'h44f;
        src8 <= 12'h8a3;
        src9 <= 12'h209;
        src10 <= 12'h6a7;
        src11 <= 12'hf2f;
        src12 <= 12'h108;
        src13 <= 12'h399;
        src14 <= 12'h507;
        src15 <= 12'hf6e;
        src16 <= 12'hf74;
        src17 <= 12'hcad;
        src18 <= 12'h53c;
        src19 <= 12'h1f0;
        src20 <= 12'hc97;
        src21 <= 12'h650;
        src22 <= 12'h36b;
        src23 <= 12'h8e1;
        src24 <= 12'h905;
        src25 <= 12'h9ab;
        src26 <= 12'h46c;
        src27 <= 12'h74d;
        src28 <= 12'h38f;
        src29 <= 12'hf9f;
        src30 <= 12'h5cd;
        src31 <= 12'hfe7;
        src32 <= 12'haf;
        src33 <= 12'h379;
        src34 <= 12'h8a5;
        src35 <= 12'h4cb;
        src36 <= 12'h3ba;
        src37 <= 12'h8ba;
        src38 <= 12'h2a7;
        src39 <= 12'h8de;
        src40 <= 12'h869;
        src41 <= 12'h6b4;
        src42 <= 12'h97a;
        src43 <= 12'h558;
        src44 <= 12'h9ff;
        src45 <= 12'h6fa;
        src46 <= 12'h842;
        src47 <= 12'h371;
        src48 <= 12'h3c2;
        src49 <= 12'h68d;
        src50 <= 12'h1a2;
        src51 <= 12'hdc0;
        src52 <= 12'h1b0;
        src53 <= 12'h675;
        src54 <= 12'h31e;
        src55 <= 12'h233;
        src56 <= 12'h89c;
        src57 <= 12'h10;
        src58 <= 12'he92;
        src59 <= 12'h3a;
        src60 <= 12'h2ad;
        src61 <= 12'h772;
        src62 <= 12'hfc0;
        src63 <= 12'h989;
        src64 <= 12'h250;
        src65 <= 12'hadb;
        src66 <= 12'hef1;
        src67 <= 12'h237;
        src68 <= 12'h2a0;
        src69 <= 12'h240;
        src70 <= 12'ha25;
        src71 <= 12'h490;
        src72 <= 12'h60;
        src73 <= 12'h25d;
        src74 <= 12'hee0;
        src75 <= 12'hf8c;
        src76 <= 12'hea6;
        src77 <= 12'he5d;
        src78 <= 12'hcea;
        src79 <= 12'hae;
        src80 <= 12'h99e;
        src81 <= 12'hc5f;
        src82 <= 12'ha84;
        src83 <= 12'hc20;
        src84 <= 12'h8ae;
        src85 <= 12'h7e8;
        src86 <= 12'h9e2;
        src87 <= 12'hfb6;
        src88 <= 12'h15e;
        src89 <= 12'hc0d;
        src90 <= 12'h41e;
        src91 <= 12'h14;
        src92 <= 12'h227;
        src93 <= 12'ha85;
        src94 <= 12'hf07;
        src95 <= 12'h58a;
        src96 <= 12'h780;
        src97 <= 12'h2cd;
        src98 <= 12'h1ff;
        src99 <= 12'hcb9;
        src100 <= 12'hb8e;
        src101 <= 12'h17;
        src102 <= 12'h49e;
        src103 <= 12'hb12;
        src104 <= 12'h581;
        src105 <= 12'h688;
        src106 <= 12'h316;
        src107 <= 12'hd6e;
        src108 <= 12'h93f;
        src109 <= 12'h9e3;
        src110 <= 12'hdb1;
        src111 <= 12'hed2;
        src112 <= 12'h4a7;
        src113 <= 12'hf5f;
        src114 <= 12'h751;
        src115 <= 12'h8e;
        src116 <= 12'hba0;
        src117 <= 12'h134;
        src118 <= 12'he38;
        src119 <= 12'hc30;
        src120 <= 12'hb95;
        src121 <= 12'h7a4;
        src122 <= 12'h538;
        src123 <= 12'h5ff;
        src124 <= 12'hcf3;
        src125 <= 12'hbe9;
        src126 <= 12'haf6;
        src127 <= 12'h80e;
        exp <= 19'h3ebd0;
        #1
        src0 <= 12'h86e;
        src1 <= 12'h31a;
        src2 <= 12'hcc8;
        src3 <= 12'h962;
        src4 <= 12'h3ec;
        src5 <= 12'h217;
        src6 <= 12'h7a6;
        src7 <= 12'h839;
        src8 <= 12'hb69;
        src9 <= 12'h701;
        src10 <= 12'h39b;
        src11 <= 12'he70;
        src12 <= 12'h79b;
        src13 <= 12'h6eb;
        src14 <= 12'h59c;
        src15 <= 12'h7c;
        src16 <= 12'hc0c;
        src17 <= 12'hbf2;
        src18 <= 12'h5a;
        src19 <= 12'hf32;
        src20 <= 12'h104;
        src21 <= 12'h598;
        src22 <= 12'hcbe;
        src23 <= 12'h9ce;
        src24 <= 12'h11c;
        src25 <= 12'h8a4;
        src26 <= 12'hd4c;
        src27 <= 12'h62e;
        src28 <= 12'hfcb;
        src29 <= 12'hebb;
        src30 <= 12'he53;
        src31 <= 12'h388;
        src32 <= 12'h846;
        src33 <= 12'heaa;
        src34 <= 12'hd4e;
        src35 <= 12'h6df;
        src36 <= 12'hc9a;
        src37 <= 12'h31b;
        src38 <= 12'h857;
        src39 <= 12'hc4b;
        src40 <= 12'h75a;
        src41 <= 12'he06;
        src42 <= 12'he8e;
        src43 <= 12'h329;
        src44 <= 12'ha16;
        src45 <= 12'h434;
        src46 <= 12'hef9;
        src47 <= 12'hc40;
        src48 <= 12'he4e;
        src49 <= 12'h94c;
        src50 <= 12'h26d;
        src51 <= 12'hc90;
        src52 <= 12'h888;
        src53 <= 12'hd69;
        src54 <= 12'h52e;
        src55 <= 12'h12f;
        src56 <= 12'h427;
        src57 <= 12'h88c;
        src58 <= 12'hd6b;
        src59 <= 12'hfd0;
        src60 <= 12'hb77;
        src61 <= 12'h4a3;
        src62 <= 12'h2bb;
        src63 <= 12'h622;
        src64 <= 12'h988;
        src65 <= 12'h68f;
        src66 <= 12'h362;
        src67 <= 12'hbc4;
        src68 <= 12'h97f;
        src69 <= 12'h47;
        src70 <= 12'hbb;
        src71 <= 12'h1df;
        src72 <= 12'h7fb;
        src73 <= 12'h7c5;
        src74 <= 12'h9e8;
        src75 <= 12'h26b;
        src76 <= 12'h3f7;
        src77 <= 12'hd72;
        src78 <= 12'hbd4;
        src79 <= 12'h2c6;
        src80 <= 12'ha2f;
        src81 <= 12'hf39;
        src82 <= 12'h969;
        src83 <= 12'h976;
        src84 <= 12'hf3c;
        src85 <= 12'hf91;
        src86 <= 12'hff4;
        src87 <= 12'h12;
        src88 <= 12'h7fe;
        src89 <= 12'hbda;
        src90 <= 12'h593;
        src91 <= 12'ha45;
        src92 <= 12'h8bb;
        src93 <= 12'h9b2;
        src94 <= 12'h509;
        src95 <= 12'h74;
        src96 <= 12'hdea;
        src97 <= 12'h18c;
        src98 <= 12'h2de;
        src99 <= 12'h626;
        src100 <= 12'h1fe;
        src101 <= 12'he91;
        src102 <= 12'h17;
        src103 <= 12'h1a5;
        src104 <= 12'h56f;
        src105 <= 12'h7f2;
        src106 <= 12'h5c8;
        src107 <= 12'hea1;
        src108 <= 12'h162;
        src109 <= 12'h289;
        src110 <= 12'hb74;
        src111 <= 12'hb48;
        src112 <= 12'hdf7;
        src113 <= 12'hc1;
        src114 <= 12'h115;
        src115 <= 12'had7;
        src116 <= 12'hba3;
        src117 <= 12'h2b;
        src118 <= 12'h12b;
        src119 <= 12'he40;
        src120 <= 12'h64f;
        src121 <= 12'h326;
        src122 <= 12'h877;
        src123 <= 12'hd0e;
        src124 <= 12'hdfd;
        src125 <= 12'h4bf;
        src126 <= 12'hd68;
        src127 <= 12'hb1f;
        exp <= 19'h40e83;
        #1
        src0 <= 12'h306;
        src1 <= 12'h17;
        src2 <= 12'h956;
        src3 <= 12'h531;
        src4 <= 12'hf7b;
        src5 <= 12'h95d;
        src6 <= 12'h215;
        src7 <= 12'h7b;
        src8 <= 12'hf7b;
        src9 <= 12'h4e9;
        src10 <= 12'h7d6;
        src11 <= 12'h53c;
        src12 <= 12'h3f7;
        src13 <= 12'h9fc;
        src14 <= 12'hd3;
        src15 <= 12'hd91;
        src16 <= 12'h49b;
        src17 <= 12'h419;
        src18 <= 12'hc0a;
        src19 <= 12'hda7;
        src20 <= 12'h7c3;
        src21 <= 12'hef9;
        src22 <= 12'hc23;
        src23 <= 12'ha33;
        src24 <= 12'hcc5;
        src25 <= 12'h62;
        src26 <= 12'h146;
        src27 <= 12'haeb;
        src28 <= 12'h2e4;
        src29 <= 12'hab6;
        src30 <= 12'h3ba;
        src31 <= 12'h648;
        src32 <= 12'hdda;
        src33 <= 12'h112;
        src34 <= 12'hb89;
        src35 <= 12'h5bf;
        src36 <= 12'h30c;
        src37 <= 12'hbf3;
        src38 <= 12'h8b;
        src39 <= 12'h9c7;
        src40 <= 12'ha19;
        src41 <= 12'h21f;
        src42 <= 12'h5c;
        src43 <= 12'h284;
        src44 <= 12'h76a;
        src45 <= 12'h8b7;
        src46 <= 12'hd0f;
        src47 <= 12'h99;
        src48 <= 12'h5b5;
        src49 <= 12'hc9a;
        src50 <= 12'h2f4;
        src51 <= 12'ha39;
        src52 <= 12'h4bb;
        src53 <= 12'ha40;
        src54 <= 12'h20b;
        src55 <= 12'h346;
        src56 <= 12'hba;
        src57 <= 12'h16;
        src58 <= 12'h4bc;
        src59 <= 12'ha8;
        src60 <= 12'h1cd;
        src61 <= 12'h49f;
        src62 <= 12'h9b7;
        src63 <= 12'h67b;
        src64 <= 12'h34f;
        src65 <= 12'h383;
        src66 <= 12'h776;
        src67 <= 12'hefd;
        src68 <= 12'h7f1;
        src69 <= 12'h545;
        src70 <= 12'h21e;
        src71 <= 12'ha9f;
        src72 <= 12'h1b;
        src73 <= 12'h95f;
        src74 <= 12'hbda;
        src75 <= 12'h25d;
        src76 <= 12'h842;
        src77 <= 12'h833;
        src78 <= 12'h710;
        src79 <= 12'h100;
        src80 <= 12'hef;
        src81 <= 12'hc6e;
        src82 <= 12'he4e;
        src83 <= 12'hb4c;
        src84 <= 12'ha60;
        src85 <= 12'h783;
        src86 <= 12'hd62;
        src87 <= 12'h38b;
        src88 <= 12'h8bb;
        src89 <= 12'hd69;
        src90 <= 12'h6c3;
        src91 <= 12'hc0a;
        src92 <= 12'hd84;
        src93 <= 12'h2c9;
        src94 <= 12'hbf2;
        src95 <= 12'h8e;
        src96 <= 12'hda9;
        src97 <= 12'h2a8;
        src98 <= 12'ha00;
        src99 <= 12'h29c;
        src100 <= 12'h5c3;
        src101 <= 12'h3fb;
        src102 <= 12'h856;
        src103 <= 12'h695;
        src104 <= 12'hca8;
        src105 <= 12'h4f7;
        src106 <= 12'ha83;
        src107 <= 12'h215;
        src108 <= 12'h54f;
        src109 <= 12'h8a2;
        src110 <= 12'h343;
        src111 <= 12'hf7;
        src112 <= 12'h339;
        src113 <= 12'h34f;
        src114 <= 12'h3c9;
        src115 <= 12'h409;
        src116 <= 12'hf6a;
        src117 <= 12'h83f;
        src118 <= 12'h261;
        src119 <= 12'h952;
        src120 <= 12'h9d5;
        src121 <= 12'h412;
        src122 <= 12'h47c;
        src123 <= 12'h1ed;
        src124 <= 12'hbfd;
        src125 <= 12'h191;
        src126 <= 12'h73b;
        src127 <= 12'hd9e;
        exp <= 19'h3679c;
        #1
        src0 <= 12'h55d;
        src1 <= 12'hdc5;
        src2 <= 12'h537;
        src3 <= 12'ha79;
        src4 <= 12'h18f;
        src5 <= 12'h770;
        src6 <= 12'h584;
        src7 <= 12'h34a;
        src8 <= 12'h850;
        src9 <= 12'h400;
        src10 <= 12'h479;
        src11 <= 12'hefd;
        src12 <= 12'h794;
        src13 <= 12'h1e0;
        src14 <= 12'h30;
        src15 <= 12'h244;
        src16 <= 12'h4e9;
        src17 <= 12'h3ec;
        src18 <= 12'h821;
        src19 <= 12'h432;
        src20 <= 12'h224;
        src21 <= 12'hffc;
        src22 <= 12'h820;
        src23 <= 12'hd00;
        src24 <= 12'heac;
        src25 <= 12'h74;
        src26 <= 12'hf18;
        src27 <= 12'hafc;
        src28 <= 12'h9e9;
        src29 <= 12'hbb;
        src30 <= 12'hee2;
        src31 <= 12'hf2f;
        src32 <= 12'hf95;
        src33 <= 12'h1ae;
        src34 <= 12'h9cb;
        src35 <= 12'h1aa;
        src36 <= 12'h63a;
        src37 <= 12'h315;
        src38 <= 12'hc7;
        src39 <= 12'hef;
        src40 <= 12'h58e;
        src41 <= 12'h918;
        src42 <= 12'h31c;
        src43 <= 12'h204;
        src44 <= 12'h2aa;
        src45 <= 12'h97d;
        src46 <= 12'hbb2;
        src47 <= 12'h788;
        src48 <= 12'h4a;
        src49 <= 12'h1b;
        src50 <= 12'h24f;
        src51 <= 12'h6c8;
        src52 <= 12'h51c;
        src53 <= 12'haba;
        src54 <= 12'ha43;
        src55 <= 12'h993;
        src56 <= 12'hc08;
        src57 <= 12'h858;
        src58 <= 12'h2eb;
        src59 <= 12'h7a6;
        src60 <= 12'h11d;
        src61 <= 12'hf7c;
        src62 <= 12'h4a4;
        src63 <= 12'h385;
        src64 <= 12'h714;
        src65 <= 12'ha2e;
        src66 <= 12'hd92;
        src67 <= 12'h519;
        src68 <= 12'hdfe;
        src69 <= 12'h764;
        src70 <= 12'h563;
        src71 <= 12'h126;
        src72 <= 12'h5af;
        src73 <= 12'hbb1;
        src74 <= 12'h41;
        src75 <= 12'hd8e;
        src76 <= 12'hf2a;
        src77 <= 12'h417;
        src78 <= 12'h685;
        src79 <= 12'hcff;
        src80 <= 12'hf4d;
        src81 <= 12'h231;
        src82 <= 12'hbc8;
        src83 <= 12'hdf0;
        src84 <= 12'hf20;
        src85 <= 12'hcb7;
        src86 <= 12'haf9;
        src87 <= 12'h561;
        src88 <= 12'h75a;
        src89 <= 12'h260;
        src90 <= 12'hfa0;
        src91 <= 12'h737;
        src92 <= 12'hecf;
        src93 <= 12'h19c;
        src94 <= 12'h474;
        src95 <= 12'h9b7;
        src96 <= 12'h773;
        src97 <= 12'hbe2;
        src98 <= 12'he1e;
        src99 <= 12'hec5;
        src100 <= 12'h7a1;
        src101 <= 12'h3ad;
        src102 <= 12'h9bc;
        src103 <= 12'h2d5;
        src104 <= 12'hee4;
        src105 <= 12'h900;
        src106 <= 12'h7f2;
        src107 <= 12'hfac;
        src108 <= 12'h411;
        src109 <= 12'hdc7;
        src110 <= 12'h363;
        src111 <= 12'hbde;
        src112 <= 12'h57;
        src113 <= 12'hd0;
        src114 <= 12'h113;
        src115 <= 12'h3e;
        src116 <= 12'he43;
        src117 <= 12'hd7f;
        src118 <= 12'h76d;
        src119 <= 12'h27;
        src120 <= 12'hcc8;
        src121 <= 12'h920;
        src122 <= 12'hea5;
        src123 <= 12'h7f1;
        src124 <= 12'hb9a;
        src125 <= 12'haa6;
        src126 <= 12'ha46;
        src127 <= 12'h40f;
        exp <= 19'h3da4a;
        #1
        src0 <= 12'h660;
        src1 <= 12'h5dd;
        src2 <= 12'h955;
        src3 <= 12'h651;
        src4 <= 12'h78f;
        src5 <= 12'he17;
        src6 <= 12'h3ff;
        src7 <= 12'h52e;
        src8 <= 12'h345;
        src9 <= 12'he17;
        src10 <= 12'h35f;
        src11 <= 12'hccc;
        src12 <= 12'h247;
        src13 <= 12'h3d0;
        src14 <= 12'h570;
        src15 <= 12'hf58;
        src16 <= 12'ha96;
        src17 <= 12'h2e7;
        src18 <= 12'h52;
        src19 <= 12'hf9;
        src20 <= 12'hcc0;
        src21 <= 12'h247;
        src22 <= 12'h5b5;
        src23 <= 12'h9fd;
        src24 <= 12'hc59;
        src25 <= 12'hf81;
        src26 <= 12'h16c;
        src27 <= 12'h983;
        src28 <= 12'h8ef;
        src29 <= 12'h4c4;
        src30 <= 12'ha3f;
        src31 <= 12'he81;
        src32 <= 12'h991;
        src33 <= 12'h453;
        src34 <= 12'h9e2;
        src35 <= 12'hf3a;
        src36 <= 12'h18b;
        src37 <= 12'hff8;
        src38 <= 12'h4b0;
        src39 <= 12'hc18;
        src40 <= 12'h388;
        src41 <= 12'h65b;
        src42 <= 12'h79;
        src43 <= 12'hbfc;
        src44 <= 12'h3b0;
        src45 <= 12'h50d;
        src46 <= 12'h7df;
        src47 <= 12'h22b;
        src48 <= 12'h344;
        src49 <= 12'h42a;
        src50 <= 12'h34e;
        src51 <= 12'h132;
        src52 <= 12'h69f;
        src53 <= 12'h8b8;
        src54 <= 12'h33;
        src55 <= 12'hb28;
        src56 <= 12'hce5;
        src57 <= 12'hd58;
        src58 <= 12'h63c;
        src59 <= 12'hded;
        src60 <= 12'h4c7;
        src61 <= 12'h891;
        src62 <= 12'h639;
        src63 <= 12'h730;
        src64 <= 12'h9f;
        src65 <= 12'hcda;
        src66 <= 12'h16a;
        src67 <= 12'h244;
        src68 <= 12'hc27;
        src69 <= 12'hc4;
        src70 <= 12'hd04;
        src71 <= 12'hacb;
        src72 <= 12'h9ff;
        src73 <= 12'hc8b;
        src74 <= 12'ha7c;
        src75 <= 12'h8c5;
        src76 <= 12'h9bc;
        src77 <= 12'h323;
        src78 <= 12'h1db;
        src79 <= 12'h19f;
        src80 <= 12'hac;
        src81 <= 12'hdb9;
        src82 <= 12'hc42;
        src83 <= 12'h368;
        src84 <= 12'h3fa;
        src85 <= 12'h47d;
        src86 <= 12'h349;
        src87 <= 12'hf2c;
        src88 <= 12'h48;
        src89 <= 12'ha85;
        src90 <= 12'hc64;
        src91 <= 12'h8db;
        src92 <= 12'hdc3;
        src93 <= 12'he89;
        src94 <= 12'h884;
        src95 <= 12'hc92;
        src96 <= 12'h9e3;
        src97 <= 12'h484;
        src98 <= 12'hfb1;
        src99 <= 12'h5a4;
        src100 <= 12'he1f;
        src101 <= 12'h33b;
        src102 <= 12'h3e6;
        src103 <= 12'h2c5;
        src104 <= 12'h140;
        src105 <= 12'h59f;
        src106 <= 12'hac;
        src107 <= 12'h43b;
        src108 <= 12'h7c5;
        src109 <= 12'h61c;
        src110 <= 12'h316;
        src111 <= 12'h2cc;
        src112 <= 12'h191;
        src113 <= 12'ha30;
        src114 <= 12'ha46;
        src115 <= 12'hd14;
        src116 <= 12'h8fd;
        src117 <= 12'h46b;
        src118 <= 12'hedb;
        src119 <= 12'hf13;
        src120 <= 12'h6b4;
        src121 <= 12'hc4e;
        src122 <= 12'hf11;
        src123 <= 12'hdb0;
        src124 <= 12'he6c;
        src125 <= 12'h209;
        src126 <= 12'h5c8;
        src127 <= 12'h447;
        exp <= 19'h3c27a;
        #1
        src0 <= 12'h81b;
        src1 <= 12'h9ad;
        src2 <= 12'h89e;
        src3 <= 12'heba;
        src4 <= 12'h558;
        src5 <= 12'heaa;
        src6 <= 12'h4e1;
        src7 <= 12'hfa;
        src8 <= 12'h9de;
        src9 <= 12'h6d4;
        src10 <= 12'h567;
        src11 <= 12'h323;
        src12 <= 12'h752;
        src13 <= 12'hbab;
        src14 <= 12'hf9f;
        src15 <= 12'h700;
        src16 <= 12'hd1;
        src17 <= 12'h8f6;
        src18 <= 12'hb5a;
        src19 <= 12'h70f;
        src20 <= 12'hdfa;
        src21 <= 12'ha80;
        src22 <= 12'h39c;
        src23 <= 12'h7f;
        src24 <= 12'h25b;
        src25 <= 12'h582;
        src26 <= 12'he55;
        src27 <= 12'hc1c;
        src28 <= 12'hadd;
        src29 <= 12'h748;
        src30 <= 12'hccd;
        src31 <= 12'h1eb;
        src32 <= 12'h1ec;
        src33 <= 12'ha23;
        src34 <= 12'h6df;
        src35 <= 12'hcc4;
        src36 <= 12'hd3a;
        src37 <= 12'ha67;
        src38 <= 12'hf2c;
        src39 <= 12'hec0;
        src40 <= 12'he63;
        src41 <= 12'h14f;
        src42 <= 12'h49d;
        src43 <= 12'h35a;
        src44 <= 12'h163;
        src45 <= 12'h48b;
        src46 <= 12'ha92;
        src47 <= 12'hfc8;
        src48 <= 12'h314;
        src49 <= 12'h427;
        src50 <= 12'h5e;
        src51 <= 12'hdc9;
        src52 <= 12'hbe4;
        src53 <= 12'h68a;
        src54 <= 12'haff;
        src55 <= 12'hdc3;
        src56 <= 12'h34;
        src57 <= 12'h65d;
        src58 <= 12'h289;
        src59 <= 12'hbc;
        src60 <= 12'hee0;
        src61 <= 12'h11;
        src62 <= 12'hfc0;
        src63 <= 12'hb91;
        src64 <= 12'h6b8;
        src65 <= 12'hbc8;
        src66 <= 12'h605;
        src67 <= 12'h161;
        src68 <= 12'hbed;
        src69 <= 12'h20d;
        src70 <= 12'hb8e;
        src71 <= 12'hff9;
        src72 <= 12'hc9;
        src73 <= 12'h927;
        src74 <= 12'habf;
        src75 <= 12'h98b;
        src76 <= 12'h5de;
        src77 <= 12'h6f2;
        src78 <= 12'h3a1;
        src79 <= 12'h877;
        src80 <= 12'ha7b;
        src81 <= 12'h392;
        src82 <= 12'hacc;
        src83 <= 12'h4f8;
        src84 <= 12'h81b;
        src85 <= 12'h6b9;
        src86 <= 12'hcfd;
        src87 <= 12'hf7;
        src88 <= 12'h32;
        src89 <= 12'hc0a;
        src90 <= 12'h60f;
        src91 <= 12'he17;
        src92 <= 12'hc52;
        src93 <= 12'hfe9;
        src94 <= 12'h27f;
        src95 <= 12'h6c4;
        src96 <= 12'h1f5;
        src97 <= 12'hecf;
        src98 <= 12'h6a1;
        src99 <= 12'h3b6;
        src100 <= 12'h2e3;
        src101 <= 12'h3e6;
        src102 <= 12'h827;
        src103 <= 12'h93;
        src104 <= 12'hd6d;
        src105 <= 12'h80c;
        src106 <= 12'h6ff;
        src107 <= 12'h60c;
        src108 <= 12'h7f3;
        src109 <= 12'hfe0;
        src110 <= 12'h3a6;
        src111 <= 12'hc03;
        src112 <= 12'h412;
        src113 <= 12'h720;
        src114 <= 12'hb85;
        src115 <= 12'h160;
        src116 <= 12'h197;
        src117 <= 12'hba6;
        src118 <= 12'h9ed;
        src119 <= 12'h66a;
        src120 <= 12'h44e;
        src121 <= 12'h86b;
        src122 <= 12'he1a;
        src123 <= 12'h445;
        src124 <= 12'h268;
        src125 <= 12'hd1f;
        src126 <= 12'h78;
        src127 <= 12'hc3c;
        exp <= 19'h3e43d;
        #1
        src0 <= 12'h1cd;
        src1 <= 12'hcc4;
        src2 <= 12'hd9a;
        src3 <= 12'h98c;
        src4 <= 12'he94;
        src5 <= 12'h47f;
        src6 <= 12'h730;
        src7 <= 12'hd15;
        src8 <= 12'h6ba;
        src9 <= 12'h2fe;
        src10 <= 12'hed;
        src11 <= 12'h806;
        src12 <= 12'h82e;
        src13 <= 12'h42e;
        src14 <= 12'h4a4;
        src15 <= 12'hcb4;
        src16 <= 12'he02;
        src17 <= 12'h9f3;
        src18 <= 12'hd08;
        src19 <= 12'h72a;
        src20 <= 12'h800;
        src21 <= 12'h395;
        src22 <= 12'h6d7;
        src23 <= 12'h298;
        src24 <= 12'he73;
        src25 <= 12'h842;
        src26 <= 12'h2a7;
        src27 <= 12'hc89;
        src28 <= 12'h9df;
        src29 <= 12'hb71;
        src30 <= 12'h4c9;
        src31 <= 12'ha35;
        src32 <= 12'h9d9;
        src33 <= 12'h7f1;
        src34 <= 12'h76f;
        src35 <= 12'h6f8;
        src36 <= 12'h9d4;
        src37 <= 12'h855;
        src38 <= 12'hd52;
        src39 <= 12'hdb;
        src40 <= 12'h23d;
        src41 <= 12'hcc7;
        src42 <= 12'hb35;
        src43 <= 12'hb03;
        src44 <= 12'h3b0;
        src45 <= 12'h559;
        src46 <= 12'h52f;
        src47 <= 12'he1d;
        src48 <= 12'h541;
        src49 <= 12'hd99;
        src50 <= 12'hddc;
        src51 <= 12'hca;
        src52 <= 12'h31a;
        src53 <= 12'h5b0;
        src54 <= 12'h42f;
        src55 <= 12'h596;
        src56 <= 12'hac3;
        src57 <= 12'hbe1;
        src58 <= 12'h2b8;
        src59 <= 12'ha6c;
        src60 <= 12'hba9;
        src61 <= 12'hb42;
        src62 <= 12'hd47;
        src63 <= 12'h28e;
        src64 <= 12'hda2;
        src65 <= 12'h24;
        src66 <= 12'ha9;
        src67 <= 12'h5ae;
        src68 <= 12'hcb7;
        src69 <= 12'h511;
        src70 <= 12'hc11;
        src71 <= 12'h6eb;
        src72 <= 12'h1bb;
        src73 <= 12'h96c;
        src74 <= 12'h42;
        src75 <= 12'h35f;
        src76 <= 12'ha5a;
        src77 <= 12'h6d1;
        src78 <= 12'h1f4;
        src79 <= 12'h169;
        src80 <= 12'hfdf;
        src81 <= 12'h879;
        src82 <= 12'h40e;
        src83 <= 12'h11;
        src84 <= 12'he14;
        src85 <= 12'h2f8;
        src86 <= 12'h1c6;
        src87 <= 12'h3f0;
        src88 <= 12'hc60;
        src89 <= 12'h607;
        src90 <= 12'h9b1;
        src91 <= 12'h90f;
        src92 <= 12'h230;
        src93 <= 12'hdd1;
        src94 <= 12'hc19;
        src95 <= 12'hfc4;
        src96 <= 12'hddd;
        src97 <= 12'h506;
        src98 <= 12'h3f9;
        src99 <= 12'hcff;
        src100 <= 12'h419;
        src101 <= 12'hb12;
        src102 <= 12'h5d9;
        src103 <= 12'hee7;
        src104 <= 12'h7d9;
        src105 <= 12'hf05;
        src106 <= 12'h8e1;
        src107 <= 12'h942;
        src108 <= 12'h46c;
        src109 <= 12'h56f;
        src110 <= 12'hde7;
        src111 <= 12'h448;
        src112 <= 12'h789;
        src113 <= 12'hbe2;
        src114 <= 12'h454;
        src115 <= 12'hbec;
        src116 <= 12'h40;
        src117 <= 12'h283;
        src118 <= 12'h86a;
        src119 <= 12'h18b;
        src120 <= 12'h3d2;
        src121 <= 12'h694;
        src122 <= 12'h2ed;
        src123 <= 12'h8c8;
        src124 <= 12'hd2b;
        src125 <= 12'hb7d;
        src126 <= 12'h82d;
        src127 <= 12'hb60;
        exp <= 19'h3e96e;
        #1
        src0 <= 12'h4aa;
        src1 <= 12'h194;
        src2 <= 12'ha35;
        src3 <= 12'h6ef;
        src4 <= 12'h178;
        src5 <= 12'h2f1;
        src6 <= 12'h7ef;
        src7 <= 12'hf9e;
        src8 <= 12'h56f;
        src9 <= 12'h679;
        src10 <= 12'hbd4;
        src11 <= 12'h140;
        src12 <= 12'h6d0;
        src13 <= 12'h57e;
        src14 <= 12'h7a8;
        src15 <= 12'h637;
        src16 <= 12'ha98;
        src17 <= 12'ha54;
        src18 <= 12'hce6;
        src19 <= 12'ha3d;
        src20 <= 12'h2e7;
        src21 <= 12'h539;
        src22 <= 12'h8dd;
        src23 <= 12'h920;
        src24 <= 12'h726;
        src25 <= 12'hf7b;
        src26 <= 12'h145;
        src27 <= 12'h9f1;
        src28 <= 12'hc87;
        src29 <= 12'h776;
        src30 <= 12'h316;
        src31 <= 12'h146;
        src32 <= 12'h57f;
        src33 <= 12'he38;
        src34 <= 12'h163;
        src35 <= 12'had2;
        src36 <= 12'h78b;
        src37 <= 12'hb7b;
        src38 <= 12'h7d2;
        src39 <= 12'ha4b;
        src40 <= 12'h5aa;
        src41 <= 12'h8de;
        src42 <= 12'h893;
        src43 <= 12'h85;
        src44 <= 12'h80e;
        src45 <= 12'h6e4;
        src46 <= 12'h5c2;
        src47 <= 12'hf9d;
        src48 <= 12'h28e;
        src49 <= 12'h128;
        src50 <= 12'hc37;
        src51 <= 12'hc01;
        src52 <= 12'h524;
        src53 <= 12'h907;
        src54 <= 12'hdf4;
        src55 <= 12'h99f;
        src56 <= 12'hb48;
        src57 <= 12'ha28;
        src58 <= 12'h10c;
        src59 <= 12'h56d;
        src60 <= 12'hc92;
        src61 <= 12'h8a5;
        src62 <= 12'h9ab;
        src63 <= 12'h4a7;
        src64 <= 12'h77a;
        src65 <= 12'hcf6;
        src66 <= 12'hbb0;
        src67 <= 12'hd7e;
        src68 <= 12'h5bc;
        src69 <= 12'h67a;
        src70 <= 12'h259;
        src71 <= 12'h83c;
        src72 <= 12'h94a;
        src73 <= 12'hf9e;
        src74 <= 12'h826;
        src75 <= 12'h7c6;
        src76 <= 12'h2c3;
        src77 <= 12'hb3e;
        src78 <= 12'h590;
        src79 <= 12'h8bb;
        src80 <= 12'h206;
        src81 <= 12'h473;
        src82 <= 12'ha47;
        src83 <= 12'hdb9;
        src84 <= 12'h75a;
        src85 <= 12'hdab;
        src86 <= 12'h49f;
        src87 <= 12'h667;
        src88 <= 12'h3bb;
        src89 <= 12'hc8a;
        src90 <= 12'hbfc;
        src91 <= 12'h497;
        src92 <= 12'h45f;
        src93 <= 12'h641;
        src94 <= 12'hfff;
        src95 <= 12'h9f3;
        src96 <= 12'hffe;
        src97 <= 12'h763;
        src98 <= 12'h7d7;
        src99 <= 12'h5b;
        src100 <= 12'h43d;
        src101 <= 12'had6;
        src102 <= 12'h265;
        src103 <= 12'h609;
        src104 <= 12'h48d;
        src105 <= 12'h442;
        src106 <= 12'h55a;
        src107 <= 12'h9a9;
        src108 <= 12'ha77;
        src109 <= 12'h99;
        src110 <= 12'h278;
        src111 <= 12'hbcb;
        src112 <= 12'hd6f;
        src113 <= 12'hfcf;
        src114 <= 12'hc24;
        src115 <= 12'hc6e;
        src116 <= 12'ha7e;
        src117 <= 12'ha0b;
        src118 <= 12'he58;
        src119 <= 12'hf07;
        src120 <= 12'h4ad;
        src121 <= 12'hf3e;
        src122 <= 12'h97b;
        src123 <= 12'hb08;
        src124 <= 12'h713;
        src125 <= 12'h893;
        src126 <= 12'hfa3;
        src127 <= 12'hcd4;
        exp <= 19'h41aee;
        #1
        src0 <= 12'h7bf;
        src1 <= 12'h917;
        src2 <= 12'h6e6;
        src3 <= 12'hb1b;
        src4 <= 12'h8c8;
        src5 <= 12'h6fd;
        src6 <= 12'hcad;
        src7 <= 12'h36c;
        src8 <= 12'h803;
        src9 <= 12'he4f;
        src10 <= 12'h6c6;
        src11 <= 12'hac8;
        src12 <= 12'hbc3;
        src13 <= 12'hc07;
        src14 <= 12'hb09;
        src15 <= 12'h3b8;
        src16 <= 12'h136;
        src17 <= 12'h62d;
        src18 <= 12'h50a;
        src19 <= 12'hffc;
        src20 <= 12'h431;
        src21 <= 12'hba1;
        src22 <= 12'h7c7;
        src23 <= 12'haa9;
        src24 <= 12'h86d;
        src25 <= 12'h3a3;
        src26 <= 12'he7e;
        src27 <= 12'haac;
        src28 <= 12'hb2f;
        src29 <= 12'h73c;
        src30 <= 12'hdd1;
        src31 <= 12'hba;
        src32 <= 12'hb08;
        src33 <= 12'ha66;
        src34 <= 12'hab8;
        src35 <= 12'h16f;
        src36 <= 12'h54e;
        src37 <= 12'hc42;
        src38 <= 12'h333;
        src39 <= 12'hb40;
        src40 <= 12'ha7b;
        src41 <= 12'h85b;
        src42 <= 12'hc13;
        src43 <= 12'hcb4;
        src44 <= 12'h5f4;
        src45 <= 12'h4a4;
        src46 <= 12'h460;
        src47 <= 12'h95f;
        src48 <= 12'hc3f;
        src49 <= 12'he09;
        src50 <= 12'h93f;
        src51 <= 12'h6df;
        src52 <= 12'h61a;
        src53 <= 12'hb71;
        src54 <= 12'ha59;
        src55 <= 12'he7c;
        src56 <= 12'h19a;
        src57 <= 12'h727;
        src58 <= 12'h474;
        src59 <= 12'he39;
        src60 <= 12'hca9;
        src61 <= 12'he19;
        src62 <= 12'h32c;
        src63 <= 12'hab;
        src64 <= 12'h68e;
        src65 <= 12'h9fe;
        src66 <= 12'hfb1;
        src67 <= 12'h586;
        src68 <= 12'h1bb;
        src69 <= 12'hbec;
        src70 <= 12'h397;
        src71 <= 12'hbcc;
        src72 <= 12'h22e;
        src73 <= 12'h1e9;
        src74 <= 12'h6d5;
        src75 <= 12'h9b6;
        src76 <= 12'hea8;
        src77 <= 12'h239;
        src78 <= 12'h6d4;
        src79 <= 12'h255;
        src80 <= 12'h53c;
        src81 <= 12'he4c;
        src82 <= 12'h568;
        src83 <= 12'h410;
        src84 <= 12'hc2d;
        src85 <= 12'h675;
        src86 <= 12'hc01;
        src87 <= 12'h6eb;
        src88 <= 12'h5e7;
        src89 <= 12'hd53;
        src90 <= 12'hd6e;
        src91 <= 12'h77d;
        src92 <= 12'hd64;
        src93 <= 12'h8db;
        src94 <= 12'h6ba;
        src95 <= 12'h48e;
        src96 <= 12'he17;
        src97 <= 12'h501;
        src98 <= 12'he26;
        src99 <= 12'ha0d;
        src100 <= 12'h4fd;
        src101 <= 12'hbd5;
        src102 <= 12'h3cf;
        src103 <= 12'h4c2;
        src104 <= 12'h740;
        src105 <= 12'h532;
        src106 <= 12'hdb4;
        src107 <= 12'h770;
        src108 <= 12'hbfa;
        src109 <= 12'hb7a;
        src110 <= 12'h73d;
        src111 <= 12'hff7;
        src112 <= 12'h2d1;
        src113 <= 12'h4e4;
        src114 <= 12'h821;
        src115 <= 12'hab8;
        src116 <= 12'ha7c;
        src117 <= 12'h1ad;
        src118 <= 12'h9a9;
        src119 <= 12'h5b0;
        src120 <= 12'h557;
        src121 <= 12'h9d6;
        src122 <= 12'h5c7;
        src123 <= 12'he27;
        src124 <= 12'h8f2;
        src125 <= 12'h3e;
        src126 <= 12'h23a;
        src127 <= 12'h4f3;
        exp <= 19'h4267b;
        #1
        src0 <= 12'h657;
        src1 <= 12'hd45;
        src2 <= 12'hb4b;
        src3 <= 12'h69;
        src4 <= 12'he4a;
        src5 <= 12'h9ee;
        src6 <= 12'h98b;
        src7 <= 12'h6bb;
        src8 <= 12'heea;
        src9 <= 12'h712;
        src10 <= 12'h300;
        src11 <= 12'hd3e;
        src12 <= 12'h7dd;
        src13 <= 12'h822;
        src14 <= 12'h32e;
        src15 <= 12'h648;
        src16 <= 12'h77;
        src17 <= 12'h814;
        src18 <= 12'hcff;
        src19 <= 12'h325;
        src20 <= 12'h48;
        src21 <= 12'he4;
        src22 <= 12'h210;
        src23 <= 12'h9ae;
        src24 <= 12'h813;
        src25 <= 12'ha0;
        src26 <= 12'hc8f;
        src27 <= 12'h7ec;
        src28 <= 12'hf12;
        src29 <= 12'h425;
        src30 <= 12'hfa4;
        src31 <= 12'h3e4;
        src32 <= 12'h5a4;
        src33 <= 12'h7a3;
        src34 <= 12'h6;
        src35 <= 12'h460;
        src36 <= 12'ha82;
        src37 <= 12'hc64;
        src38 <= 12'hc90;
        src39 <= 12'h991;
        src40 <= 12'h3fa;
        src41 <= 12'ha33;
        src42 <= 12'ha23;
        src43 <= 12'h4e;
        src44 <= 12'h738;
        src45 <= 12'h7bf;
        src46 <= 12'h4a2;
        src47 <= 12'hd4c;
        src48 <= 12'hd90;
        src49 <= 12'h494;
        src50 <= 12'hd8f;
        src51 <= 12'h7f;
        src52 <= 12'hcb0;
        src53 <= 12'h40b;
        src54 <= 12'h296;
        src55 <= 12'haec;
        src56 <= 12'h113;
        src57 <= 12'h9b6;
        src58 <= 12'h6db;
        src59 <= 12'h899;
        src60 <= 12'had4;
        src61 <= 12'hdf2;
        src62 <= 12'hc46;
        src63 <= 12'hab2;
        src64 <= 12'ha1d;
        src65 <= 12'h3e;
        src66 <= 12'h251;
        src67 <= 12'h438;
        src68 <= 12'h885;
        src69 <= 12'h2f;
        src70 <= 12'h105;
        src71 <= 12'h7c1;
        src72 <= 12'hd6b;
        src73 <= 12'ha45;
        src74 <= 12'h60;
        src75 <= 12'ha9d;
        src76 <= 12'hafb;
        src77 <= 12'h5ae;
        src78 <= 12'h69;
        src79 <= 12'h33f;
        src80 <= 12'h27d;
        src81 <= 12'he67;
        src82 <= 12'hfbc;
        src83 <= 12'h3bf;
        src84 <= 12'h49;
        src85 <= 12'he04;
        src86 <= 12'h537;
        src87 <= 12'hb28;
        src88 <= 12'h27a;
        src89 <= 12'h172;
        src90 <= 12'h1ce;
        src91 <= 12'h5a7;
        src92 <= 12'hada;
        src93 <= 12'hf8;
        src94 <= 12'hf70;
        src95 <= 12'h3c4;
        src96 <= 12'hfef;
        src97 <= 12'h56e;
        src98 <= 12'ha5c;
        src99 <= 12'h8af;
        src100 <= 12'h251;
        src101 <= 12'h82;
        src102 <= 12'h538;
        src103 <= 12'h546;
        src104 <= 12'h585;
        src105 <= 12'ha1;
        src106 <= 12'h991;
        src107 <= 12'h44b;
        src108 <= 12'h6d4;
        src109 <= 12'h97c;
        src110 <= 12'h3db;
        src111 <= 12'h39;
        src112 <= 12'ha2e;
        src113 <= 12'h6d4;
        src114 <= 12'h644;
        src115 <= 12'h363;
        src116 <= 12'hfb1;
        src117 <= 12'h159;
        src118 <= 12'h265;
        src119 <= 12'h16c;
        src120 <= 12'h42b;
        src121 <= 12'h4b7;
        src122 <= 12'haf4;
        src123 <= 12'h115;
        src124 <= 12'hb61;
        src125 <= 12'he1f;
        src126 <= 12'h61b;
        src127 <= 12'hda4;
        exp <= 19'h3883f;
        #1
        src0 <= 12'ha71;
        src1 <= 12'h9b3;
        src2 <= 12'h748;
        src3 <= 12'h34;
        src4 <= 12'hdfd;
        src5 <= 12'h760;
        src6 <= 12'h2e9;
        src7 <= 12'h475;
        src8 <= 12'h719;
        src9 <= 12'h73f;
        src10 <= 12'hbbc;
        src11 <= 12'hf91;
        src12 <= 12'hf41;
        src13 <= 12'hb20;
        src14 <= 12'h3f7;
        src15 <= 12'h710;
        src16 <= 12'heec;
        src17 <= 12'h84a;
        src18 <= 12'h57c;
        src19 <= 12'hf1;
        src20 <= 12'he5c;
        src21 <= 12'h2d;
        src22 <= 12'h8dc;
        src23 <= 12'h64d;
        src24 <= 12'h1d9;
        src25 <= 12'hbfb;
        src26 <= 12'h923;
        src27 <= 12'h257;
        src28 <= 12'h86;
        src29 <= 12'ha34;
        src30 <= 12'hb7a;
        src31 <= 12'hf42;
        src32 <= 12'h95b;
        src33 <= 12'hb18;
        src34 <= 12'h941;
        src35 <= 12'h50;
        src36 <= 12'h58f;
        src37 <= 12'h517;
        src38 <= 12'h40b;
        src39 <= 12'h6ec;
        src40 <= 12'h5f8;
        src41 <= 12'ha38;
        src42 <= 12'hb5f;
        src43 <= 12'hb3c;
        src44 <= 12'h604;
        src45 <= 12'hc27;
        src46 <= 12'h832;
        src47 <= 12'hc8e;
        src48 <= 12'ha32;
        src49 <= 12'hd11;
        src50 <= 12'h799;
        src51 <= 12'h1f8;
        src52 <= 12'h430;
        src53 <= 12'hdbf;
        src54 <= 12'hfc8;
        src55 <= 12'h45b;
        src56 <= 12'hecb;
        src57 <= 12'h233;
        src58 <= 12'h9df;
        src59 <= 12'h9b7;
        src60 <= 12'ha89;
        src61 <= 12'hf64;
        src62 <= 12'h730;
        src63 <= 12'heba;
        src64 <= 12'h8b1;
        src65 <= 12'hffd;
        src66 <= 12'he60;
        src67 <= 12'hf99;
        src68 <= 12'h11d;
        src69 <= 12'hcf3;
        src70 <= 12'hadf;
        src71 <= 12'ha8;
        src72 <= 12'hcb6;
        src73 <= 12'h512;
        src74 <= 12'h605;
        src75 <= 12'h1a3;
        src76 <= 12'h705;
        src77 <= 12'hbf8;
        src78 <= 12'h97a;
        src79 <= 12'hd44;
        src80 <= 12'h5fd;
        src81 <= 12'h95f;
        src82 <= 12'hf55;
        src83 <= 12'h6b4;
        src84 <= 12'h45f;
        src85 <= 12'h2a4;
        src86 <= 12'h227;
        src87 <= 12'he1a;
        src88 <= 12'hd28;
        src89 <= 12'h411;
        src90 <= 12'h22f;
        src91 <= 12'hf59;
        src92 <= 12'h54d;
        src93 <= 12'h4fd;
        src94 <= 12'h4fb;
        src95 <= 12'h91f;
        src96 <= 12'h5cc;
        src97 <= 12'hf82;
        src98 <= 12'hbc7;
        src99 <= 12'h6f6;
        src100 <= 12'hb25;
        src101 <= 12'h822;
        src102 <= 12'h4d6;
        src103 <= 12'h2ea;
        src104 <= 12'h1cc;
        src105 <= 12'h12a;
        src106 <= 12'h8e7;
        src107 <= 12'hd6b;
        src108 <= 12'hc37;
        src109 <= 12'h6ce;
        src110 <= 12'h5dd;
        src111 <= 12'h92;
        src112 <= 12'h46d;
        src113 <= 12'h726;
        src114 <= 12'hd21;
        src115 <= 12'hcad;
        src116 <= 12'hf6;
        src117 <= 12'hf5a;
        src118 <= 12'h85a;
        src119 <= 12'hea7;
        src120 <= 12'h496;
        src121 <= 12'h2ab;
        src122 <= 12'h3cc;
        src123 <= 12'h381;
        src124 <= 12'h5f2;
        src125 <= 12'h860;
        src126 <= 12'h6ed;
        src127 <= 12'h87a;
        exp <= 19'h41827;
        #1
        src0 <= 12'hdc7;
        src1 <= 12'hf69;
        src2 <= 12'h541;
        src3 <= 12'hf0e;
        src4 <= 12'hbd1;
        src5 <= 12'h1e1;
        src6 <= 12'hee4;
        src7 <= 12'h6af;
        src8 <= 12'h7dd;
        src9 <= 12'h6e9;
        src10 <= 12'h8f1;
        src11 <= 12'h820;
        src12 <= 12'h6ec;
        src13 <= 12'he17;
        src14 <= 12'h3ce;
        src15 <= 12'hf21;
        src16 <= 12'h35b;
        src17 <= 12'hfab;
        src18 <= 12'h1c3;
        src19 <= 12'h2ca;
        src20 <= 12'h5ec;
        src21 <= 12'hd36;
        src22 <= 12'h90a;
        src23 <= 12'hc5c;
        src24 <= 12'h13c;
        src25 <= 12'h377;
        src26 <= 12'h474;
        src27 <= 12'hb83;
        src28 <= 12'hadd;
        src29 <= 12'h33a;
        src30 <= 12'h600;
        src31 <= 12'h3df;
        src32 <= 12'h6d4;
        src33 <= 12'h19b;
        src34 <= 12'h661;
        src35 <= 12'hccb;
        src36 <= 12'hcf6;
        src37 <= 12'h22b;
        src38 <= 12'he53;
        src39 <= 12'h546;
        src40 <= 12'h6b;
        src41 <= 12'hbb6;
        src42 <= 12'h448;
        src43 <= 12'h326;
        src44 <= 12'hfd5;
        src45 <= 12'h5ac;
        src46 <= 12'h247;
        src47 <= 12'h148;
        src48 <= 12'ha2f;
        src49 <= 12'h25c;
        src50 <= 12'h7a8;
        src51 <= 12'h848;
        src52 <= 12'h6c1;
        src53 <= 12'h1a1;
        src54 <= 12'h4db;
        src55 <= 12'h841;
        src56 <= 12'h2d7;
        src57 <= 12'hfaf;
        src58 <= 12'h8ef;
        src59 <= 12'hff3;
        src60 <= 12'h5cd;
        src61 <= 12'h5f0;
        src62 <= 12'h599;
        src63 <= 12'h11e;
        src64 <= 12'h658;
        src65 <= 12'hca8;
        src66 <= 12'h30a;
        src67 <= 12'hcc3;
        src68 <= 12'h2ae;
        src69 <= 12'h9b5;
        src70 <= 12'h458;
        src71 <= 12'ha88;
        src72 <= 12'haf9;
        src73 <= 12'h2a5;
        src74 <= 12'ha8c;
        src75 <= 12'h807;
        src76 <= 12'hff4;
        src77 <= 12'ha7d;
        src78 <= 12'ha22;
        src79 <= 12'hb95;
        src80 <= 12'h9d1;
        src81 <= 12'h3a7;
        src82 <= 12'ha45;
        src83 <= 12'ha01;
        src84 <= 12'hc04;
        src85 <= 12'hb5e;
        src86 <= 12'h517;
        src87 <= 12'h20d;
        src88 <= 12'hb15;
        src89 <= 12'hf54;
        src90 <= 12'h7ea;
        src91 <= 12'h2c8;
        src92 <= 12'hf27;
        src93 <= 12'h5a9;
        src94 <= 12'h793;
        src95 <= 12'h659;
        src96 <= 12'h129;
        src97 <= 12'h73a;
        src98 <= 12'h7ec;
        src99 <= 12'he8a;
        src100 <= 12'ha47;
        src101 <= 12'hc59;
        src102 <= 12'h3ee;
        src103 <= 12'hdc3;
        src104 <= 12'hd8b;
        src105 <= 12'he18;
        src106 <= 12'hd15;
        src107 <= 12'h975;
        src108 <= 12'he3;
        src109 <= 12'hb4;
        src110 <= 12'he47;
        src111 <= 12'hfeb;
        src112 <= 12'hc91;
        src113 <= 12'ha4f;
        src114 <= 12'h5b6;
        src115 <= 12'h8c8;
        src116 <= 12'h946;
        src117 <= 12'h756;
        src118 <= 12'h510;
        src119 <= 12'h59a;
        src120 <= 12'h309;
        src121 <= 12'he38;
        src122 <= 12'h914;
        src123 <= 12'h93e;
        src124 <= 12'hb0f;
        src125 <= 12'h681;
        src126 <= 12'h8;
        src127 <= 12'ha99;
        exp <= 19'h4141d;
        #1
        src0 <= 12'he36;
        src1 <= 12'h5c5;
        src2 <= 12'h5f4;
        src3 <= 12'h885;
        src4 <= 12'h2a6;
        src5 <= 12'h7b0;
        src6 <= 12'h8b2;
        src7 <= 12'h44;
        src8 <= 12'h94a;
        src9 <= 12'hd65;
        src10 <= 12'h858;
        src11 <= 12'h3a5;
        src12 <= 12'hecd;
        src13 <= 12'h4f2;
        src14 <= 12'hbba;
        src15 <= 12'he88;
        src16 <= 12'hb03;
        src17 <= 12'h205;
        src18 <= 12'h553;
        src19 <= 12'h72e;
        src20 <= 12'h3cc;
        src21 <= 12'h32e;
        src22 <= 12'hfc;
        src23 <= 12'hac2;
        src24 <= 12'hd57;
        src25 <= 12'h578;
        src26 <= 12'hb75;
        src27 <= 12'he10;
        src28 <= 12'h3f4;
        src29 <= 12'h2d5;
        src30 <= 12'h6a8;
        src31 <= 12'h454;
        src32 <= 12'hbb8;
        src33 <= 12'h3c1;
        src34 <= 12'h7f6;
        src35 <= 12'hedb;
        src36 <= 12'h6a8;
        src37 <= 12'h3b7;
        src38 <= 12'hbef;
        src39 <= 12'ha6f;
        src40 <= 12'h6ba;
        src41 <= 12'h671;
        src42 <= 12'h24d;
        src43 <= 12'h36f;
        src44 <= 12'h3e1;
        src45 <= 12'h9ce;
        src46 <= 12'h222;
        src47 <= 12'hd59;
        src48 <= 12'h670;
        src49 <= 12'h61c;
        src50 <= 12'hc48;
        src51 <= 12'hf3e;
        src52 <= 12'hc3d;
        src53 <= 12'h883;
        src54 <= 12'hb2e;
        src55 <= 12'hb32;
        src56 <= 12'hc9b;
        src57 <= 12'h2f4;
        src58 <= 12'h55c;
        src59 <= 12'h749;
        src60 <= 12'hf77;
        src61 <= 12'hd54;
        src62 <= 12'hc53;
        src63 <= 12'haf0;
        src64 <= 12'hf13;
        src65 <= 12'h7ae;
        src66 <= 12'ha8f;
        src67 <= 12'h43b;
        src68 <= 12'hc7d;
        src69 <= 12'hef3;
        src70 <= 12'h84a;
        src71 <= 12'ha84;
        src72 <= 12'h410;
        src73 <= 12'ha7c;
        src74 <= 12'hc36;
        src75 <= 12'h957;
        src76 <= 12'h7b;
        src77 <= 12'h3a9;
        src78 <= 12'h9c;
        src79 <= 12'he22;
        src80 <= 12'heb5;
        src81 <= 12'h1fd;
        src82 <= 12'hb;
        src83 <= 12'haf2;
        src84 <= 12'h340;
        src85 <= 12'h843;
        src86 <= 12'h31;
        src87 <= 12'hd7e;
        src88 <= 12'h4d0;
        src89 <= 12'he4b;
        src90 <= 12'hdd0;
        src91 <= 12'h28d;
        src92 <= 12'hf0b;
        src93 <= 12'h305;
        src94 <= 12'h7bb;
        src95 <= 12'haa6;
        src96 <= 12'h4ee;
        src97 <= 12'hb32;
        src98 <= 12'hc42;
        src99 <= 12'h988;
        src100 <= 12'h8e;
        src101 <= 12'h18e;
        src102 <= 12'hf70;
        src103 <= 12'h10e;
        src104 <= 12'he4f;
        src105 <= 12'h782;
        src106 <= 12'hd7;
        src107 <= 12'h978;
        src108 <= 12'hcaa;
        src109 <= 12'h3db;
        src110 <= 12'hb36;
        src111 <= 12'hc9e;
        src112 <= 12'hb0c;
        src113 <= 12'h63d;
        src114 <= 12'ha88;
        src115 <= 12'h956;
        src116 <= 12'hd5d;
        src117 <= 12'h71c;
        src118 <= 12'h1a2;
        src119 <= 12'h746;
        src120 <= 12'hdcb;
        src121 <= 12'h750;
        src122 <= 12'h8d7;
        src123 <= 12'h372;
        src124 <= 12'h127;
        src125 <= 12'h6c2;
        src126 <= 12'hf69;
        src127 <= 12'h956;
        exp <= 19'h41872;
        #1
        src0 <= 12'hcad;
        src1 <= 12'h5a;
        src2 <= 12'hd32;
        src3 <= 12'h9f9;
        src4 <= 12'h5b;
        src5 <= 12'h5df;
        src6 <= 12'ha99;
        src7 <= 12'ha6;
        src8 <= 12'hc6e;
        src9 <= 12'h4bd;
        src10 <= 12'ha53;
        src11 <= 12'haeb;
        src12 <= 12'h27c;
        src13 <= 12'hf20;
        src14 <= 12'h3fd;
        src15 <= 12'h4c3;
        src16 <= 12'h9c6;
        src17 <= 12'h226;
        src18 <= 12'h617;
        src19 <= 12'h4e9;
        src20 <= 12'h519;
        src21 <= 12'hb76;
        src22 <= 12'he4a;
        src23 <= 12'h9a3;
        src24 <= 12'hc2d;
        src25 <= 12'h334;
        src26 <= 12'ha29;
        src27 <= 12'h459;
        src28 <= 12'h7c1;
        src29 <= 12'h2a5;
        src30 <= 12'h4b7;
        src31 <= 12'hbb4;
        src32 <= 12'h26e;
        src33 <= 12'h4f;
        src34 <= 12'h83b;
        src35 <= 12'h13c;
        src36 <= 12'h34a;
        src37 <= 12'ha77;
        src38 <= 12'h71d;
        src39 <= 12'h83d;
        src40 <= 12'hb74;
        src41 <= 12'hd27;
        src42 <= 12'h9d9;
        src43 <= 12'h38f;
        src44 <= 12'hc35;
        src45 <= 12'hdd9;
        src46 <= 12'h844;
        src47 <= 12'h4b;
        src48 <= 12'h397;
        src49 <= 12'h6fa;
        src50 <= 12'he27;
        src51 <= 12'h2d4;
        src52 <= 12'h55e;
        src53 <= 12'hdc5;
        src54 <= 12'h2fb;
        src55 <= 12'h285;
        src56 <= 12'h147;
        src57 <= 12'ha6;
        src58 <= 12'h4d6;
        src59 <= 12'hd21;
        src60 <= 12'h204;
        src61 <= 12'h179;
        src62 <= 12'hec;
        src63 <= 12'h51f;
        src64 <= 12'h228;
        src65 <= 12'hc15;
        src66 <= 12'h1c6;
        src67 <= 12'h6e8;
        src68 <= 12'h803;
        src69 <= 12'he61;
        src70 <= 12'h519;
        src71 <= 12'h16f;
        src72 <= 12'h34d;
        src73 <= 12'h4a9;
        src74 <= 12'hce7;
        src75 <= 12'h361;
        src76 <= 12'h112;
        src77 <= 12'hd47;
        src78 <= 12'h70;
        src79 <= 12'h934;
        src80 <= 12'h2b3;
        src81 <= 12'h858;
        src82 <= 12'h474;
        src83 <= 12'h6ba;
        src84 <= 12'h533;
        src85 <= 12'h981;
        src86 <= 12'h2f9;
        src87 <= 12'h88a;
        src88 <= 12'hb99;
        src89 <= 12'h5ba;
        src90 <= 12'h9ab;
        src91 <= 12'h9ca;
        src92 <= 12'h478;
        src93 <= 12'hc9d;
        src94 <= 12'ha81;
        src95 <= 12'h4c2;
        src96 <= 12'h86;
        src97 <= 12'hfae;
        src98 <= 12'h11e;
        src99 <= 12'h315;
        src100 <= 12'h234;
        src101 <= 12'h58;
        src102 <= 12'h811;
        src103 <= 12'hc32;
        src104 <= 12'h1d4;
        src105 <= 12'h657;
        src106 <= 12'h752;
        src107 <= 12'h89f;
        src108 <= 12'hf41;
        src109 <= 12'h8ad;
        src110 <= 12'h10a;
        src111 <= 12'hc4b;
        src112 <= 12'h75f;
        src113 <= 12'h6f5;
        src114 <= 12'h53c;
        src115 <= 12'hb01;
        src116 <= 12'ha30;
        src117 <= 12'hc4a;
        src118 <= 12'ha97;
        src119 <= 12'h7e;
        src120 <= 12'h77a;
        src121 <= 12'h2c9;
        src122 <= 12'h2da;
        src123 <= 12'h99d;
        src124 <= 12'h932;
        src125 <= 12'h7c1;
        src126 <= 12'he57;
        src127 <= 12'hc6;
        exp <= 19'h36b37;
        #1
        src0 <= 12'h2e3;
        src1 <= 12'hc89;
        src2 <= 12'h97d;
        src3 <= 12'hdab;
        src4 <= 12'hb83;
        src5 <= 12'he3a;
        src6 <= 12'hb7a;
        src7 <= 12'h2a9;
        src8 <= 12'h226;
        src9 <= 12'hf01;
        src10 <= 12'hc75;
        src11 <= 12'h521;
        src12 <= 12'h2;
        src13 <= 12'h1db;
        src14 <= 12'h4fa;
        src15 <= 12'hb8b;
        src16 <= 12'ha4a;
        src17 <= 12'h704;
        src18 <= 12'h376;
        src19 <= 12'h449;
        src20 <= 12'h2e;
        src21 <= 12'h50e;
        src22 <= 12'hd0a;
        src23 <= 12'hbe0;
        src24 <= 12'hf76;
        src25 <= 12'heb7;
        src26 <= 12'h367;
        src27 <= 12'hd8c;
        src28 <= 12'hfc0;
        src29 <= 12'hf1a;
        src30 <= 12'hf5;
        src31 <= 12'hded;
        src32 <= 12'hd3c;
        src33 <= 12'h33d;
        src34 <= 12'h78e;
        src35 <= 12'h5e6;
        src36 <= 12'h327;
        src37 <= 12'ha6f;
        src38 <= 12'hae;
        src39 <= 12'h4a3;
        src40 <= 12'h49;
        src41 <= 12'h573;
        src42 <= 12'h89a;
        src43 <= 12'h228;
        src44 <= 12'h91b;
        src45 <= 12'hf17;
        src46 <= 12'h5ca;
        src47 <= 12'hc3b;
        src48 <= 12'hd8c;
        src49 <= 12'hde6;
        src50 <= 12'h362;
        src51 <= 12'hd8b;
        src52 <= 12'hf9e;
        src53 <= 12'hc1;
        src54 <= 12'h9ec;
        src55 <= 12'h5d4;
        src56 <= 12'hb1f;
        src57 <= 12'ha01;
        src58 <= 12'h857;
        src59 <= 12'h6ec;
        src60 <= 12'h497;
        src61 <= 12'ha60;
        src62 <= 12'hafa;
        src63 <= 12'h835;
        src64 <= 12'h450;
        src65 <= 12'h86f;
        src66 <= 12'hb5b;
        src67 <= 12'h475;
        src68 <= 12'h2c9;
        src69 <= 12'h125;
        src70 <= 12'h164;
        src71 <= 12'h526;
        src72 <= 12'h806;
        src73 <= 12'h60f;
        src74 <= 12'h9d7;
        src75 <= 12'hfcc;
        src76 <= 12'ha8b;
        src77 <= 12'h30;
        src78 <= 12'hec0;
        src79 <= 12'hc1d;
        src80 <= 12'h48e;
        src81 <= 12'hcb0;
        src82 <= 12'h4ac;
        src83 <= 12'h50b;
        src84 <= 12'h5cb;
        src85 <= 12'h8c7;
        src86 <= 12'h6ca;
        src87 <= 12'haef;
        src88 <= 12'h9dc;
        src89 <= 12'h8b7;
        src90 <= 12'h490;
        src91 <= 12'hb0c;
        src92 <= 12'h505;
        src93 <= 12'h777;
        src94 <= 12'hf2f;
        src95 <= 12'h183;
        src96 <= 12'hf9a;
        src97 <= 12'h85;
        src98 <= 12'h292;
        src99 <= 12'he9f;
        src100 <= 12'hefd;
        src101 <= 12'h140;
        src102 <= 12'h14c;
        src103 <= 12'h93e;
        src104 <= 12'hb4e;
        src105 <= 12'h69c;
        src106 <= 12'h289;
        src107 <= 12'hb16;
        src108 <= 12'h36a;
        src109 <= 12'he30;
        src110 <= 12'hdb5;
        src111 <= 12'h64b;
        src112 <= 12'hcd0;
        src113 <= 12'he6c;
        src114 <= 12'he5b;
        src115 <= 12'h7a8;
        src116 <= 12'hd66;
        src117 <= 12'h658;
        src118 <= 12'hdc0;
        src119 <= 12'h9cc;
        src120 <= 12'h46d;
        src121 <= 12'hdd7;
        src122 <= 12'hdb1;
        src123 <= 12'h5d8;
        src124 <= 12'h36;
        src125 <= 12'h1cb;
        src126 <= 12'hdc8;
        src127 <= 12'h1b4;
        exp <= 19'h41a33;
        #1
        src0 <= 12'he52;
        src1 <= 12'h938;
        src2 <= 12'hd66;
        src3 <= 12'h93d;
        src4 <= 12'h7e2;
        src5 <= 12'h158;
        src6 <= 12'h763;
        src7 <= 12'haf;
        src8 <= 12'hcfd;
        src9 <= 12'hd49;
        src10 <= 12'h21c;
        src11 <= 12'h403;
        src12 <= 12'ha10;
        src13 <= 12'haec;
        src14 <= 12'h1e;
        src15 <= 12'hff2;
        src16 <= 12'h92e;
        src17 <= 12'hbb;
        src18 <= 12'hd41;
        src19 <= 12'hf41;
        src20 <= 12'hd10;
        src21 <= 12'hcd3;
        src22 <= 12'hf82;
        src23 <= 12'hea6;
        src24 <= 12'h90b;
        src25 <= 12'h7d4;
        src26 <= 12'hc80;
        src27 <= 12'h92d;
        src28 <= 12'hc92;
        src29 <= 12'hc0a;
        src30 <= 12'ha41;
        src31 <= 12'h955;
        src32 <= 12'h91d;
        src33 <= 12'h346;
        src34 <= 12'hfe;
        src35 <= 12'h9da;
        src36 <= 12'hb74;
        src37 <= 12'h6c;
        src38 <= 12'h81d;
        src39 <= 12'h14e;
        src40 <= 12'h38;
        src41 <= 12'h33e;
        src42 <= 12'hba9;
        src43 <= 12'ha1b;
        src44 <= 12'hfec;
        src45 <= 12'hcff;
        src46 <= 12'h31c;
        src47 <= 12'h9f6;
        src48 <= 12'h8f9;
        src49 <= 12'h3e9;
        src50 <= 12'h9e8;
        src51 <= 12'h3f0;
        src52 <= 12'hb7b;
        src53 <= 12'h279;
        src54 <= 12'h6a7;
        src55 <= 12'hf2a;
        src56 <= 12'hb91;
        src57 <= 12'hd7d;
        src58 <= 12'h8be;
        src59 <= 12'h2f1;
        src60 <= 12'h930;
        src61 <= 12'h1bc;
        src62 <= 12'h3a4;
        src63 <= 12'h4fe;
        src64 <= 12'hd76;
        src65 <= 12'h6b4;
        src66 <= 12'he8e;
        src67 <= 12'h3de;
        src68 <= 12'hbec;
        src69 <= 12'h1;
        src70 <= 12'h13f;
        src71 <= 12'h428;
        src72 <= 12'hb5e;
        src73 <= 12'h312;
        src74 <= 12'hb1a;
        src75 <= 12'hd8a;
        src76 <= 12'h395;
        src77 <= 12'hb1c;
        src78 <= 12'h526;
        src79 <= 12'h905;
        src80 <= 12'hd08;
        src81 <= 12'h6dc;
        src82 <= 12'h305;
        src83 <= 12'h800;
        src84 <= 12'h3b0;
        src85 <= 12'he44;
        src86 <= 12'he;
        src87 <= 12'hb54;
        src88 <= 12'hd3a;
        src89 <= 12'he4b;
        src90 <= 12'h117;
        src91 <= 12'ha48;
        src92 <= 12'hab1;
        src93 <= 12'h808;
        src94 <= 12'h35c;
        src95 <= 12'ha3f;
        src96 <= 12'h687;
        src97 <= 12'h583;
        src98 <= 12'hc58;
        src99 <= 12'h21f;
        src100 <= 12'h95d;
        src101 <= 12'hd4f;
        src102 <= 12'hfd4;
        src103 <= 12'hc76;
        src104 <= 12'ha73;
        src105 <= 12'h90b;
        src106 <= 12'h151;
        src107 <= 12'hbca;
        src108 <= 12'ha1e;
        src109 <= 12'h701;
        src110 <= 12'hba6;
        src111 <= 12'hc8;
        src112 <= 12'h4e0;
        src113 <= 12'h5f0;
        src114 <= 12'h66e;
        src115 <= 12'h540;
        src116 <= 12'h8d6;
        src117 <= 12'hfd9;
        src118 <= 12'h10e;
        src119 <= 12'ha3f;
        src120 <= 12'hb81;
        src121 <= 12'h4aa;
        src122 <= 12'hcb;
        src123 <= 12'hed1;
        src124 <= 12'hf90;
        src125 <= 12'hffc;
        src126 <= 12'he74;
        src127 <= 12'h2bc;
        exp <= 19'h43290;
        #1
        src0 <= 12'h176;
        src1 <= 12'h6b0;
        src2 <= 12'hc68;
        src3 <= 12'hd9d;
        src4 <= 12'hc00;
        src5 <= 12'h237;
        src6 <= 12'hc4a;
        src7 <= 12'h575;
        src8 <= 12'hfb4;
        src9 <= 12'h633;
        src10 <= 12'h66e;
        src11 <= 12'h530;
        src12 <= 12'h787;
        src13 <= 12'hca8;
        src14 <= 12'hf1d;
        src15 <= 12'h8d0;
        src16 <= 12'ha9c;
        src17 <= 12'hf57;
        src18 <= 12'h6d2;
        src19 <= 12'h178;
        src20 <= 12'h557;
        src21 <= 12'h153;
        src22 <= 12'hdcc;
        src23 <= 12'h572;
        src24 <= 12'h32c;
        src25 <= 12'h45a;
        src26 <= 12'h4a;
        src27 <= 12'h3ab;
        src28 <= 12'heeb;
        src29 <= 12'hf1f;
        src30 <= 12'h8be;
        src31 <= 12'hbba;
        src32 <= 12'h940;
        src33 <= 12'h47d;
        src34 <= 12'hecc;
        src35 <= 12'h4ef;
        src36 <= 12'h4a0;
        src37 <= 12'h970;
        src38 <= 12'ha88;
        src39 <= 12'h407;
        src40 <= 12'h50d;
        src41 <= 12'h385;
        src42 <= 12'h749;
        src43 <= 12'h8e0;
        src44 <= 12'h2a2;
        src45 <= 12'he77;
        src46 <= 12'h219;
        src47 <= 12'h980;
        src48 <= 12'hbab;
        src49 <= 12'h568;
        src50 <= 12'hfa3;
        src51 <= 12'h387;
        src52 <= 12'h1a8;
        src53 <= 12'hfb4;
        src54 <= 12'h95a;
        src55 <= 12'hdb3;
        src56 <= 12'h151;
        src57 <= 12'h4e6;
        src58 <= 12'h7c0;
        src59 <= 12'h9ba;
        src60 <= 12'h75f;
        src61 <= 12'h822;
        src62 <= 12'hce5;
        src63 <= 12'hb8a;
        src64 <= 12'hfb6;
        src65 <= 12'h1f9;
        src66 <= 12'h53a;
        src67 <= 12'hc7d;
        src68 <= 12'h393;
        src69 <= 12'h9a0;
        src70 <= 12'h8cf;
        src71 <= 12'h8fa;
        src72 <= 12'hc17;
        src73 <= 12'h909;
        src74 <= 12'h526;
        src75 <= 12'hb8f;
        src76 <= 12'h120;
        src77 <= 12'he77;
        src78 <= 12'he5d;
        src79 <= 12'h701;
        src80 <= 12'h726;
        src81 <= 12'h540;
        src82 <= 12'hd31;
        src83 <= 12'hcc2;
        src84 <= 12'hae1;
        src85 <= 12'ha9b;
        src86 <= 12'hfe8;
        src87 <= 12'h56e;
        src88 <= 12'h472;
        src89 <= 12'hb19;
        src90 <= 12'h186;
        src91 <= 12'hb8c;
        src92 <= 12'h634;
        src93 <= 12'h6a7;
        src94 <= 12'h830;
        src95 <= 12'h257;
        src96 <= 12'h6f0;
        src97 <= 12'hb59;
        src98 <= 12'h5e1;
        src99 <= 12'had;
        src100 <= 12'h83a;
        src101 <= 12'hb4a;
        src102 <= 12'h33e;
        src103 <= 12'h7d7;
        src104 <= 12'h740;
        src105 <= 12'h1f7;
        src106 <= 12'h6e5;
        src107 <= 12'haa;
        src108 <= 12'h16;
        src109 <= 12'h69a;
        src110 <= 12'hc08;
        src111 <= 12'he5f;
        src112 <= 12'h4fc;
        src113 <= 12'h813;
        src114 <= 12'haaa;
        src115 <= 12'h773;
        src116 <= 12'h1c;
        src117 <= 12'h91c;
        src118 <= 12'h243;
        src119 <= 12'h9d5;
        src120 <= 12'h436;
        src121 <= 12'h9c4;
        src122 <= 12'hecf;
        src123 <= 12'haa3;
        src124 <= 12'h3b4;
        src125 <= 12'h95;
        src126 <= 12'h7c2;
        src127 <= 12'h680;
        exp <= 19'h3f3c5;
        #1
        src0 <= 12'hb72;
        src1 <= 12'h1d4;
        src2 <= 12'hc8f;
        src3 <= 12'he0f;
        src4 <= 12'hb8c;
        src5 <= 12'h5bf;
        src6 <= 12'hfe;
        src7 <= 12'h876;
        src8 <= 12'h692;
        src9 <= 12'hcbd;
        src10 <= 12'h419;
        src11 <= 12'hc5e;
        src12 <= 12'h4bc;
        src13 <= 12'hc90;
        src14 <= 12'hae0;
        src15 <= 12'ha43;
        src16 <= 12'h26c;
        src17 <= 12'h91f;
        src18 <= 12'hc8a;
        src19 <= 12'hc14;
        src20 <= 12'h87f;
        src21 <= 12'hdbb;
        src22 <= 12'h364;
        src23 <= 12'h4d8;
        src24 <= 12'h143;
        src25 <= 12'hc6a;
        src26 <= 12'h15f;
        src27 <= 12'h6e5;
        src28 <= 12'hb95;
        src29 <= 12'h9d6;
        src30 <= 12'h8dc;
        src31 <= 12'h94c;
        src32 <= 12'h6f1;
        src33 <= 12'h17f;
        src34 <= 12'h22b;
        src35 <= 12'h499;
        src36 <= 12'h262;
        src37 <= 12'h7bd;
        src38 <= 12'h4e3;
        src39 <= 12'h66f;
        src40 <= 12'h51d;
        src41 <= 12'h4f9;
        src42 <= 12'hdee;
        src43 <= 12'hd7b;
        src44 <= 12'h7c4;
        src45 <= 12'h8f4;
        src46 <= 12'hdc4;
        src47 <= 12'hc2;
        src48 <= 12'hf54;
        src49 <= 12'h101;
        src50 <= 12'h5f1;
        src51 <= 12'h47a;
        src52 <= 12'hd9e;
        src53 <= 12'hdeb;
        src54 <= 12'hb1e;
        src55 <= 12'hd11;
        src56 <= 12'h8f4;
        src57 <= 12'h43;
        src58 <= 12'h706;
        src59 <= 12'h241;
        src60 <= 12'hab6;
        src61 <= 12'heae;
        src62 <= 12'hc2a;
        src63 <= 12'h20;
        src64 <= 12'h217;
        src65 <= 12'haa2;
        src66 <= 12'h2f3;
        src67 <= 12'h8ab;
        src68 <= 12'hed1;
        src69 <= 12'h367;
        src70 <= 12'h8a4;
        src71 <= 12'hcc5;
        src72 <= 12'he38;
        src73 <= 12'hf9c;
        src74 <= 12'h9f4;
        src75 <= 12'h7d3;
        src76 <= 12'h950;
        src77 <= 12'h2c6;
        src78 <= 12'h6a0;
        src79 <= 12'ha97;
        src80 <= 12'hcf4;
        src81 <= 12'he12;
        src82 <= 12'h929;
        src83 <= 12'h1b6;
        src84 <= 12'h619;
        src85 <= 12'had3;
        src86 <= 12'hc63;
        src87 <= 12'hcb4;
        src88 <= 12'h2dc;
        src89 <= 12'h5f1;
        src90 <= 12'h394;
        src91 <= 12'h93a;
        src92 <= 12'h98f;
        src93 <= 12'h38a;
        src94 <= 12'ha50;
        src95 <= 12'hd11;
        src96 <= 12'hfd7;
        src97 <= 12'h74b;
        src98 <= 12'hcfc;
        src99 <= 12'h2e7;
        src100 <= 12'h79a;
        src101 <= 12'h1e3;
        src102 <= 12'haff;
        src103 <= 12'h4d;
        src104 <= 12'haf7;
        src105 <= 12'h831;
        src106 <= 12'h60a;
        src107 <= 12'h6ba;
        src108 <= 12'hf4c;
        src109 <= 12'h3ae;
        src110 <= 12'h70;
        src111 <= 12'h315;
        src112 <= 12'h3;
        src113 <= 12'hccc;
        src114 <= 12'h146;
        src115 <= 12'h633;
        src116 <= 12'hfc3;
        src117 <= 12'h2db;
        src118 <= 12'h66a;
        src119 <= 12'h93;
        src120 <= 12'ha7b;
        src121 <= 12'hedd;
        src122 <= 12'h262;
        src123 <= 12'h831;
        src124 <= 12'h503;
        src125 <= 12'h738;
        src126 <= 12'hec5;
        src127 <= 12'h512;
        exp <= 19'h3f7f7;
        #1
        src0 <= 12'hbd3;
        src1 <= 12'hd8d;
        src2 <= 12'h220;
        src3 <= 12'hc3;
        src4 <= 12'h4d9;
        src5 <= 12'h6f1;
        src6 <= 12'h885;
        src7 <= 12'hc89;
        src8 <= 12'habd;
        src9 <= 12'h6d6;
        src10 <= 12'ha3c;
        src11 <= 12'hfcf;
        src12 <= 12'h8fd;
        src13 <= 12'hf05;
        src14 <= 12'hf9f;
        src15 <= 12'hd1c;
        src16 <= 12'h4ca;
        src17 <= 12'h47a;
        src18 <= 12'hac5;
        src19 <= 12'h8c9;
        src20 <= 12'hc4e;
        src21 <= 12'h75c;
        src22 <= 12'hdf9;
        src23 <= 12'h8b2;
        src24 <= 12'h782;
        src25 <= 12'h494;
        src26 <= 12'h66e;
        src27 <= 12'h940;
        src28 <= 12'h50a;
        src29 <= 12'hfa8;
        src30 <= 12'hb6;
        src31 <= 12'h408;
        src32 <= 12'hbd9;
        src33 <= 12'h467;
        src34 <= 12'h78f;
        src35 <= 12'ha23;
        src36 <= 12'h418;
        src37 <= 12'h3e2;
        src38 <= 12'h9fd;
        src39 <= 12'h74f;
        src40 <= 12'hdfe;
        src41 <= 12'hdd3;
        src42 <= 12'h2ab;
        src43 <= 12'heb2;
        src44 <= 12'hd72;
        src45 <= 12'h6da;
        src46 <= 12'h94e;
        src47 <= 12'h24c;
        src48 <= 12'h116;
        src49 <= 12'h47;
        src50 <= 12'hafc;
        src51 <= 12'h59e;
        src52 <= 12'h40e;
        src53 <= 12'h1e7;
        src54 <= 12'h30f;
        src55 <= 12'h9f1;
        src56 <= 12'h222;
        src57 <= 12'hceb;
        src58 <= 12'h41f;
        src59 <= 12'hc08;
        src60 <= 12'he89;
        src61 <= 12'h903;
        src62 <= 12'hec;
        src63 <= 12'h418;
        src64 <= 12'hcbd;
        src65 <= 12'h2f;
        src66 <= 12'h73;
        src67 <= 12'hce5;
        src68 <= 12'h7ab;
        src69 <= 12'h917;
        src70 <= 12'h9a3;
        src71 <= 12'hafc;
        src72 <= 12'hf11;
        src73 <= 12'h74d;
        src74 <= 12'h292;
        src75 <= 12'hb89;
        src76 <= 12'hc4b;
        src77 <= 12'he7c;
        src78 <= 12'h4c;
        src79 <= 12'h9c5;
        src80 <= 12'hf96;
        src81 <= 12'h347;
        src82 <= 12'h5ce;
        src83 <= 12'heb8;
        src84 <= 12'he6b;
        src85 <= 12'hc0f;
        src86 <= 12'hd73;
        src87 <= 12'h1c0;
        src88 <= 12'hdc0;
        src89 <= 12'hb98;
        src90 <= 12'he0d;
        src91 <= 12'h625;
        src92 <= 12'hed4;
        src93 <= 12'h62c;
        src94 <= 12'h24d;
        src95 <= 12'h5ea;
        src96 <= 12'hf84;
        src97 <= 12'he77;
        src98 <= 12'h841;
        src99 <= 12'hf5f;
        src100 <= 12'h79e;
        src101 <= 12'ha35;
        src102 <= 12'h53c;
        src103 <= 12'h4cd;
        src104 <= 12'h838;
        src105 <= 12'h875;
        src106 <= 12'h49d;
        src107 <= 12'h379;
        src108 <= 12'hf5d;
        src109 <= 12'h2b2;
        src110 <= 12'hb41;
        src111 <= 12'h1d9;
        src112 <= 12'hb02;
        src113 <= 12'had8;
        src114 <= 12'hb08;
        src115 <= 12'h3a5;
        src116 <= 12'hf09;
        src117 <= 12'he78;
        src118 <= 12'h277;
        src119 <= 12'h45;
        src120 <= 12'hcfc;
        src121 <= 12'h7b4;
        src122 <= 12'h3c3;
        src123 <= 12'hd79;
        src124 <= 12'hf82;
        src125 <= 12'h5cb;
        src126 <= 12'hf1b;
        src127 <= 12'h8a1;
        exp <= 19'h448b0;
        #1
        src0 <= 12'h74a;
        src1 <= 12'h881;
        src2 <= 12'h8ba;
        src3 <= 12'h71d;
        src4 <= 12'h4c9;
        src5 <= 12'hd5b;
        src6 <= 12'hf29;
        src7 <= 12'hce5;
        src8 <= 12'hd0a;
        src9 <= 12'hdc8;
        src10 <= 12'hd2b;
        src11 <= 12'h395;
        src12 <= 12'hd13;
        src13 <= 12'hcf1;
        src14 <= 12'h61d;
        src15 <= 12'h597;
        src16 <= 12'ha69;
        src17 <= 12'h68a;
        src18 <= 12'h76b;
        src19 <= 12'hd90;
        src20 <= 12'h49;
        src21 <= 12'hc07;
        src22 <= 12'h7f3;
        src23 <= 12'hb7c;
        src24 <= 12'hd85;
        src25 <= 12'ha6e;
        src26 <= 12'h514;
        src27 <= 12'hb5b;
        src28 <= 12'hf76;
        src29 <= 12'h64c;
        src30 <= 12'h5c9;
        src31 <= 12'h1e6;
        src32 <= 12'hebe;
        src33 <= 12'h113;
        src34 <= 12'h4c6;
        src35 <= 12'hbcf;
        src36 <= 12'h6c4;
        src37 <= 12'hac4;
        src38 <= 12'hfb0;
        src39 <= 12'ha26;
        src40 <= 12'hba0;
        src41 <= 12'h2e3;
        src42 <= 12'h392;
        src43 <= 12'h173;
        src44 <= 12'hb42;
        src45 <= 12'h4c3;
        src46 <= 12'h1a1;
        src47 <= 12'hdbd;
        src48 <= 12'ha37;
        src49 <= 12'hd54;
        src50 <= 12'hda2;
        src51 <= 12'hc51;
        src52 <= 12'h25b;
        src53 <= 12'h5d8;
        src54 <= 12'ha32;
        src55 <= 12'h323;
        src56 <= 12'h265;
        src57 <= 12'hd0;
        src58 <= 12'h706;
        src59 <= 12'h284;
        src60 <= 12'he2d;
        src61 <= 12'h404;
        src62 <= 12'h5f4;
        src63 <= 12'h934;
        src64 <= 12'h4bd;
        src65 <= 12'hcd1;
        src66 <= 12'h5c1;
        src67 <= 12'hf89;
        src68 <= 12'h21a;
        src69 <= 12'hd96;
        src70 <= 12'h197;
        src71 <= 12'ha45;
        src72 <= 12'h9c6;
        src73 <= 12'h171;
        src74 <= 12'h4c;
        src75 <= 12'h1be;
        src76 <= 12'h40c;
        src77 <= 12'had2;
        src78 <= 12'h74f;
        src79 <= 12'h112;
        src80 <= 12'hebb;
        src81 <= 12'hbe3;
        src82 <= 12'h8e2;
        src83 <= 12'h675;
        src84 <= 12'h902;
        src85 <= 12'hd91;
        src86 <= 12'h813;
        src87 <= 12'h3ee;
        src88 <= 12'h1db;
        src89 <= 12'h199;
        src90 <= 12'h2cf;
        src91 <= 12'hc20;
        src92 <= 12'hee5;
        src93 <= 12'hb5d;
        src94 <= 12'hb05;
        src95 <= 12'hd2e;
        src96 <= 12'h4df;
        src97 <= 12'hccd;
        src98 <= 12'h748;
        src99 <= 12'h245;
        src100 <= 12'h74f;
        src101 <= 12'hb74;
        src102 <= 12'heba;
        src103 <= 12'h1;
        src104 <= 12'h97b;
        src105 <= 12'h25b;
        src106 <= 12'hf1b;
        src107 <= 12'h8e3;
        src108 <= 12'h62c;
        src109 <= 12'he94;
        src110 <= 12'hbf6;
        src111 <= 12'h430;
        src112 <= 12'hb21;
        src113 <= 12'he10;
        src114 <= 12'h51b;
        src115 <= 12'ha03;
        src116 <= 12'hcc7;
        src117 <= 12'h604;
        src118 <= 12'hbb3;
        src119 <= 12'h5e1;
        src120 <= 12'h85e;
        src121 <= 12'haae;
        src122 <= 12'h339;
        src123 <= 12'hd8d;
        src124 <= 12'h280;
        src125 <= 12'h21;
        src126 <= 12'he52;
        src127 <= 12'h8aa;
        exp <= 19'h4263e;
        #1
        src0 <= 12'h394;
        src1 <= 12'h9f9;
        src2 <= 12'ha69;
        src3 <= 12'haf6;
        src4 <= 12'h1ed;
        src5 <= 12'h685;
        src6 <= 12'h375;
        src7 <= 12'hb75;
        src8 <= 12'he9;
        src9 <= 12'h100;
        src10 <= 12'h5b8;
        src11 <= 12'h9b4;
        src12 <= 12'h438;
        src13 <= 12'h7d2;
        src14 <= 12'h669;
        src15 <= 12'h752;
        src16 <= 12'h44d;
        src17 <= 12'h2af;
        src18 <= 12'h7cc;
        src19 <= 12'hfd5;
        src20 <= 12'h624;
        src21 <= 12'he5f;
        src22 <= 12'hade;
        src23 <= 12'haa2;
        src24 <= 12'ha07;
        src25 <= 12'hab4;
        src26 <= 12'h483;
        src27 <= 12'h15;
        src28 <= 12'h5f6;
        src29 <= 12'h763;
        src30 <= 12'h49a;
        src31 <= 12'h145;
        src32 <= 12'h615;
        src33 <= 12'h86c;
        src34 <= 12'h8ac;
        src35 <= 12'h218;
        src36 <= 12'h784;
        src37 <= 12'h7e9;
        src38 <= 12'hf66;
        src39 <= 12'hb0b;
        src40 <= 12'hfc9;
        src41 <= 12'h40c;
        src42 <= 12'h5fe;
        src43 <= 12'hfa6;
        src44 <= 12'h168;
        src45 <= 12'had7;
        src46 <= 12'h66e;
        src47 <= 12'habf;
        src48 <= 12'h410;
        src49 <= 12'he08;
        src50 <= 12'h4f6;
        src51 <= 12'h561;
        src52 <= 12'h38b;
        src53 <= 12'h747;
        src54 <= 12'h560;
        src55 <= 12'h635;
        src56 <= 12'hdc6;
        src57 <= 12'ha5d;
        src58 <= 12'ha42;
        src59 <= 12'h768;
        src60 <= 12'hd06;
        src61 <= 12'h218;
        src62 <= 12'h6a4;
        src63 <= 12'h22a;
        src64 <= 12'h99d;
        src65 <= 12'hd50;
        src66 <= 12'h653;
        src67 <= 12'h555;
        src68 <= 12'h8eb;
        src69 <= 12'h87b;
        src70 <= 12'hdcb;
        src71 <= 12'hd79;
        src72 <= 12'h9e4;
        src73 <= 12'h6d1;
        src74 <= 12'h990;
        src75 <= 12'h499;
        src76 <= 12'h1f0;
        src77 <= 12'h459;
        src78 <= 12'h6f7;
        src79 <= 12'hd9f;
        src80 <= 12'he1c;
        src81 <= 12'h9b1;
        src82 <= 12'h427;
        src83 <= 12'h77e;
        src84 <= 12'h53f;
        src85 <= 12'hcfc;
        src86 <= 12'h3ba;
        src87 <= 12'h59;
        src88 <= 12'he5e;
        src89 <= 12'h55d;
        src90 <= 12'hf0a;
        src91 <= 12'hf79;
        src92 <= 12'h89d;
        src93 <= 12'hb11;
        src94 <= 12'h765;
        src95 <= 12'h756;
        src96 <= 12'h778;
        src97 <= 12'hefa;
        src98 <= 12'hb8;
        src99 <= 12'h67e;
        src100 <= 12'hd2;
        src101 <= 12'h724;
        src102 <= 12'h3ab;
        src103 <= 12'h17f;
        src104 <= 12'h88;
        src105 <= 12'h21b;
        src106 <= 12'hf48;
        src107 <= 12'h50a;
        src108 <= 12'h9d9;
        src109 <= 12'h33c;
        src110 <= 12'h3b;
        src111 <= 12'hcdc;
        src112 <= 12'hb4;
        src113 <= 12'h6d8;
        src114 <= 12'hd00;
        src115 <= 12'h281;
        src116 <= 12'h2ff;
        src117 <= 12'ha9f;
        src118 <= 12'h478;
        src119 <= 12'h543;
        src120 <= 12'h46;
        src121 <= 12'ha78;
        src122 <= 12'ha7c;
        src123 <= 12'h91b;
        src124 <= 12'hbb4;
        src125 <= 12'h56f;
        src126 <= 12'h15e;
        src127 <= 12'h137;
        exp <= 19'h3ace3;
        #1
        src0 <= 12'h8e6;
        src1 <= 12'h70e;
        src2 <= 12'h604;
        src3 <= 12'h96e;
        src4 <= 12'ha54;
        src5 <= 12'h876;
        src6 <= 12'h8db;
        src7 <= 12'h1c7;
        src8 <= 12'h454;
        src9 <= 12'hbf1;
        src10 <= 12'h460;
        src11 <= 12'hd51;
        src12 <= 12'h6c8;
        src13 <= 12'h90;
        src14 <= 12'he21;
        src15 <= 12'hd1e;
        src16 <= 12'h259;
        src17 <= 12'h3f4;
        src18 <= 12'hc2f;
        src19 <= 12'hca;
        src20 <= 12'hd00;
        src21 <= 12'h94a;
        src22 <= 12'h6e9;
        src23 <= 12'h920;
        src24 <= 12'hb78;
        src25 <= 12'h65e;
        src26 <= 12'h50;
        src27 <= 12'h34e;
        src28 <= 12'hfe8;
        src29 <= 12'h640;
        src30 <= 12'h37e;
        src31 <= 12'hf7f;
        src32 <= 12'h85e;
        src33 <= 12'he42;
        src34 <= 12'h84b;
        src35 <= 12'h549;
        src36 <= 12'h86e;
        src37 <= 12'ha19;
        src38 <= 12'h50e;
        src39 <= 12'h5d7;
        src40 <= 12'h4d4;
        src41 <= 12'hf97;
        src42 <= 12'he7f;
        src43 <= 12'h899;
        src44 <= 12'hf53;
        src45 <= 12'h260;
        src46 <= 12'head;
        src47 <= 12'he8d;
        src48 <= 12'ha9c;
        src49 <= 12'h8be;
        src50 <= 12'h1bc;
        src51 <= 12'hf2c;
        src52 <= 12'h873;
        src53 <= 12'h348;
        src54 <= 12'h360;
        src55 <= 12'hf60;
        src56 <= 12'h46a;
        src57 <= 12'hfc7;
        src58 <= 12'h283;
        src59 <= 12'h970;
        src60 <= 12'hbc4;
        src61 <= 12'hc35;
        src62 <= 12'hb85;
        src63 <= 12'hffb;
        src64 <= 12'hce9;
        src65 <= 12'h5b;
        src66 <= 12'hb06;
        src67 <= 12'hd21;
        src68 <= 12'hdc1;
        src69 <= 12'hc54;
        src70 <= 12'h52a;
        src71 <= 12'h799;
        src72 <= 12'hab2;
        src73 <= 12'h5c7;
        src74 <= 12'h654;
        src75 <= 12'h81f;
        src76 <= 12'ha78;
        src77 <= 12'h36e;
        src78 <= 12'h48a;
        src79 <= 12'h3d5;
        src80 <= 12'hc08;
        src81 <= 12'h1e5;
        src82 <= 12'h5f4;
        src83 <= 12'hc86;
        src84 <= 12'hb8e;
        src85 <= 12'h615;
        src86 <= 12'h1ea;
        src87 <= 12'h888;
        src88 <= 12'h994;
        src89 <= 12'h20;
        src90 <= 12'he03;
        src91 <= 12'h78d;
        src92 <= 12'hc15;
        src93 <= 12'h7b6;
        src94 <= 12'h1d5;
        src95 <= 12'h330;
        src96 <= 12'hc76;
        src97 <= 12'h96c;
        src98 <= 12'hfc8;
        src99 <= 12'h28a;
        src100 <= 12'h146;
        src101 <= 12'h5b7;
        src102 <= 12'h8b6;
        src103 <= 12'h4de;
        src104 <= 12'hffb;
        src105 <= 12'h40d;
        src106 <= 12'hca1;
        src107 <= 12'hb62;
        src108 <= 12'hcd5;
        src109 <= 12'hb23;
        src110 <= 12'h853;
        src111 <= 12'hb21;
        src112 <= 12'h275;
        src113 <= 12'he6d;
        src114 <= 12'hd76;
        src115 <= 12'hac0;
        src116 <= 12'hb43;
        src117 <= 12'he88;
        src118 <= 12'h33d;
        src119 <= 12'ha42;
        src120 <= 12'h26a;
        src121 <= 12'hc8c;
        src122 <= 12'h58b;
        src123 <= 12'h961;
        src124 <= 12'h114;
        src125 <= 12'h110;
        src126 <= 12'h30b;
        src127 <= 12'h32f;
        exp <= 19'h42cdd;
        #1
        src0 <= 12'hf5;
        src1 <= 12'h903;
        src2 <= 12'h526;
        src3 <= 12'hdfb;
        src4 <= 12'h724;
        src5 <= 12'hde5;
        src6 <= 12'h7c1;
        src7 <= 12'he81;
        src8 <= 12'h959;
        src9 <= 12'ha5f;
        src10 <= 12'h160;
        src11 <= 12'hdf2;
        src12 <= 12'h689;
        src13 <= 12'h271;
        src14 <= 12'h92c;
        src15 <= 12'h7a9;
        src16 <= 12'h6a;
        src17 <= 12'h63;
        src18 <= 12'h82c;
        src19 <= 12'hb2a;
        src20 <= 12'h13d;
        src21 <= 12'ha08;
        src22 <= 12'h11f;
        src23 <= 12'h123;
        src24 <= 12'h2e6;
        src25 <= 12'h971;
        src26 <= 12'hf92;
        src27 <= 12'h58c;
        src28 <= 12'h94a;
        src29 <= 12'hf1;
        src30 <= 12'h88a;
        src31 <= 12'hd46;
        src32 <= 12'h33;
        src33 <= 12'h32f;
        src34 <= 12'h794;
        src35 <= 12'h46;
        src36 <= 12'h4fc;
        src37 <= 12'h587;
        src38 <= 12'h95d;
        src39 <= 12'he2a;
        src40 <= 12'h148;
        src41 <= 12'hff0;
        src42 <= 12'hbd8;
        src43 <= 12'hd0b;
        src44 <= 12'h84c;
        src45 <= 12'hea1;
        src46 <= 12'h7da;
        src47 <= 12'hd5d;
        src48 <= 12'h54a;
        src49 <= 12'haa0;
        src50 <= 12'h958;
        src51 <= 12'h60;
        src52 <= 12'hb80;
        src53 <= 12'h20a;
        src54 <= 12'h853;
        src55 <= 12'h1ff;
        src56 <= 12'h15c;
        src57 <= 12'h84;
        src58 <= 12'h9c7;
        src59 <= 12'hae6;
        src60 <= 12'hd27;
        src61 <= 12'h137;
        src62 <= 12'h716;
        src63 <= 12'hf76;
        src64 <= 12'h4d7;
        src65 <= 12'h614;
        src66 <= 12'h835;
        src67 <= 12'hb96;
        src68 <= 12'he45;
        src69 <= 12'hba1;
        src70 <= 12'h43f;
        src71 <= 12'hee1;
        src72 <= 12'hf13;
        src73 <= 12'h33d;
        src74 <= 12'h641;
        src75 <= 12'h853;
        src76 <= 12'h299;
        src77 <= 12'hc0d;
        src78 <= 12'hb59;
        src79 <= 12'h9e5;
        src80 <= 12'ha9a;
        src81 <= 12'h34a;
        src82 <= 12'h6aa;
        src83 <= 12'h71c;
        src84 <= 12'h87;
        src85 <= 12'hcd3;
        src86 <= 12'h6eb;
        src87 <= 12'hebe;
        src88 <= 12'h784;
        src89 <= 12'h8d2;
        src90 <= 12'h6cb;
        src91 <= 12'h76c;
        src92 <= 12'hf50;
        src93 <= 12'hba2;
        src94 <= 12'h2f7;
        src95 <= 12'h9b7;
        src96 <= 12'h9fc;
        src97 <= 12'h495;
        src98 <= 12'h7f0;
        src99 <= 12'h910;
        src100 <= 12'h55b;
        src101 <= 12'h184;
        src102 <= 12'h66;
        src103 <= 12'ha0c;
        src104 <= 12'h47;
        src105 <= 12'ha24;
        src106 <= 12'hab9;
        src107 <= 12'h4de;
        src108 <= 12'hb02;
        src109 <= 12'h3eb;
        src110 <= 12'had9;
        src111 <= 12'heda;
        src112 <= 12'h22a;
        src113 <= 12'h309;
        src114 <= 12'h6aa;
        src115 <= 12'hb42;
        src116 <= 12'h106;
        src117 <= 12'h211;
        src118 <= 12'h334;
        src119 <= 12'h200;
        src120 <= 12'h63c;
        src121 <= 12'h7eb;
        src122 <= 12'h10a;
        src123 <= 12'h66c;
        src124 <= 12'hdb8;
        src125 <= 12'h850;
        src126 <= 12'he18;
        src127 <= 12'h3ab;
        exp <= 19'h3be95;
        #1
        src0 <= 12'h49d;
        src1 <= 12'h262;
        src2 <= 12'h53f;
        src3 <= 12'hc2a;
        src4 <= 12'h5f;
        src5 <= 12'hc60;
        src6 <= 12'hc7e;
        src7 <= 12'hddd;
        src8 <= 12'hf1f;
        src9 <= 12'h6b6;
        src10 <= 12'hd32;
        src11 <= 12'h646;
        src12 <= 12'h958;
        src13 <= 12'hd1d;
        src14 <= 12'h821;
        src15 <= 12'h81b;
        src16 <= 12'h326;
        src17 <= 12'hd0;
        src18 <= 12'hb32;
        src19 <= 12'hb9b;
        src20 <= 12'h889;
        src21 <= 12'h5a5;
        src22 <= 12'h5a5;
        src23 <= 12'h9b1;
        src24 <= 12'h995;
        src25 <= 12'h1fd;
        src26 <= 12'h710;
        src27 <= 12'h7b5;
        src28 <= 12'he6d;
        src29 <= 12'hd1b;
        src30 <= 12'hd7;
        src31 <= 12'he71;
        src32 <= 12'h3f8;
        src33 <= 12'h246;
        src34 <= 12'hbfb;
        src35 <= 12'h26;
        src36 <= 12'hc05;
        src37 <= 12'hd3b;
        src38 <= 12'h52e;
        src39 <= 12'h27d;
        src40 <= 12'hf12;
        src41 <= 12'h7cb;
        src42 <= 12'hee;
        src43 <= 12'h781;
        src44 <= 12'h750;
        src45 <= 12'hdef;
        src46 <= 12'h156;
        src47 <= 12'h8c7;
        src48 <= 12'hf24;
        src49 <= 12'hc5;
        src50 <= 12'h941;
        src51 <= 12'h149;
        src52 <= 12'h6be;
        src53 <= 12'h5d8;
        src54 <= 12'hfa8;
        src55 <= 12'hf;
        src56 <= 12'h39a;
        src57 <= 12'h4f6;
        src58 <= 12'hee1;
        src59 <= 12'h961;
        src60 <= 12'h630;
        src61 <= 12'h769;
        src62 <= 12'hb5d;
        src63 <= 12'h258;
        src64 <= 12'h9af;
        src65 <= 12'hca0;
        src66 <= 12'hdef;
        src67 <= 12'ha3b;
        src68 <= 12'h3bb;
        src69 <= 12'ha23;
        src70 <= 12'h1ea;
        src71 <= 12'he30;
        src72 <= 12'h126;
        src73 <= 12'hdc5;
        src74 <= 12'h4af;
        src75 <= 12'h187;
        src76 <= 12'h363;
        src77 <= 12'h1be;
        src78 <= 12'he37;
        src79 <= 12'hdde;
        src80 <= 12'h4c;
        src81 <= 12'h1a6;
        src82 <= 12'h2e7;
        src83 <= 12'hcbf;
        src84 <= 12'ha7;
        src85 <= 12'hc55;
        src86 <= 12'h6d7;
        src87 <= 12'hc12;
        src88 <= 12'h760;
        src89 <= 12'hbc9;
        src90 <= 12'hc83;
        src91 <= 12'h49e;
        src92 <= 12'ha54;
        src93 <= 12'h6d;
        src94 <= 12'h8c6;
        src95 <= 12'h621;
        src96 <= 12'hfb6;
        src97 <= 12'h1fd;
        src98 <= 12'he4c;
        src99 <= 12'h769;
        src100 <= 12'h72e;
        src101 <= 12'h9d9;
        src102 <= 12'h36d;
        src103 <= 12'h112;
        src104 <= 12'hc42;
        src105 <= 12'hb4;
        src106 <= 12'hcd;
        src107 <= 12'he48;
        src108 <= 12'hcf2;
        src109 <= 12'h2bf;
        src110 <= 12'h80c;
        src111 <= 12'hf7d;
        src112 <= 12'h7a2;
        src113 <= 12'hc6a;
        src114 <= 12'h965;
        src115 <= 12'h366;
        src116 <= 12'h35c;
        src117 <= 12'habb;
        src118 <= 12'h730;
        src119 <= 12'h5b6;
        src120 <= 12'h536;
        src121 <= 12'hb19;
        src122 <= 12'h436;
        src123 <= 12'h923;
        src124 <= 12'ha00;
        src125 <= 12'h4ff;
        src126 <= 12'he24;
        src127 <= 12'hd83;
        exp <= 19'h3e84c;
        #1
        src0 <= 12'hb56;
        src1 <= 12'h18c;
        src2 <= 12'hde5;
        src3 <= 12'hded;
        src4 <= 12'h3e4;
        src5 <= 12'h5a9;
        src6 <= 12'h4a7;
        src7 <= 12'hddd;
        src8 <= 12'hf4;
        src9 <= 12'hfe6;
        src10 <= 12'he73;
        src11 <= 12'h4e3;
        src12 <= 12'h2f8;
        src13 <= 12'hd35;
        src14 <= 12'h77;
        src15 <= 12'hd4c;
        src16 <= 12'he0e;
        src17 <= 12'hd11;
        src18 <= 12'hf2e;
        src19 <= 12'h781;
        src20 <= 12'hc35;
        src21 <= 12'hbf0;
        src22 <= 12'h460;
        src23 <= 12'hb83;
        src24 <= 12'h3f8;
        src25 <= 12'h89;
        src26 <= 12'ha17;
        src27 <= 12'hed6;
        src28 <= 12'h7a9;
        src29 <= 12'h917;
        src30 <= 12'h802;
        src31 <= 12'he21;
        src32 <= 12'h268;
        src33 <= 12'heab;
        src34 <= 12'h719;
        src35 <= 12'h893;
        src36 <= 12'h720;
        src37 <= 12'ha1d;
        src38 <= 12'h909;
        src39 <= 12'h5fc;
        src40 <= 12'hc7;
        src41 <= 12'haf0;
        src42 <= 12'h71f;
        src43 <= 12'h2a9;
        src44 <= 12'h336;
        src45 <= 12'h2d3;
        src46 <= 12'h981;
        src47 <= 12'hc6b;
        src48 <= 12'h29a;
        src49 <= 12'hd96;
        src50 <= 12'hb76;
        src51 <= 12'hba0;
        src52 <= 12'h209;
        src53 <= 12'h2b7;
        src54 <= 12'h636;
        src55 <= 12'hbe6;
        src56 <= 12'hd79;
        src57 <= 12'h445;
        src58 <= 12'hfc0;
        src59 <= 12'h92e;
        src60 <= 12'h2cf;
        src61 <= 12'hd3e;
        src62 <= 12'h3a4;
        src63 <= 12'h910;
        src64 <= 12'h6c3;
        src65 <= 12'he15;
        src66 <= 12'h151;
        src67 <= 12'h2b5;
        src68 <= 12'he2e;
        src69 <= 12'hab6;
        src70 <= 12'hcec;
        src71 <= 12'h875;
        src72 <= 12'hebe;
        src73 <= 12'hed7;
        src74 <= 12'hb8a;
        src75 <= 12'hfb0;
        src76 <= 12'h4e8;
        src77 <= 12'h9f4;
        src78 <= 12'hde8;
        src79 <= 12'h2b2;
        src80 <= 12'h81a;
        src81 <= 12'h70a;
        src82 <= 12'h83a;
        src83 <= 12'hee2;
        src84 <= 12'h8b7;
        src85 <= 12'h7af;
        src86 <= 12'h159;
        src87 <= 12'h2dc;
        src88 <= 12'hb90;
        src89 <= 12'h53f;
        src90 <= 12'heb;
        src91 <= 12'h743;
        src92 <= 12'hf30;
        src93 <= 12'ha93;
        src94 <= 12'h52a;
        src95 <= 12'h601;
        src96 <= 12'hbdc;
        src97 <= 12'h7df;
        src98 <= 12'h1fb;
        src99 <= 12'h3f9;
        src100 <= 12'h2d9;
        src101 <= 12'h316;
        src102 <= 12'h47c;
        src103 <= 12'h7b2;
        src104 <= 12'ha9;
        src105 <= 12'hd1b;
        src106 <= 12'hf15;
        src107 <= 12'hf07;
        src108 <= 12'h446;
        src109 <= 12'h8b9;
        src110 <= 12'hb8d;
        src111 <= 12'h65;
        src112 <= 12'hdf0;
        src113 <= 12'h1d0;
        src114 <= 12'h5bb;
        src115 <= 12'h1a7;
        src116 <= 12'ha2;
        src117 <= 12'ha17;
        src118 <= 12'hcc9;
        src119 <= 12'h272;
        src120 <= 12'h200;
        src121 <= 12'h48;
        src122 <= 12'h445;
        src123 <= 12'h551;
        src124 <= 12'h3fb;
        src125 <= 12'hec2;
        src126 <= 12'hd36;
        src127 <= 12'h7ad;
        exp <= 19'h40a6f;
        #1
        src0 <= 12'hafc;
        src1 <= 12'haeb;
        src2 <= 12'h61;
        src3 <= 12'h6cd;
        src4 <= 12'h6cb;
        src5 <= 12'hd74;
        src6 <= 12'hc50;
        src7 <= 12'h812;
        src8 <= 12'h4f8;
        src9 <= 12'h73;
        src10 <= 12'hdbe;
        src11 <= 12'h68a;
        src12 <= 12'h1e;
        src13 <= 12'h4ad;
        src14 <= 12'h740;
        src15 <= 12'hbf6;
        src16 <= 12'h82e;
        src17 <= 12'h9ae;
        src18 <= 12'h401;
        src19 <= 12'h6bc;
        src20 <= 12'he63;
        src21 <= 12'h1bb;
        src22 <= 12'hb46;
        src23 <= 12'hae;
        src24 <= 12'hfa0;
        src25 <= 12'h5c4;
        src26 <= 12'hbf7;
        src27 <= 12'hec0;
        src28 <= 12'hac8;
        src29 <= 12'h97f;
        src30 <= 12'h89e;
        src31 <= 12'h8a7;
        src32 <= 12'hc1d;
        src33 <= 12'h150;
        src34 <= 12'he64;
        src35 <= 12'ha6b;
        src36 <= 12'h5ba;
        src37 <= 12'hc8a;
        src38 <= 12'h6;
        src39 <= 12'h204;
        src40 <= 12'h678;
        src41 <= 12'h108;
        src42 <= 12'ha58;
        src43 <= 12'h18c;
        src44 <= 12'h6;
        src45 <= 12'hae1;
        src46 <= 12'h6ef;
        src47 <= 12'h95f;
        src48 <= 12'hc05;
        src49 <= 12'h49;
        src50 <= 12'h109;
        src51 <= 12'h11;
        src52 <= 12'hdd9;
        src53 <= 12'h349;
        src54 <= 12'hcc3;
        src55 <= 12'h43;
        src56 <= 12'h58c;
        src57 <= 12'hab1;
        src58 <= 12'h10d;
        src59 <= 12'h98c;
        src60 <= 12'h2e0;
        src61 <= 12'h53b;
        src62 <= 12'h9a9;
        src63 <= 12'h742;
        src64 <= 12'hcbd;
        src65 <= 12'h118;
        src66 <= 12'hfec;
        src67 <= 12'h248;
        src68 <= 12'h7e1;
        src69 <= 12'hdb1;
        src70 <= 12'h3e9;
        src71 <= 12'h680;
        src72 <= 12'h2e4;
        src73 <= 12'h3b6;
        src74 <= 12'he85;
        src75 <= 12'h62c;
        src76 <= 12'h114;
        src77 <= 12'hc72;
        src78 <= 12'h2ef;
        src79 <= 12'h219;
        src80 <= 12'h348;
        src81 <= 12'h391;
        src82 <= 12'h84c;
        src83 <= 12'h927;
        src84 <= 12'hebe;
        src85 <= 12'hb83;
        src86 <= 12'h4fb;
        src87 <= 12'hbb8;
        src88 <= 12'h67c;
        src89 <= 12'hf8a;
        src90 <= 12'h524;
        src91 <= 12'hf31;
        src92 <= 12'h921;
        src93 <= 12'h97b;
        src94 <= 12'hbb0;
        src95 <= 12'h605;
        src96 <= 12'hedf;
        src97 <= 12'h7b7;
        src98 <= 12'he95;
        src99 <= 12'hfe9;
        src100 <= 12'h878;
        src101 <= 12'h8a3;
        src102 <= 12'h519;
        src103 <= 12'h99d;
        src104 <= 12'h427;
        src105 <= 12'h9fd;
        src106 <= 12'h47b;
        src107 <= 12'hc1e;
        src108 <= 12'h50e;
        src109 <= 12'h5fb;
        src110 <= 12'h946;
        src111 <= 12'h1bd;
        src112 <= 12'h95e;
        src113 <= 12'h327;
        src114 <= 12'h493;
        src115 <= 12'h4d9;
        src116 <= 12'hec2;
        src117 <= 12'hc3c;
        src118 <= 12'h87f;
        src119 <= 12'hc7d;
        src120 <= 12'hbd0;
        src121 <= 12'h53c;
        src122 <= 12'h3a9;
        src123 <= 12'hc33;
        src124 <= 12'h8a8;
        src125 <= 12'hafe;
        src126 <= 12'hac;
        src127 <= 12'haa2;
        exp <= 19'h3dd89;
        #1
        src0 <= 12'h2b1;
        src1 <= 12'he5;
        src2 <= 12'h976;
        src3 <= 12'hb56;
        src4 <= 12'hb2f;
        src5 <= 12'h9cd;
        src6 <= 12'hbfd;
        src7 <= 12'h454;
        src8 <= 12'had;
        src9 <= 12'h4d7;
        src10 <= 12'h6;
        src11 <= 12'h443;
        src12 <= 12'h5d3;
        src13 <= 12'h2c2;
        src14 <= 12'hf18;
        src15 <= 12'ha64;
        src16 <= 12'h431;
        src17 <= 12'hcf2;
        src18 <= 12'h55f;
        src19 <= 12'hc89;
        src20 <= 12'h481;
        src21 <= 12'h984;
        src22 <= 12'hfcd;
        src23 <= 12'hcac;
        src24 <= 12'h11d;
        src25 <= 12'h31f;
        src26 <= 12'h8b8;
        src27 <= 12'hdd2;
        src28 <= 12'hadc;
        src29 <= 12'h17;
        src30 <= 12'h17;
        src31 <= 12'hed4;
        src32 <= 12'h6fa;
        src33 <= 12'hec5;
        src34 <= 12'h8;
        src35 <= 12'hcd1;
        src36 <= 12'hf9c;
        src37 <= 12'h549;
        src38 <= 12'ha78;
        src39 <= 12'h261;
        src40 <= 12'hdc7;
        src41 <= 12'h620;
        src42 <= 12'h584;
        src43 <= 12'hca1;
        src44 <= 12'hb7c;
        src45 <= 12'h4db;
        src46 <= 12'h339;
        src47 <= 12'h9c;
        src48 <= 12'h41;
        src49 <= 12'h652;
        src50 <= 12'h149;
        src51 <= 12'he47;
        src52 <= 12'hcd4;
        src53 <= 12'h146;
        src54 <= 12'h8c6;
        src55 <= 12'ha80;
        src56 <= 12'h679;
        src57 <= 12'hcee;
        src58 <= 12'hbe;
        src59 <= 12'h30c;
        src60 <= 12'h358;
        src61 <= 12'h24e;
        src62 <= 12'h213;
        src63 <= 12'h182;
        src64 <= 12'h31c;
        src65 <= 12'h473;
        src66 <= 12'h2bc;
        src67 <= 12'hcb8;
        src68 <= 12'h79e;
        src69 <= 12'h8f2;
        src70 <= 12'h76d;
        src71 <= 12'h6d5;
        src72 <= 12'hc4;
        src73 <= 12'hafc;
        src74 <= 12'ha72;
        src75 <= 12'h7bd;
        src76 <= 12'h18b;
        src77 <= 12'h48b;
        src78 <= 12'hc81;
        src79 <= 12'h6c4;
        src80 <= 12'hf2a;
        src81 <= 12'h759;
        src82 <= 12'h1e4;
        src83 <= 12'h85;
        src84 <= 12'heba;
        src85 <= 12'h8ce;
        src86 <= 12'h81;
        src87 <= 12'he12;
        src88 <= 12'hb00;
        src89 <= 12'h97a;
        src90 <= 12'hfb;
        src91 <= 12'hfb9;
        src92 <= 12'h172;
        src93 <= 12'hf4;
        src94 <= 12'h929;
        src95 <= 12'hfbf;
        src96 <= 12'h505;
        src97 <= 12'hc69;
        src98 <= 12'hd80;
        src99 <= 12'hbab;
        src100 <= 12'h5c5;
        src101 <= 12'hb74;
        src102 <= 12'hb86;
        src103 <= 12'hbae;
        src104 <= 12'h19d;
        src105 <= 12'h45b;
        src106 <= 12'h7d0;
        src107 <= 12'h514;
        src108 <= 12'hebb;
        src109 <= 12'hbdf;
        src110 <= 12'h97d;
        src111 <= 12'h72d;
        src112 <= 12'he3e;
        src113 <= 12'h577;
        src114 <= 12'hfc0;
        src115 <= 12'h6a6;
        src116 <= 12'h80c;
        src117 <= 12'hdb7;
        src118 <= 12'hcad;
        src119 <= 12'h464;
        src120 <= 12'he59;
        src121 <= 12'hf14;
        src122 <= 12'hf1d;
        src123 <= 12'h711;
        src124 <= 12'h830;
        src125 <= 12'h6ee;
        src126 <= 12'hae9;
        src127 <= 12'h7d6;
        exp <= 19'h3e666;
        #1
        src0 <= 12'h41f;
        src1 <= 12'hff8;
        src2 <= 12'hb5e;
        src3 <= 12'h63e;
        src4 <= 12'ha79;
        src5 <= 12'h5e;
        src6 <= 12'h154;
        src7 <= 12'h4ba;
        src8 <= 12'h4b3;
        src9 <= 12'hd30;
        src10 <= 12'he8b;
        src11 <= 12'h2f4;
        src12 <= 12'h267;
        src13 <= 12'h828;
        src14 <= 12'h3a;
        src15 <= 12'h6a7;
        src16 <= 12'h178;
        src17 <= 12'he24;
        src18 <= 12'h12f;
        src19 <= 12'h86c;
        src20 <= 12'h79b;
        src21 <= 12'hd10;
        src22 <= 12'h542;
        src23 <= 12'h579;
        src24 <= 12'hae3;
        src25 <= 12'h945;
        src26 <= 12'h11e;
        src27 <= 12'h965;
        src28 <= 12'hd07;
        src29 <= 12'ha5a;
        src30 <= 12'hdd4;
        src31 <= 12'hb31;
        src32 <= 12'hbcd;
        src33 <= 12'hea3;
        src34 <= 12'h17d;
        src35 <= 12'hea0;
        src36 <= 12'hc0b;
        src37 <= 12'h95a;
        src38 <= 12'hd2e;
        src39 <= 12'hb11;
        src40 <= 12'h200;
        src41 <= 12'h6c6;
        src42 <= 12'hada;
        src43 <= 12'h6d5;
        src44 <= 12'h1fc;
        src45 <= 12'h520;
        src46 <= 12'h603;
        src47 <= 12'hc61;
        src48 <= 12'h5b8;
        src49 <= 12'hea0;
        src50 <= 12'hf8b;
        src51 <= 12'hdda;
        src52 <= 12'h918;
        src53 <= 12'h6d;
        src54 <= 12'h668;
        src55 <= 12'hfff;
        src56 <= 12'h14d;
        src57 <= 12'h7e5;
        src58 <= 12'heda;
        src59 <= 12'h5f7;
        src60 <= 12'hbc5;
        src61 <= 12'h9c6;
        src62 <= 12'h2a7;
        src63 <= 12'h1ee;
        src64 <= 12'hc02;
        src65 <= 12'h717;
        src66 <= 12'h7ae;
        src67 <= 12'hc22;
        src68 <= 12'h1d5;
        src69 <= 12'h653;
        src70 <= 12'h4bf;
        src71 <= 12'h10b;
        src72 <= 12'he8;
        src73 <= 12'hbe8;
        src74 <= 12'h576;
        src75 <= 12'h411;
        src76 <= 12'h2fa;
        src77 <= 12'hbb7;
        src78 <= 12'h382;
        src79 <= 12'h867;
        src80 <= 12'haf4;
        src81 <= 12'hdb8;
        src82 <= 12'h18;
        src83 <= 12'h4f;
        src84 <= 12'h507;
        src85 <= 12'h6ed;
        src86 <= 12'h5ab;
        src87 <= 12'h935;
        src88 <= 12'h60c;
        src89 <= 12'h9f6;
        src90 <= 12'hd2f;
        src91 <= 12'hd92;
        src92 <= 12'hb6b;
        src93 <= 12'h653;
        src94 <= 12'hd59;
        src95 <= 12'h13d;
        src96 <= 12'hab8;
        src97 <= 12'h335;
        src98 <= 12'hedd;
        src99 <= 12'hb50;
        src100 <= 12'h14b;
        src101 <= 12'hc86;
        src102 <= 12'h375;
        src103 <= 12'h3c5;
        src104 <= 12'h414;
        src105 <= 12'hf08;
        src106 <= 12'h836;
        src107 <= 12'he06;
        src108 <= 12'ha4;
        src109 <= 12'hcfa;
        src110 <= 12'h805;
        src111 <= 12'h1ce;
        src112 <= 12'h649;
        src113 <= 12'ha7b;
        src114 <= 12'h1f7;
        src115 <= 12'h33a;
        src116 <= 12'h9d5;
        src117 <= 12'h1e5;
        src118 <= 12'h441;
        src119 <= 12'hdb3;
        src120 <= 12'h451;
        src121 <= 12'hafd;
        src122 <= 12'h4c;
        src123 <= 12'hf4d;
        src124 <= 12'hf7;
        src125 <= 12'hd46;
        src126 <= 12'he09;
        src127 <= 12'hc5e;
        exp <= 19'h3e6f0;
        #1
        src0 <= 12'hf1e;
        src1 <= 12'ha1a;
        src2 <= 12'hd67;
        src3 <= 12'h752;
        src4 <= 12'haca;
        src5 <= 12'h822;
        src6 <= 12'h149;
        src7 <= 12'hef0;
        src8 <= 12'ha35;
        src9 <= 12'ha32;
        src10 <= 12'h319;
        src11 <= 12'h15b;
        src12 <= 12'h7d8;
        src13 <= 12'ha20;
        src14 <= 12'h6b5;
        src15 <= 12'hc8d;
        src16 <= 12'hd1d;
        src17 <= 12'h72;
        src18 <= 12'h601;
        src19 <= 12'h520;
        src20 <= 12'heda;
        src21 <= 12'hb27;
        src22 <= 12'h1b;
        src23 <= 12'h95d;
        src24 <= 12'he41;
        src25 <= 12'h302;
        src26 <= 12'hd8d;
        src27 <= 12'hea5;
        src28 <= 12'h189;
        src29 <= 12'h1d4;
        src30 <= 12'h79;
        src31 <= 12'h765;
        src32 <= 12'haff;
        src33 <= 12'hfc3;
        src34 <= 12'h85f;
        src35 <= 12'h43c;
        src36 <= 12'h1d9;
        src37 <= 12'h6f2;
        src38 <= 12'hfdd;
        src39 <= 12'hb27;
        src40 <= 12'hdd0;
        src41 <= 12'ha24;
        src42 <= 12'h1bf;
        src43 <= 12'h247;
        src44 <= 12'he4a;
        src45 <= 12'he9;
        src46 <= 12'he40;
        src47 <= 12'h620;
        src48 <= 12'h8e2;
        src49 <= 12'h49c;
        src50 <= 12'h15d;
        src51 <= 12'h9fc;
        src52 <= 12'h596;
        src53 <= 12'he20;
        src54 <= 12'habf;
        src55 <= 12'h9cc;
        src56 <= 12'h23c;
        src57 <= 12'h94c;
        src58 <= 12'hc2f;
        src59 <= 12'hd04;
        src60 <= 12'h1b9;
        src61 <= 12'hed4;
        src62 <= 12'he2d;
        src63 <= 12'he52;
        src64 <= 12'hdba;
        src65 <= 12'hea7;
        src66 <= 12'hd8;
        src67 <= 12'hcae;
        src68 <= 12'h671;
        src69 <= 12'hf7;
        src70 <= 12'hcda;
        src71 <= 12'h68d;
        src72 <= 12'h267;
        src73 <= 12'h6ca;
        src74 <= 12'h3d0;
        src75 <= 12'hfb0;
        src76 <= 12'hf77;
        src77 <= 12'h2e1;
        src78 <= 12'h455;
        src79 <= 12'h600;
        src80 <= 12'h704;
        src81 <= 12'hab;
        src82 <= 12'ha3b;
        src83 <= 12'h242;
        src84 <= 12'hac5;
        src85 <= 12'h5c0;
        src86 <= 12'h719;
        src87 <= 12'h805;
        src88 <= 12'hf3c;
        src89 <= 12'h67e;
        src90 <= 12'hacd;
        src91 <= 12'hb6;
        src92 <= 12'hf8a;
        src93 <= 12'h792;
        src94 <= 12'hb1;
        src95 <= 12'h272;
        src96 <= 12'hed6;
        src97 <= 12'h5dc;
        src98 <= 12'h94f;
        src99 <= 12'hefc;
        src100 <= 12'h644;
        src101 <= 12'hc3a;
        src102 <= 12'h3bd;
        src103 <= 12'h34;
        src104 <= 12'h717;
        src105 <= 12'h6c5;
        src106 <= 12'h9c6;
        src107 <= 12'h2bb;
        src108 <= 12'hbcd;
        src109 <= 12'hdda;
        src110 <= 12'h31c;
        src111 <= 12'hc6c;
        src112 <= 12'h7ef;
        src113 <= 12'h125;
        src114 <= 12'hc43;
        src115 <= 12'ha37;
        src116 <= 12'h548;
        src117 <= 12'ha78;
        src118 <= 12'h116;
        src119 <= 12'he7a;
        src120 <= 12'h814;
        src121 <= 12'h398;
        src122 <= 12'h1e1;
        src123 <= 12'h512;
        src124 <= 12'h3e8;
        src125 <= 12'h472;
        src126 <= 12'hda;
        src127 <= 12'he1b;
        exp <= 19'h3febf;
        #1
        src0 <= 12'h8e4;
        src1 <= 12'h9d;
        src2 <= 12'h4b3;
        src3 <= 12'hd4c;
        src4 <= 12'h1c0;
        src5 <= 12'h693;
        src6 <= 12'h2fd;
        src7 <= 12'hbd5;
        src8 <= 12'h856;
        src9 <= 12'hbfb;
        src10 <= 12'hef6;
        src11 <= 12'h88f;
        src12 <= 12'h483;
        src13 <= 12'h364;
        src14 <= 12'h43a;
        src15 <= 12'h71b;
        src16 <= 12'h1f;
        src17 <= 12'h22b;
        src18 <= 12'h126;
        src19 <= 12'h7e4;
        src20 <= 12'hab8;
        src21 <= 12'h5cd;
        src22 <= 12'h219;
        src23 <= 12'h8ee;
        src24 <= 12'hc23;
        src25 <= 12'h490;
        src26 <= 12'h1d9;
        src27 <= 12'h6e6;
        src28 <= 12'h853;
        src29 <= 12'hcaa;
        src30 <= 12'h5b4;
        src31 <= 12'hcd2;
        src32 <= 12'h670;
        src33 <= 12'h6dd;
        src34 <= 12'h697;
        src35 <= 12'h29f;
        src36 <= 12'hed1;
        src37 <= 12'h44d;
        src38 <= 12'hd8a;
        src39 <= 12'hd2b;
        src40 <= 12'h8f9;
        src41 <= 12'hce2;
        src42 <= 12'h192;
        src43 <= 12'hf7f;
        src44 <= 12'h1e5;
        src45 <= 12'hc54;
        src46 <= 12'hf53;
        src47 <= 12'ha5c;
        src48 <= 12'h1bc;
        src49 <= 12'hb7d;
        src50 <= 12'haec;
        src51 <= 12'hbb8;
        src52 <= 12'h536;
        src53 <= 12'h885;
        src54 <= 12'h52d;
        src55 <= 12'hfcb;
        src56 <= 12'hbcb;
        src57 <= 12'ha6e;
        src58 <= 12'h659;
        src59 <= 12'hc17;
        src60 <= 12'hdae;
        src61 <= 12'hd53;
        src62 <= 12'h40a;
        src63 <= 12'hc45;
        src64 <= 12'h85f;
        src65 <= 12'ha1;
        src66 <= 12'h634;
        src67 <= 12'hecc;
        src68 <= 12'hbb0;
        src69 <= 12'h4fb;
        src70 <= 12'hcf6;
        src71 <= 12'hf2a;
        src72 <= 12'he96;
        src73 <= 12'he7;
        src74 <= 12'h83a;
        src75 <= 12'hb15;
        src76 <= 12'h1fd;
        src77 <= 12'h312;
        src78 <= 12'h134;
        src79 <= 12'hf0d;
        src80 <= 12'h1ae;
        src81 <= 12'hfe;
        src82 <= 12'h649;
        src83 <= 12'h70e;
        src84 <= 12'h9a9;
        src85 <= 12'h4fd;
        src86 <= 12'h1d0;
        src87 <= 12'ha2d;
        src88 <= 12'ha1e;
        src89 <= 12'h6fa;
        src90 <= 12'hed0;
        src91 <= 12'heb3;
        src92 <= 12'h3e1;
        src93 <= 12'h22c;
        src94 <= 12'he7;
        src95 <= 12'hf65;
        src96 <= 12'hff4;
        src97 <= 12'hac9;
        src98 <= 12'h8ee;
        src99 <= 12'h729;
        src100 <= 12'h21d;
        src101 <= 12'h4ca;
        src102 <= 12'he7e;
        src103 <= 12'hd86;
        src104 <= 12'h656;
        src105 <= 12'ha24;
        src106 <= 12'h7c5;
        src107 <= 12'h347;
        src108 <= 12'ha5b;
        src109 <= 12'hf53;
        src110 <= 12'h86;
        src111 <= 12'h881;
        src112 <= 12'h27b;
        src113 <= 12'h5cd;
        src114 <= 12'h66e;
        src115 <= 12'h5ff;
        src116 <= 12'h22b;
        src117 <= 12'he3c;
        src118 <= 12'h698;
        src119 <= 12'he2f;
        src120 <= 12'h859;
        src121 <= 12'hf32;
        src122 <= 12'hc2;
        src123 <= 12'h4c7;
        src124 <= 12'h687;
        src125 <= 12'h20;
        src126 <= 12'hed2;
        src127 <= 12'h685;
        exp <= 19'h3f8af;
        #1
        src0 <= 12'had0;
        src1 <= 12'h342;
        src2 <= 12'hb57;
        src3 <= 12'h45e;
        src4 <= 12'h85c;
        src5 <= 12'hda6;
        src6 <= 12'h5d;
        src7 <= 12'h36c;
        src8 <= 12'h4f;
        src9 <= 12'h9ec;
        src10 <= 12'hf37;
        src11 <= 12'h4f5;
        src12 <= 12'hd0a;
        src13 <= 12'hdc1;
        src14 <= 12'h703;
        src15 <= 12'h7eb;
        src16 <= 12'h12b;
        src17 <= 12'h52d;
        src18 <= 12'hae7;
        src19 <= 12'hf6;
        src20 <= 12'he6d;
        src21 <= 12'h389;
        src22 <= 12'h533;
        src23 <= 12'h12c;
        src24 <= 12'h50e;
        src25 <= 12'h84c;
        src26 <= 12'h1cc;
        src27 <= 12'ha98;
        src28 <= 12'hbf7;
        src29 <= 12'hfeb;
        src30 <= 12'h1f2;
        src31 <= 12'h6dc;
        src32 <= 12'h1b8;
        src33 <= 12'hf40;
        src34 <= 12'h8fb;
        src35 <= 12'hb73;
        src36 <= 12'h5c4;
        src37 <= 12'h116;
        src38 <= 12'h392;
        src39 <= 12'h41;
        src40 <= 12'hd0;
        src41 <= 12'h9f2;
        src42 <= 12'hf93;
        src43 <= 12'h4a;
        src44 <= 12'h8f5;
        src45 <= 12'h140;
        src46 <= 12'h6c2;
        src47 <= 12'hca4;
        src48 <= 12'h783;
        src49 <= 12'ha78;
        src50 <= 12'h2f6;
        src51 <= 12'h4ab;
        src52 <= 12'h7da;
        src53 <= 12'hb04;
        src54 <= 12'he6e;
        src55 <= 12'hefe;
        src56 <= 12'h26b;
        src57 <= 12'hb8c;
        src58 <= 12'hdd1;
        src59 <= 12'hcca;
        src60 <= 12'h48c;
        src61 <= 12'h38b;
        src62 <= 12'hfab;
        src63 <= 12'hcc7;
        src64 <= 12'hb04;
        src65 <= 12'h32b;
        src66 <= 12'hf8;
        src67 <= 12'h509;
        src68 <= 12'hc09;
        src69 <= 12'he18;
        src70 <= 12'h122;
        src71 <= 12'hfd0;
        src72 <= 12'h83e;
        src73 <= 12'h326;
        src74 <= 12'h4ce;
        src75 <= 12'hc8e;
        src76 <= 12'hcaf;
        src77 <= 12'h158;
        src78 <= 12'h38;
        src79 <= 12'h79d;
        src80 <= 12'hb78;
        src81 <= 12'h5c5;
        src82 <= 12'hec3;
        src83 <= 12'hfb9;
        src84 <= 12'he40;
        src85 <= 12'hca6;
        src86 <= 12'hf43;
        src87 <= 12'h79b;
        src88 <= 12'hc68;
        src89 <= 12'h2e9;
        src90 <= 12'h4f2;
        src91 <= 12'h774;
        src92 <= 12'h4dd;
        src93 <= 12'hbe;
        src94 <= 12'h919;
        src95 <= 12'h721;
        src96 <= 12'h3cc;
        src97 <= 12'hc05;
        src98 <= 12'h906;
        src99 <= 12'h667;
        src100 <= 12'h3bd;
        src101 <= 12'h187;
        src102 <= 12'h2f8;
        src103 <= 12'h6e4;
        src104 <= 12'hd26;
        src105 <= 12'h7d2;
        src106 <= 12'hddb;
        src107 <= 12'h6e;
        src108 <= 12'hed0;
        src109 <= 12'hcaa;
        src110 <= 12'h413;
        src111 <= 12'hdd;
        src112 <= 12'hba2;
        src113 <= 12'hd4c;
        src114 <= 12'hfd0;
        src115 <= 12'hc90;
        src116 <= 12'heb6;
        src117 <= 12'hf7;
        src118 <= 12'h690;
        src119 <= 12'hb34;
        src120 <= 12'h6bb;
        src121 <= 12'hcb;
        src122 <= 12'hb2b;
        src123 <= 12'hcfb;
        src124 <= 12'h65f;
        src125 <= 12'hbae;
        src126 <= 12'hf90;
        src127 <= 12'hd08;
        exp <= 19'h403f9;
        #1
        src0 <= 12'h4a6;
        src1 <= 12'hd19;
        src2 <= 12'hc9a;
        src3 <= 12'h775;
        src4 <= 12'h5d9;
        src5 <= 12'h399;
        src6 <= 12'hed4;
        src7 <= 12'h3f;
        src8 <= 12'h140;
        src9 <= 12'h77b;
        src10 <= 12'h7cb;
        src11 <= 12'h715;
        src12 <= 12'hdc3;
        src13 <= 12'hace;
        src14 <= 12'h229;
        src15 <= 12'h795;
        src16 <= 12'he62;
        src17 <= 12'h4a5;
        src18 <= 12'h211;
        src19 <= 12'h426;
        src20 <= 12'h53d;
        src21 <= 12'h939;
        src22 <= 12'h1a8;
        src23 <= 12'hb95;
        src24 <= 12'h3be;
        src25 <= 12'h1ca;
        src26 <= 12'hda7;
        src27 <= 12'hd10;
        src28 <= 12'h930;
        src29 <= 12'haba;
        src30 <= 12'h4c3;
        src31 <= 12'h637;
        src32 <= 12'h6fe;
        src33 <= 12'h34a;
        src34 <= 12'ha04;
        src35 <= 12'h6a9;
        src36 <= 12'hb10;
        src37 <= 12'hc14;
        src38 <= 12'h693;
        src39 <= 12'h337;
        src40 <= 12'h5ae;
        src41 <= 12'hd3a;
        src42 <= 12'he6a;
        src43 <= 12'h759;
        src44 <= 12'h77c;
        src45 <= 12'he44;
        src46 <= 12'h331;
        src47 <= 12'h5d5;
        src48 <= 12'h218;
        src49 <= 12'hffe;
        src50 <= 12'h236;
        src51 <= 12'h86a;
        src52 <= 12'hd9;
        src53 <= 12'hff9;
        src54 <= 12'h968;
        src55 <= 12'h8ff;
        src56 <= 12'hcda;
        src57 <= 12'heb7;
        src58 <= 12'hbdd;
        src59 <= 12'h9cd;
        src60 <= 12'hf41;
        src61 <= 12'h43d;
        src62 <= 12'h719;
        src63 <= 12'h3cd;
        src64 <= 12'hc67;
        src65 <= 12'h469;
        src66 <= 12'h8c9;
        src67 <= 12'h8ee;
        src68 <= 12'hd3;
        src69 <= 12'h375;
        src70 <= 12'h4d1;
        src71 <= 12'hf55;
        src72 <= 12'h5ce;
        src73 <= 12'hfdb;
        src74 <= 12'h1b3;
        src75 <= 12'h947;
        src76 <= 12'h508;
        src77 <= 12'h2b0;
        src78 <= 12'hae5;
        src79 <= 12'ha00;
        src80 <= 12'ha50;
        src81 <= 12'h26a;
        src82 <= 12'h76b;
        src83 <= 12'h384;
        src84 <= 12'h370;
        src85 <= 12'h5a2;
        src86 <= 12'he88;
        src87 <= 12'h7f1;
        src88 <= 12'h76c;
        src89 <= 12'h99d;
        src90 <= 12'hcdd;
        src91 <= 12'hf86;
        src92 <= 12'he24;
        src93 <= 12'h206;
        src94 <= 12'h474;
        src95 <= 12'hdbd;
        src96 <= 12'hf96;
        src97 <= 12'h464;
        src98 <= 12'h7e9;
        src99 <= 12'h24c;
        src100 <= 12'hd1e;
        src101 <= 12'h71d;
        src102 <= 12'hd4a;
        src103 <= 12'h3cf;
        src104 <= 12'h97f;
        src105 <= 12'hdbf;
        src106 <= 12'h9c4;
        src107 <= 12'h1e3;
        src108 <= 12'h830;
        src109 <= 12'h35c;
        src110 <= 12'heaf;
        src111 <= 12'hd08;
        src112 <= 12'h365;
        src113 <= 12'h6c6;
        src114 <= 12'hcc;
        src115 <= 12'hf46;
        src116 <= 12'h21c;
        src117 <= 12'ha55;
        src118 <= 12'h81c;
        src119 <= 12'hd4e;
        src120 <= 12'h90e;
        src121 <= 12'h81e;
        src122 <= 12'hadc;
        src123 <= 12'h57a;
        src124 <= 12'h46;
        src125 <= 12'h7c6;
        src126 <= 12'h2ee;
        src127 <= 12'h58f;
        exp <= 19'h3fa31;
        #1
        src0 <= 12'h99e;
        src1 <= 12'h1f9;
        src2 <= 12'h6b5;
        src3 <= 12'hf66;
        src4 <= 12'h95;
        src5 <= 12'h18;
        src6 <= 12'h5a3;
        src7 <= 12'hfd1;
        src8 <= 12'h68f;
        src9 <= 12'h3c;
        src10 <= 12'h478;
        src11 <= 12'h8af;
        src12 <= 12'hb39;
        src13 <= 12'hb08;
        src14 <= 12'h764;
        src15 <= 12'hade;
        src16 <= 12'h43a;
        src17 <= 12'hdef;
        src18 <= 12'hc2;
        src19 <= 12'hd4c;
        src20 <= 12'h237;
        src21 <= 12'h5fa;
        src22 <= 12'h329;
        src23 <= 12'h1a8;
        src24 <= 12'hf3a;
        src25 <= 12'h538;
        src26 <= 12'ha46;
        src27 <= 12'h3d0;
        src28 <= 12'h74a;
        src29 <= 12'haf3;
        src30 <= 12'h65d;
        src31 <= 12'h97e;
        src32 <= 12'hb0f;
        src33 <= 12'hea8;
        src34 <= 12'hbbd;
        src35 <= 12'h115;
        src36 <= 12'had7;
        src37 <= 12'h77d;
        src38 <= 12'hb9c;
        src39 <= 12'h808;
        src40 <= 12'h573;
        src41 <= 12'hdc8;
        src42 <= 12'h92e;
        src43 <= 12'h760;
        src44 <= 12'ha4a;
        src45 <= 12'hf54;
        src46 <= 12'h6e4;
        src47 <= 12'h830;
        src48 <= 12'he96;
        src49 <= 12'hbf5;
        src50 <= 12'h42e;
        src51 <= 12'h4d8;
        src52 <= 12'h76f;
        src53 <= 12'h3ad;
        src54 <= 12'h99f;
        src55 <= 12'h50b;
        src56 <= 12'h967;
        src57 <= 12'h638;
        src58 <= 12'h777;
        src59 <= 12'he7c;
        src60 <= 12'h393;
        src61 <= 12'h433;
        src62 <= 12'h187;
        src63 <= 12'h43a;
        src64 <= 12'h2c7;
        src65 <= 12'hf73;
        src66 <= 12'hf51;
        src67 <= 12'h1ac;
        src68 <= 12'h651;
        src69 <= 12'hcdd;
        src70 <= 12'hacd;
        src71 <= 12'h719;
        src72 <= 12'h3f3;
        src73 <= 12'h578;
        src74 <= 12'he22;
        src75 <= 12'h9f3;
        src76 <= 12'h31b;
        src77 <= 12'hb6c;
        src78 <= 12'h419;
        src79 <= 12'h8a4;
        src80 <= 12'h4fe;
        src81 <= 12'had0;
        src82 <= 12'hc4a;
        src83 <= 12'h23c;
        src84 <= 12'hb2a;
        src85 <= 12'h345;
        src86 <= 12'h207;
        src87 <= 12'h83a;
        src88 <= 12'hdf0;
        src89 <= 12'hc5f;
        src90 <= 12'h4ba;
        src91 <= 12'hc00;
        src92 <= 12'he82;
        src93 <= 12'hcc0;
        src94 <= 12'hd42;
        src95 <= 12'hb0b;
        src96 <= 12'h47b;
        src97 <= 12'h9e8;
        src98 <= 12'hc75;
        src99 <= 12'h102;
        src100 <= 12'he90;
        src101 <= 12'hb33;
        src102 <= 12'h150;
        src103 <= 12'h876;
        src104 <= 12'h33;
        src105 <= 12'h5c3;
        src106 <= 12'h171;
        src107 <= 12'hc8e;
        src108 <= 12'hdf6;
        src109 <= 12'hca2;
        src110 <= 12'hd41;
        src111 <= 12'hb0b;
        src112 <= 12'hdaa;
        src113 <= 12'h3f3;
        src114 <= 12'h75c;
        src115 <= 12'hb33;
        src116 <= 12'h30b;
        src117 <= 12'h6f5;
        src118 <= 12'h52e;
        src119 <= 12'hc53;
        src120 <= 12'h1f;
        src121 <= 12'h644;
        src122 <= 12'h7c7;
        src123 <= 12'hb0b;
        src124 <= 12'hdb9;
        src125 <= 12'heac;
        src126 <= 12'ha7d;
        src127 <= 12'h40f;
        exp <= 19'h41447;
        #1
        src0 <= 12'h587;
        src1 <= 12'h669;
        src2 <= 12'he00;
        src3 <= 12'h3e9;
        src4 <= 12'h4b1;
        src5 <= 12'h275;
        src6 <= 12'hec3;
        src7 <= 12'h27a;
        src8 <= 12'ha8f;
        src9 <= 12'h43d;
        src10 <= 12'h921;
        src11 <= 12'hd5f;
        src12 <= 12'hd60;
        src13 <= 12'he17;
        src14 <= 12'h61a;
        src15 <= 12'h748;
        src16 <= 12'h8cd;
        src17 <= 12'he1d;
        src18 <= 12'h812;
        src19 <= 12'hd92;
        src20 <= 12'h267;
        src21 <= 12'h3fc;
        src22 <= 12'hba9;
        src23 <= 12'h2b8;
        src24 <= 12'h72f;
        src25 <= 12'h1a1;
        src26 <= 12'he93;
        src27 <= 12'h85e;
        src28 <= 12'ha3f;
        src29 <= 12'h48a;
        src30 <= 12'h5e8;
        src31 <= 12'h45e;
        src32 <= 12'he09;
        src33 <= 12'hf3c;
        src34 <= 12'h26f;
        src35 <= 12'he62;
        src36 <= 12'hbba;
        src37 <= 12'h23d;
        src38 <= 12'h6bf;
        src39 <= 12'h92;
        src40 <= 12'h8bf;
        src41 <= 12'hc3d;
        src42 <= 12'hf24;
        src43 <= 12'h6c2;
        src44 <= 12'h9bc;
        src45 <= 12'h749;
        src46 <= 12'h1a6;
        src47 <= 12'h84c;
        src48 <= 12'h1da;
        src49 <= 12'hf18;
        src50 <= 12'hb07;
        src51 <= 12'h852;
        src52 <= 12'h547;
        src53 <= 12'h1a9;
        src54 <= 12'h256;
        src55 <= 12'h2d;
        src56 <= 12'h1f5;
        src57 <= 12'h89b;
        src58 <= 12'h758;
        src59 <= 12'hf36;
        src60 <= 12'h5ab;
        src61 <= 12'haee;
        src62 <= 12'h60f;
        src63 <= 12'h2f2;
        src64 <= 12'h3bf;
        src65 <= 12'h760;
        src66 <= 12'h9e3;
        src67 <= 12'h17c;
        src68 <= 12'ha1b;
        src69 <= 12'h75c;
        src70 <= 12'haa3;
        src71 <= 12'hd20;
        src72 <= 12'hf48;
        src73 <= 12'h83f;
        src74 <= 12'haf5;
        src75 <= 12'h3a3;
        src76 <= 12'h40f;
        src77 <= 12'h2e6;
        src78 <= 12'hc08;
        src79 <= 12'h81f;
        src80 <= 12'h743;
        src81 <= 12'h8f8;
        src82 <= 12'h173;
        src83 <= 12'haf5;
        src84 <= 12'h68a;
        src85 <= 12'h667;
        src86 <= 12'h9c7;
        src87 <= 12'h929;
        src88 <= 12'hbf7;
        src89 <= 12'hfc7;
        src90 <= 12'hb9a;
        src91 <= 12'h64b;
        src92 <= 12'h9f3;
        src93 <= 12'hd64;
        src94 <= 12'h9e3;
        src95 <= 12'hc28;
        src96 <= 12'h66b;
        src97 <= 12'he37;
        src98 <= 12'hc3e;
        src99 <= 12'h100;
        src100 <= 12'h549;
        src101 <= 12'h5c;
        src102 <= 12'hed9;
        src103 <= 12'hae0;
        src104 <= 12'hc97;
        src105 <= 12'hf1;
        src106 <= 12'ha44;
        src107 <= 12'h8db;
        src108 <= 12'h935;
        src109 <= 12'h867;
        src110 <= 12'h501;
        src111 <= 12'h481;
        src112 <= 12'hbce;
        src113 <= 12'h132;
        src114 <= 12'h8f2;
        src115 <= 12'hdca;
        src116 <= 12'h3aa;
        src117 <= 12'h32c;
        src118 <= 12'hef8;
        src119 <= 12'hcbd;
        src120 <= 12'hd65;
        src121 <= 12'h1a6;
        src122 <= 12'h714;
        src123 <= 12'h8ad;
        src124 <= 12'h712;
        src125 <= 12'hfe8;
        src126 <= 12'hc2f;
        src127 <= 12'h2a9;
        exp <= 19'h41094;
        #1
        src0 <= 12'hfb3;
        src1 <= 12'h1ea;
        src2 <= 12'h5c9;
        src3 <= 12'h154;
        src4 <= 12'he9e;
        src5 <= 12'h9ae;
        src6 <= 12'hc6c;
        src7 <= 12'h4f7;
        src8 <= 12'h564;
        src9 <= 12'h9e1;
        src10 <= 12'hac7;
        src11 <= 12'h4b8;
        src12 <= 12'h12e;
        src13 <= 12'he78;
        src14 <= 12'ha3d;
        src15 <= 12'h384;
        src16 <= 12'hc6;
        src17 <= 12'h181;
        src18 <= 12'h7dd;
        src19 <= 12'hda6;
        src20 <= 12'h733;
        src21 <= 12'hcd2;
        src22 <= 12'hd69;
        src23 <= 12'h667;
        src24 <= 12'h866;
        src25 <= 12'h9c3;
        src26 <= 12'hb48;
        src27 <= 12'hef6;
        src28 <= 12'h699;
        src29 <= 12'h5ec;
        src30 <= 12'hc7c;
        src31 <= 12'hfc;
        src32 <= 12'hb27;
        src33 <= 12'hb8e;
        src34 <= 12'hb4e;
        src35 <= 12'hb7;
        src36 <= 12'hbca;
        src37 <= 12'h936;
        src38 <= 12'h4c8;
        src39 <= 12'h194;
        src40 <= 12'h7a4;
        src41 <= 12'h1f6;
        src42 <= 12'h82b;
        src43 <= 12'h943;
        src44 <= 12'hc54;
        src45 <= 12'h649;
        src46 <= 12'h98b;
        src47 <= 12'h89a;
        src48 <= 12'hc88;
        src49 <= 12'h819;
        src50 <= 12'h44a;
        src51 <= 12'hfec;
        src52 <= 12'h6f2;
        src53 <= 12'hbe6;
        src54 <= 12'h28d;
        src55 <= 12'h330;
        src56 <= 12'hbfd;
        src57 <= 12'h140;
        src58 <= 12'h9c5;
        src59 <= 12'hb73;
        src60 <= 12'h17;
        src61 <= 12'he81;
        src62 <= 12'h2c7;
        src63 <= 12'hc43;
        src64 <= 12'hc13;
        src65 <= 12'h6f5;
        src66 <= 12'h286;
        src67 <= 12'hbe6;
        src68 <= 12'h682;
        src69 <= 12'h9;
        src70 <= 12'hd72;
        src71 <= 12'h8dd;
        src72 <= 12'hb20;
        src73 <= 12'h8d8;
        src74 <= 12'hfaa;
        src75 <= 12'h311;
        src76 <= 12'h303;
        src77 <= 12'h776;
        src78 <= 12'hac0;
        src79 <= 12'h557;
        src80 <= 12'h5e1;
        src81 <= 12'hfda;
        src82 <= 12'h7e3;
        src83 <= 12'ha28;
        src84 <= 12'h280;
        src85 <= 12'h229;
        src86 <= 12'h5c;
        src87 <= 12'h73e;
        src88 <= 12'h497;
        src89 <= 12'h9ab;
        src90 <= 12'h365;
        src91 <= 12'h869;
        src92 <= 12'haff;
        src93 <= 12'h778;
        src94 <= 12'hf4d;
        src95 <= 12'h97a;
        src96 <= 12'h1a4;
        src97 <= 12'h96c;
        src98 <= 12'h59d;
        src99 <= 12'h2eb;
        src100 <= 12'h500;
        src101 <= 12'hdc3;
        src102 <= 12'h9d8;
        src103 <= 12'h6c5;
        src104 <= 12'h87b;
        src105 <= 12'h89b;
        src106 <= 12'hf00;
        src107 <= 12'h407;
        src108 <= 12'hecc;
        src109 <= 12'hc8;
        src110 <= 12'h226;
        src111 <= 12'hfc3;
        src112 <= 12'hd3b;
        src113 <= 12'h7bc;
        src114 <= 12'h10d;
        src115 <= 12'h720;
        src116 <= 12'h83e;
        src117 <= 12'h52e;
        src118 <= 12'he76;
        src119 <= 12'h8ea;
        src120 <= 12'h2c0;
        src121 <= 12'hb43;
        src122 <= 12'h219;
        src123 <= 12'hf08;
        src124 <= 12'hfed;
        src125 <= 12'h1e1;
        src126 <= 12'hd6a;
        src127 <= 12'hf16;
        exp <= 19'h408d6;
        #1
        src0 <= 12'h1ed;
        src1 <= 12'ha49;
        src2 <= 12'h96c;
        src3 <= 12'hb2a;
        src4 <= 12'h9cb;
        src5 <= 12'h8e2;
        src6 <= 12'hf79;
        src7 <= 12'hf45;
        src8 <= 12'hc2a;
        src9 <= 12'h6db;
        src10 <= 12'hf06;
        src11 <= 12'h796;
        src12 <= 12'h603;
        src13 <= 12'hff5;
        src14 <= 12'h894;
        src15 <= 12'h91a;
        src16 <= 12'h3ba;
        src17 <= 12'hd;
        src18 <= 12'hd8c;
        src19 <= 12'h10f;
        src20 <= 12'h892;
        src21 <= 12'h71c;
        src22 <= 12'hc84;
        src23 <= 12'h2f5;
        src24 <= 12'hb1e;
        src25 <= 12'hd75;
        src26 <= 12'h892;
        src27 <= 12'h10f;
        src28 <= 12'hf98;
        src29 <= 12'h80f;
        src30 <= 12'h2ef;
        src31 <= 12'hd0;
        src32 <= 12'h947;
        src33 <= 12'hba8;
        src34 <= 12'h87a;
        src35 <= 12'h211;
        src36 <= 12'hcd6;
        src37 <= 12'h95a;
        src38 <= 12'hec4;
        src39 <= 12'h68b;
        src40 <= 12'h672;
        src41 <= 12'hb80;
        src42 <= 12'hdcc;
        src43 <= 12'h89e;
        src44 <= 12'he98;
        src45 <= 12'h2e5;
        src46 <= 12'h285;
        src47 <= 12'h556;
        src48 <= 12'he56;
        src49 <= 12'hbd6;
        src50 <= 12'h95d;
        src51 <= 12'he43;
        src52 <= 12'h656;
        src53 <= 12'h48e;
        src54 <= 12'he9a;
        src55 <= 12'h2a3;
        src56 <= 12'h8c9;
        src57 <= 12'h547;
        src58 <= 12'he0c;
        src59 <= 12'h2f0;
        src60 <= 12'h5e9;
        src61 <= 12'h93f;
        src62 <= 12'h705;
        src63 <= 12'h5da;
        src64 <= 12'ha3e;
        src65 <= 12'h9de;
        src66 <= 12'h581;
        src67 <= 12'h2bb;
        src68 <= 12'h409;
        src69 <= 12'hf42;
        src70 <= 12'heea;
        src71 <= 12'hbe9;
        src72 <= 12'he2f;
        src73 <= 12'h40a;
        src74 <= 12'hbcf;
        src75 <= 12'h49b;
        src76 <= 12'hd7c;
        src77 <= 12'h7e4;
        src78 <= 12'h514;
        src79 <= 12'hebc;
        src80 <= 12'h926;
        src81 <= 12'haa4;
        src82 <= 12'h419;
        src83 <= 12'h978;
        src84 <= 12'h1d5;
        src85 <= 12'h35e;
        src86 <= 12'h8a2;
        src87 <= 12'h1f1;
        src88 <= 12'h846;
        src89 <= 12'hfb5;
        src90 <= 12'h175;
        src91 <= 12'h379;
        src92 <= 12'h222;
        src93 <= 12'h6a9;
        src94 <= 12'hd1a;
        src95 <= 12'h59b;
        src96 <= 12'h328;
        src97 <= 12'hba2;
        src98 <= 12'h2fb;
        src99 <= 12'hb23;
        src100 <= 12'h489;
        src101 <= 12'had1;
        src102 <= 12'h679;
        src103 <= 12'hb66;
        src104 <= 12'h77c;
        src105 <= 12'hdab;
        src106 <= 12'heb0;
        src107 <= 12'ha23;
        src108 <= 12'hff5;
        src109 <= 12'h35d;
        src110 <= 12'h472;
        src111 <= 12'hc2;
        src112 <= 12'hd8f;
        src113 <= 12'h444;
        src114 <= 12'h5f3;
        src115 <= 12'h638;
        src116 <= 12'h837;
        src117 <= 12'hccd;
        src118 <= 12'hd84;
        src119 <= 12'h84b;
        src120 <= 12'h9d4;
        src121 <= 12'h758;
        src122 <= 12'hbfa;
        src123 <= 12'he52;
        src124 <= 12'hda4;
        src125 <= 12'h513;
        src126 <= 12'h979;
        src127 <= 12'h4b2;
        exp <= 19'h441ed;
        #1
        src0 <= 12'h227;
        src1 <= 12'hc93;
        src2 <= 12'h4a5;
        src3 <= 12'hef7;
        src4 <= 12'h9f5;
        src5 <= 12'h776;
        src6 <= 12'h64;
        src7 <= 12'h87d;
        src8 <= 12'h385;
        src9 <= 12'he0f;
        src10 <= 12'hae;
        src11 <= 12'h60e;
        src12 <= 12'hcc4;
        src13 <= 12'he6;
        src14 <= 12'h349;
        src15 <= 12'h703;
        src16 <= 12'h83d;
        src17 <= 12'hff8;
        src18 <= 12'ha19;
        src19 <= 12'hed0;
        src20 <= 12'h3c4;
        src21 <= 12'h7b2;
        src22 <= 12'h5da;
        src23 <= 12'h1f4;
        src24 <= 12'h550;
        src25 <= 12'h678;
        src26 <= 12'hd9b;
        src27 <= 12'hd60;
        src28 <= 12'h385;
        src29 <= 12'h2fa;
        src30 <= 12'h1c9;
        src31 <= 12'h1f0;
        src32 <= 12'h8a1;
        src33 <= 12'h4c5;
        src34 <= 12'h7e1;
        src35 <= 12'h27e;
        src36 <= 12'hceb;
        src37 <= 12'hf35;
        src38 <= 12'h638;
        src39 <= 12'h688;
        src40 <= 12'h5fe;
        src41 <= 12'h2ac;
        src42 <= 12'h5cb;
        src43 <= 12'h348;
        src44 <= 12'h418;
        src45 <= 12'h7ca;
        src46 <= 12'hf60;
        src47 <= 12'h159;
        src48 <= 12'hc03;
        src49 <= 12'ha64;
        src50 <= 12'hac3;
        src51 <= 12'hc4f;
        src52 <= 12'h9d3;
        src53 <= 12'hc0e;
        src54 <= 12'h85c;
        src55 <= 12'h936;
        src56 <= 12'h6fc;
        src57 <= 12'h937;
        src58 <= 12'h6a9;
        src59 <= 12'h71c;
        src60 <= 12'h1e2;
        src61 <= 12'h3a1;
        src62 <= 12'he73;
        src63 <= 12'hde7;
        src64 <= 12'h389;
        src65 <= 12'h2b0;
        src66 <= 12'hfed;
        src67 <= 12'hc83;
        src68 <= 12'h49e;
        src69 <= 12'hfc0;
        src70 <= 12'haca;
        src71 <= 12'h149;
        src72 <= 12'h5b8;
        src73 <= 12'h79b;
        src74 <= 12'hbe7;
        src75 <= 12'hd8a;
        src76 <= 12'h916;
        src77 <= 12'h609;
        src78 <= 12'h76e;
        src79 <= 12'hf6f;
        src80 <= 12'h7ee;
        src81 <= 12'h969;
        src82 <= 12'h9ed;
        src83 <= 12'ha5d;
        src84 <= 12'h629;
        src85 <= 12'hde7;
        src86 <= 12'ha06;
        src87 <= 12'hf45;
        src88 <= 12'h741;
        src89 <= 12'he56;
        src90 <= 12'heaa;
        src91 <= 12'hd6d;
        src92 <= 12'h820;
        src93 <= 12'h369;
        src94 <= 12'hd6a;
        src95 <= 12'h9af;
        src96 <= 12'h398;
        src97 <= 12'h17c;
        src98 <= 12'hd27;
        src99 <= 12'h6bd;
        src100 <= 12'h8e5;
        src101 <= 12'h2bf;
        src102 <= 12'hdc8;
        src103 <= 12'h7a9;
        src104 <= 12'he61;
        src105 <= 12'hc90;
        src106 <= 12'h543;
        src107 <= 12'hc43;
        src108 <= 12'hf4;
        src109 <= 12'h6a9;
        src110 <= 12'haa5;
        src111 <= 12'h64e;
        src112 <= 12'hfca;
        src113 <= 12'h237;
        src114 <= 12'h8e9;
        src115 <= 12'hd87;
        src116 <= 12'h76;
        src117 <= 12'hd3f;
        src118 <= 12'h414;
        src119 <= 12'hd1a;
        src120 <= 12'h9fd;
        src121 <= 12'h51f;
        src122 <= 12'h93f;
        src123 <= 12'h5b1;
        src124 <= 12'h8c5;
        src125 <= 12'ha40;
        src126 <= 12'hf70;
        src127 <= 12'hdc9;
        exp <= 19'h431db;
        #1
        src0 <= 12'hedf;
        src1 <= 12'hc3;
        src2 <= 12'h402;
        src3 <= 12'h8fa;
        src4 <= 12'hd69;
        src5 <= 12'ha5a;
        src6 <= 12'hc5;
        src7 <= 12'h996;
        src8 <= 12'h8af;
        src9 <= 12'h216;
        src10 <= 12'h3af;
        src11 <= 12'h767;
        src12 <= 12'h3e6;
        src13 <= 12'hcc5;
        src14 <= 12'h9f2;
        src15 <= 12'h12;
        src16 <= 12'h13a;
        src17 <= 12'h371;
        src18 <= 12'h406;
        src19 <= 12'hbdd;
        src20 <= 12'h511;
        src21 <= 12'h404;
        src22 <= 12'h19b;
        src23 <= 12'h5e8;
        src24 <= 12'h335;
        src25 <= 12'h98a;
        src26 <= 12'h73f;
        src27 <= 12'hf74;
        src28 <= 12'h8a8;
        src29 <= 12'hb2b;
        src30 <= 12'h6d2;
        src31 <= 12'h49b;
        src32 <= 12'h2e;
        src33 <= 12'h20;
        src34 <= 12'h616;
        src35 <= 12'hb06;
        src36 <= 12'hd4b;
        src37 <= 12'h82b;
        src38 <= 12'h11a;
        src39 <= 12'hc56;
        src40 <= 12'hec9;
        src41 <= 12'h5a6;
        src42 <= 12'h4ad;
        src43 <= 12'ha82;
        src44 <= 12'he10;
        src45 <= 12'h6bd;
        src46 <= 12'hd57;
        src47 <= 12'h905;
        src48 <= 12'hb4e;
        src49 <= 12'h711;
        src50 <= 12'h5f4;
        src51 <= 12'h165;
        src52 <= 12'hd52;
        src53 <= 12'hb46;
        src54 <= 12'hb2b;
        src55 <= 12'hc84;
        src56 <= 12'h834;
        src57 <= 12'h82b;
        src58 <= 12'h323;
        src59 <= 12'h1b5;
        src60 <= 12'h580;
        src61 <= 12'hc11;
        src62 <= 12'h7ac;
        src63 <= 12'h603;
        src64 <= 12'h769;
        src65 <= 12'h662;
        src66 <= 12'h550;
        src67 <= 12'hd83;
        src68 <= 12'hcc;
        src69 <= 12'h53b;
        src70 <= 12'hb5;
        src71 <= 12'h6a3;
        src72 <= 12'h268;
        src73 <= 12'ha4e;
        src74 <= 12'hc47;
        src75 <= 12'h8a7;
        src76 <= 12'h7e7;
        src77 <= 12'hb97;
        src78 <= 12'h41f;
        src79 <= 12'hcbb;
        src80 <= 12'h57c;
        src81 <= 12'h68;
        src82 <= 12'h37d;
        src83 <= 12'h8a6;
        src84 <= 12'hca0;
        src85 <= 12'h85b;
        src86 <= 12'hed1;
        src87 <= 12'hd13;
        src88 <= 12'h71f;
        src89 <= 12'h5e8;
        src90 <= 12'h7;
        src91 <= 12'hefd;
        src92 <= 12'hf3b;
        src93 <= 12'h95f;
        src94 <= 12'h23b;
        src95 <= 12'hfb2;
        src96 <= 12'hff;
        src97 <= 12'h994;
        src98 <= 12'hfe5;
        src99 <= 12'h168;
        src100 <= 12'h765;
        src101 <= 12'h4b9;
        src102 <= 12'hd63;
        src103 <= 12'hb3f;
        src104 <= 12'h140;
        src105 <= 12'hbc1;
        src106 <= 12'hf6f;
        src107 <= 12'h97a;
        src108 <= 12'h1c9;
        src109 <= 12'h57;
        src110 <= 12'h5f0;
        src111 <= 12'hcc7;
        src112 <= 12'ha1b;
        src113 <= 12'h1fe;
        src114 <= 12'h385;
        src115 <= 12'h586;
        src116 <= 12'h3ac;
        src117 <= 12'h697;
        src118 <= 12'h6d4;
        src119 <= 12'h5b7;
        src120 <= 12'h9f5;
        src121 <= 12'h491;
        src122 <= 12'h246;
        src123 <= 12'hde9;
        src124 <= 12'heaf;
        src125 <= 12'he6f;
        src126 <= 12'haee;
        src127 <= 12'h2a3;
        exp <= 19'h3c6d3;
        #1
        src0 <= 12'h698;
        src1 <= 12'hc9e;
        src2 <= 12'hdcf;
        src3 <= 12'h304;
        src4 <= 12'hb27;
        src5 <= 12'h5a7;
        src6 <= 12'h1be;
        src7 <= 12'h5db;
        src8 <= 12'h957;
        src9 <= 12'hc6a;
        src10 <= 12'h33e;
        src11 <= 12'h423;
        src12 <= 12'h740;
        src13 <= 12'h312;
        src14 <= 12'hd09;
        src15 <= 12'he6a;
        src16 <= 12'h52a;
        src17 <= 12'hc05;
        src18 <= 12'h7d8;
        src19 <= 12'he64;
        src20 <= 12'h8c2;
        src21 <= 12'hb4c;
        src22 <= 12'h678;
        src23 <= 12'hb89;
        src24 <= 12'h5c4;
        src25 <= 12'hd5a;
        src26 <= 12'h9ff;
        src27 <= 12'h644;
        src28 <= 12'hfdf;
        src29 <= 12'hd69;
        src30 <= 12'hdac;
        src31 <= 12'hdd4;
        src32 <= 12'h19b;
        src33 <= 12'hbdb;
        src34 <= 12'h3c7;
        src35 <= 12'hfb7;
        src36 <= 12'h3c;
        src37 <= 12'h270;
        src38 <= 12'h2cb;
        src39 <= 12'hbff;
        src40 <= 12'h565;
        src41 <= 12'ha5;
        src42 <= 12'h5ee;
        src43 <= 12'h7ad;
        src44 <= 12'h5eb;
        src45 <= 12'he30;
        src46 <= 12'hab3;
        src47 <= 12'had8;
        src48 <= 12'hbe7;
        src49 <= 12'h582;
        src50 <= 12'hab6;
        src51 <= 12'h178;
        src52 <= 12'h46f;
        src53 <= 12'hd1a;
        src54 <= 12'hff2;
        src55 <= 12'hd1d;
        src56 <= 12'h9da;
        src57 <= 12'hb7d;
        src58 <= 12'h757;
        src59 <= 12'h62b;
        src60 <= 12'h1bd;
        src61 <= 12'h448;
        src62 <= 12'hb2c;
        src63 <= 12'h9cf;
        src64 <= 12'h711;
        src65 <= 12'h3b6;
        src66 <= 12'h27a;
        src67 <= 12'h12f;
        src68 <= 12'h671;
        src69 <= 12'h3d4;
        src70 <= 12'h319;
        src71 <= 12'h33b;
        src72 <= 12'h388;
        src73 <= 12'h8c6;
        src74 <= 12'h74c;
        src75 <= 12'hc6;
        src76 <= 12'hb4b;
        src77 <= 12'h7cf;
        src78 <= 12'he9a;
        src79 <= 12'hdee;
        src80 <= 12'h6e0;
        src81 <= 12'h91e;
        src82 <= 12'h3b0;
        src83 <= 12'h40c;
        src84 <= 12'h7a9;
        src85 <= 12'haf6;
        src86 <= 12'h2b5;
        src87 <= 12'hc40;
        src88 <= 12'h58f;
        src89 <= 12'h47e;
        src90 <= 12'haf5;
        src91 <= 12'hec3;
        src92 <= 12'h8fe;
        src93 <= 12'h529;
        src94 <= 12'h148;
        src95 <= 12'h4dd;
        src96 <= 12'h826;
        src97 <= 12'h297;
        src98 <= 12'hff0;
        src99 <= 12'h944;
        src100 <= 12'hcda;
        src101 <= 12'h98a;
        src102 <= 12'h7cd;
        src103 <= 12'h552;
        src104 <= 12'h26f;
        src105 <= 12'hc46;
        src106 <= 12'hbe4;
        src107 <= 12'h3ff;
        src108 <= 12'hd2a;
        src109 <= 12'ha1d;
        src110 <= 12'h629;
        src111 <= 12'hf32;
        src112 <= 12'hd35;
        src113 <= 12'h2a6;
        src114 <= 12'h5f6;
        src115 <= 12'hc9f;
        src116 <= 12'h585;
        src117 <= 12'h979;
        src118 <= 12'hda5;
        src119 <= 12'hebc;
        src120 <= 12'h1b;
        src121 <= 12'hc84;
        src122 <= 12'h37c;
        src123 <= 12'h853;
        src124 <= 12'hb0;
        src125 <= 12'he5f;
        src126 <= 12'h49a;
        src127 <= 12'h86f;
        exp <= 19'h40c24;
        #1
        src0 <= 12'ha67;
        src1 <= 12'h3fc;
        src2 <= 12'h25e;
        src3 <= 12'h592;
        src4 <= 12'h1e3;
        src5 <= 12'h24d;
        src6 <= 12'h3c2;
        src7 <= 12'hcf2;
        src8 <= 12'hf79;
        src9 <= 12'h286;
        src10 <= 12'hf34;
        src11 <= 12'h978;
        src12 <= 12'hc65;
        src13 <= 12'h5f9;
        src14 <= 12'h5b2;
        src15 <= 12'h1c;
        src16 <= 12'h9cc;
        src17 <= 12'hac9;
        src18 <= 12'h378;
        src19 <= 12'h303;
        src20 <= 12'h964;
        src21 <= 12'h1c1;
        src22 <= 12'hc6b;
        src23 <= 12'h88e;
        src24 <= 12'hdaf;
        src25 <= 12'hcfb;
        src26 <= 12'h58;
        src27 <= 12'h7aa;
        src28 <= 12'h6e1;
        src29 <= 12'h9e;
        src30 <= 12'ha0d;
        src31 <= 12'had3;
        src32 <= 12'h6c1;
        src33 <= 12'ha9d;
        src34 <= 12'hecf;
        src35 <= 12'h212;
        src36 <= 12'h620;
        src37 <= 12'h731;
        src38 <= 12'haa6;
        src39 <= 12'h43d;
        src40 <= 12'h285;
        src41 <= 12'h870;
        src42 <= 12'h9ce;
        src43 <= 12'h55e;
        src44 <= 12'h16a;
        src45 <= 12'he5f;
        src46 <= 12'hcba;
        src47 <= 12'h9c0;
        src48 <= 12'h8c;
        src49 <= 12'h690;
        src50 <= 12'hb90;
        src51 <= 12'h3fb;
        src52 <= 12'haa8;
        src53 <= 12'heed;
        src54 <= 12'h638;
        src55 <= 12'h2e2;
        src56 <= 12'hf63;
        src57 <= 12'h883;
        src58 <= 12'h958;
        src59 <= 12'h9ae;
        src60 <= 12'hd92;
        src61 <= 12'h4c5;
        src62 <= 12'h24a;
        src63 <= 12'h705;
        src64 <= 12'hf21;
        src65 <= 12'h1cf;
        src66 <= 12'h706;
        src67 <= 12'h256;
        src68 <= 12'hc72;
        src69 <= 12'hd08;
        src70 <= 12'h474;
        src71 <= 12'h3a6;
        src72 <= 12'h197;
        src73 <= 12'h217;
        src74 <= 12'h524;
        src75 <= 12'h3b5;
        src76 <= 12'h8ed;
        src77 <= 12'h8e3;
        src78 <= 12'h7b9;
        src79 <= 12'hc54;
        src80 <= 12'h306;
        src81 <= 12'h50e;
        src82 <= 12'hd13;
        src83 <= 12'h7ce;
        src84 <= 12'hb39;
        src85 <= 12'h55a;
        src86 <= 12'h5a2;
        src87 <= 12'haa5;
        src88 <= 12'hd06;
        src89 <= 12'h30e;
        src90 <= 12'h9c9;
        src91 <= 12'he2c;
        src92 <= 12'hea1;
        src93 <= 12'h755;
        src94 <= 12'hebe;
        src95 <= 12'h43a;
        src96 <= 12'h7fd;
        src97 <= 12'h8c8;
        src98 <= 12'hc3e;
        src99 <= 12'h770;
        src100 <= 12'h1cc;
        src101 <= 12'h900;
        src102 <= 12'hdc6;
        src103 <= 12'h7f1;
        src104 <= 12'ha08;
        src105 <= 12'hd06;
        src106 <= 12'h75;
        src107 <= 12'h483;
        src108 <= 12'h569;
        src109 <= 12'h526;
        src110 <= 12'h17a;
        src111 <= 12'h54b;
        src112 <= 12'h71b;
        src113 <= 12'ha8c;
        src114 <= 12'h22f;
        src115 <= 12'hbbf;
        src116 <= 12'hbc0;
        src117 <= 12'h828;
        src118 <= 12'h117;
        src119 <= 12'h8c0;
        src120 <= 12'h466;
        src121 <= 12'ha1d;
        src122 <= 12'h4e2;
        src123 <= 12'hcba;
        src124 <= 12'h562;
        src125 <= 12'h67e;
        src126 <= 12'hf5f;
        src127 <= 12'h17;
        exp <= 19'h3cf29;
        #1
        src0 <= 12'h694;
        src1 <= 12'h4b4;
        src2 <= 12'h195;
        src3 <= 12'h5b8;
        src4 <= 12'h6f5;
        src5 <= 12'h9f9;
        src6 <= 12'he6e;
        src7 <= 12'h880;
        src8 <= 12'heed;
        src9 <= 12'h1d6;
        src10 <= 12'hd38;
        src11 <= 12'hd40;
        src12 <= 12'h24d;
        src13 <= 12'h644;
        src14 <= 12'h375;
        src15 <= 12'h59;
        src16 <= 12'hd6f;
        src17 <= 12'h44;
        src18 <= 12'h5a7;
        src19 <= 12'h841;
        src20 <= 12'h78a;
        src21 <= 12'hbfb;
        src22 <= 12'hc00;
        src23 <= 12'h828;
        src24 <= 12'hf4f;
        src25 <= 12'ha2a;
        src26 <= 12'h35e;
        src27 <= 12'hb80;
        src28 <= 12'h938;
        src29 <= 12'h3ce;
        src30 <= 12'h775;
        src31 <= 12'hb4f;
        src32 <= 12'h509;
        src33 <= 12'h37d;
        src34 <= 12'ha79;
        src35 <= 12'he6c;
        src36 <= 12'hb79;
        src37 <= 12'hdaf;
        src38 <= 12'h91a;
        src39 <= 12'h9be;
        src40 <= 12'hb3b;
        src41 <= 12'h71;
        src42 <= 12'h72e;
        src43 <= 12'h465;
        src44 <= 12'h97d;
        src45 <= 12'h29b;
        src46 <= 12'h6de;
        src47 <= 12'h2d8;
        src48 <= 12'h268;
        src49 <= 12'he7e;
        src50 <= 12'h7eb;
        src51 <= 12'h190;
        src52 <= 12'hb03;
        src53 <= 12'h370;
        src54 <= 12'h4aa;
        src55 <= 12'h1e7;
        src56 <= 12'h9e8;
        src57 <= 12'h448;
        src58 <= 12'h7ff;
        src59 <= 12'h8c3;
        src60 <= 12'hfee;
        src61 <= 12'ha8d;
        src62 <= 12'he11;
        src63 <= 12'hd86;
        src64 <= 12'he38;
        src65 <= 12'h8ce;
        src66 <= 12'hf8b;
        src67 <= 12'h20e;
        src68 <= 12'heb0;
        src69 <= 12'he32;
        src70 <= 12'hd34;
        src71 <= 12'h3f2;
        src72 <= 12'h3b6;
        src73 <= 12'h95b;
        src74 <= 12'he32;
        src75 <= 12'h98c;
        src76 <= 12'h3d1;
        src77 <= 12'h1d9;
        src78 <= 12'hd83;
        src79 <= 12'h446;
        src80 <= 12'h63e;
        src81 <= 12'h11a;
        src82 <= 12'h1a4;
        src83 <= 12'hac7;
        src84 <= 12'h87e;
        src85 <= 12'h849;
        src86 <= 12'h35b;
        src87 <= 12'h345;
        src88 <= 12'hb89;
        src89 <= 12'hf4c;
        src90 <= 12'hda;
        src91 <= 12'hce2;
        src92 <= 12'ha55;
        src93 <= 12'h2ec;
        src94 <= 12'hf21;
        src95 <= 12'h67a;
        src96 <= 12'hc47;
        src97 <= 12'h655;
        src98 <= 12'hdff;
        src99 <= 12'h81d;
        src100 <= 12'h35c;
        src101 <= 12'h850;
        src102 <= 12'h59f;
        src103 <= 12'hae2;
        src104 <= 12'h6b4;
        src105 <= 12'h465;
        src106 <= 12'hc7f;
        src107 <= 12'heb8;
        src108 <= 12'h692;
        src109 <= 12'hb6b;
        src110 <= 12'hbf9;
        src111 <= 12'he41;
        src112 <= 12'hae4;
        src113 <= 12'h892;
        src114 <= 12'he47;
        src115 <= 12'hbf7;
        src116 <= 12'hda4;
        src117 <= 12'hcbb;
        src118 <= 12'hb1d;
        src119 <= 12'h773;
        src120 <= 12'h7b5;
        src121 <= 12'hb22;
        src122 <= 12'h2dc;
        src123 <= 12'h956;
        src124 <= 12'h1b4;
        src125 <= 12'h9bb;
        src126 <= 12'h820;
        src127 <= 12'h168;
        exp <= 19'h42be4;
        #1
        src0 <= 12'h551;
        src1 <= 12'h263;
        src2 <= 12'h284;
        src3 <= 12'h116;
        src4 <= 12'he12;
        src5 <= 12'ha08;
        src6 <= 12'h7c;
        src7 <= 12'hef3;
        src8 <= 12'h7ec;
        src9 <= 12'hd2a;
        src10 <= 12'h8a6;
        src11 <= 12'h896;
        src12 <= 12'h907;
        src13 <= 12'h88e;
        src14 <= 12'h822;
        src15 <= 12'h252;
        src16 <= 12'hf71;
        src17 <= 12'he04;
        src18 <= 12'hd68;
        src19 <= 12'h9a2;
        src20 <= 12'h94e;
        src21 <= 12'hb7b;
        src22 <= 12'h4c1;
        src23 <= 12'hdc4;
        src24 <= 12'h377;
        src25 <= 12'hb45;
        src26 <= 12'h5f6;
        src27 <= 12'h4f8;
        src28 <= 12'h7ee;
        src29 <= 12'h72c;
        src30 <= 12'hb23;
        src31 <= 12'hb8f;
        src32 <= 12'h5ac;
        src33 <= 12'h896;
        src34 <= 12'h28e;
        src35 <= 12'h46b;
        src36 <= 12'hae7;
        src37 <= 12'h58c;
        src38 <= 12'hd76;
        src39 <= 12'h1ea;
        src40 <= 12'h38e;
        src41 <= 12'h243;
        src42 <= 12'h9d6;
        src43 <= 12'h1dc;
        src44 <= 12'h152;
        src45 <= 12'h88e;
        src46 <= 12'hadc;
        src47 <= 12'h19a;
        src48 <= 12'hc52;
        src49 <= 12'he0a;
        src50 <= 12'h945;
        src51 <= 12'h8c;
        src52 <= 12'h260;
        src53 <= 12'ha3e;
        src54 <= 12'h8a0;
        src55 <= 12'h61;
        src56 <= 12'h61b;
        src57 <= 12'hc7b;
        src58 <= 12'hdf6;
        src59 <= 12'h5d2;
        src60 <= 12'h225;
        src61 <= 12'hd6e;
        src62 <= 12'hfc4;
        src63 <= 12'h22;
        src64 <= 12'h3cb;
        src65 <= 12'h337;
        src66 <= 12'h40c;
        src67 <= 12'h1d6;
        src68 <= 12'h24a;
        src69 <= 12'h8ec;
        src70 <= 12'hada;
        src71 <= 12'h5cb;
        src72 <= 12'hbb6;
        src73 <= 12'hdbe;
        src74 <= 12'hab;
        src75 <= 12'h9f6;
        src76 <= 12'hd8b;
        src77 <= 12'h155;
        src78 <= 12'h828;
        src79 <= 12'hed6;
        src80 <= 12'h236;
        src81 <= 12'hb92;
        src82 <= 12'h18a;
        src83 <= 12'h551;
        src84 <= 12'h77e;
        src85 <= 12'hcdf;
        src86 <= 12'hda5;
        src87 <= 12'hf9d;
        src88 <= 12'ha07;
        src89 <= 12'h135;
        src90 <= 12'h7e0;
        src91 <= 12'h48c;
        src92 <= 12'h8b1;
        src93 <= 12'hccb;
        src94 <= 12'h8ba;
        src95 <= 12'h717;
        src96 <= 12'h83a;
        src97 <= 12'h1b4;
        src98 <= 12'h958;
        src99 <= 12'hebc;
        src100 <= 12'h86b;
        src101 <= 12'hab2;
        src102 <= 12'hdb4;
        src103 <= 12'h1d5;
        src104 <= 12'h8c0;
        src105 <= 12'hf41;
        src106 <= 12'h3ba;
        src107 <= 12'h58c;
        src108 <= 12'h126;
        src109 <= 12'ha74;
        src110 <= 12'hd0d;
        src111 <= 12'hf3e;
        src112 <= 12'ha96;
        src113 <= 12'hfb7;
        src114 <= 12'h694;
        src115 <= 12'h86e;
        src116 <= 12'h32f;
        src117 <= 12'h516;
        src118 <= 12'h102;
        src119 <= 12'h5f4;
        src120 <= 12'h63d;
        src121 <= 12'h7d7;
        src122 <= 12'hac;
        src123 <= 12'hc15;
        src124 <= 12'h89c;
        src125 <= 12'h42d;
        src126 <= 12'h62c;
        src127 <= 12'hba2;
        exp <= 19'h3e2b2;
        #1
        src0 <= 12'h1bc;
        src1 <= 12'h633;
        src2 <= 12'h510;
        src3 <= 12'h256;
        src4 <= 12'hb05;
        src5 <= 12'h501;
        src6 <= 12'h596;
        src7 <= 12'h6be;
        src8 <= 12'hc15;
        src9 <= 12'h1f0;
        src10 <= 12'h2f0;
        src11 <= 12'h501;
        src12 <= 12'h7e4;
        src13 <= 12'h9c8;
        src14 <= 12'he2a;
        src15 <= 12'h23f;
        src16 <= 12'h859;
        src17 <= 12'h4e2;
        src18 <= 12'h235;
        src19 <= 12'h742;
        src20 <= 12'h748;
        src21 <= 12'ha27;
        src22 <= 12'haba;
        src23 <= 12'h324;
        src24 <= 12'h3b8;
        src25 <= 12'h9d3;
        src26 <= 12'h332;
        src27 <= 12'h75;
        src28 <= 12'h7db;
        src29 <= 12'hc04;
        src30 <= 12'h1dc;
        src31 <= 12'ha8b;
        src32 <= 12'h8e6;
        src33 <= 12'hac2;
        src34 <= 12'ha4c;
        src35 <= 12'h46e;
        src36 <= 12'ha80;
        src37 <= 12'hd83;
        src38 <= 12'hd59;
        src39 <= 12'h7e8;
        src40 <= 12'hb7d;
        src41 <= 12'hb19;
        src42 <= 12'h29a;
        src43 <= 12'hcc4;
        src44 <= 12'hddf;
        src45 <= 12'h6a3;
        src46 <= 12'h498;
        src47 <= 12'h588;
        src48 <= 12'h936;
        src49 <= 12'h163;
        src50 <= 12'hf63;
        src51 <= 12'hb78;
        src52 <= 12'heb5;
        src53 <= 12'h5cb;
        src54 <= 12'h87d;
        src55 <= 12'h23d;
        src56 <= 12'ha0;
        src57 <= 12'hc9;
        src58 <= 12'hd88;
        src59 <= 12'hba1;
        src60 <= 12'hf6a;
        src61 <= 12'hce7;
        src62 <= 12'hd4b;
        src63 <= 12'he65;
        src64 <= 12'h105;
        src65 <= 12'h3b4;
        src66 <= 12'h88d;
        src67 <= 12'h840;
        src68 <= 12'hec4;
        src69 <= 12'hdb7;
        src70 <= 12'h2d5;
        src71 <= 12'hcaa;
        src72 <= 12'h58c;
        src73 <= 12'h635;
        src74 <= 12'h903;
        src75 <= 12'h206;
        src76 <= 12'hdcf;
        src77 <= 12'h657;
        src78 <= 12'h909;
        src79 <= 12'hf6e;
        src80 <= 12'h965;
        src81 <= 12'h472;
        src82 <= 12'h313;
        src83 <= 12'he7d;
        src84 <= 12'h11e;
        src85 <= 12'hece;
        src86 <= 12'hb54;
        src87 <= 12'hfdc;
        src88 <= 12'h79b;
        src89 <= 12'h21e;
        src90 <= 12'h2be;
        src91 <= 12'h6f0;
        src92 <= 12'h1d5;
        src93 <= 12'h55a;
        src94 <= 12'h503;
        src95 <= 12'he77;
        src96 <= 12'hc04;
        src97 <= 12'h90c;
        src98 <= 12'he43;
        src99 <= 12'h695;
        src100 <= 12'h4f0;
        src101 <= 12'h92;
        src102 <= 12'h1f8;
        src103 <= 12'h333;
        src104 <= 12'hd60;
        src105 <= 12'hd91;
        src106 <= 12'h342;
        src107 <= 12'h39f;
        src108 <= 12'ha88;
        src109 <= 12'haed;
        src110 <= 12'h559;
        src111 <= 12'h8b7;
        src112 <= 12'hbfd;
        src113 <= 12'hdd;
        src114 <= 12'h156;
        src115 <= 12'h683;
        src116 <= 12'hf67;
        src117 <= 12'hca2;
        src118 <= 12'hdc4;
        src119 <= 12'hb3d;
        src120 <= 12'ha8e;
        src121 <= 12'hf04;
        src122 <= 12'hcd0;
        src123 <= 12'hd69;
        src124 <= 12'hd5;
        src125 <= 12'h47a;
        src126 <= 12'h47b;
        src127 <= 12'h69;
        exp <= 19'h3f5cf;
        #1
        src0 <= 12'h3b;
        src1 <= 12'h8b3;
        src2 <= 12'h8c7;
        src3 <= 12'h695;
        src4 <= 12'hd92;
        src5 <= 12'h101;
        src6 <= 12'hda4;
        src7 <= 12'he3a;
        src8 <= 12'h68;
        src9 <= 12'h570;
        src10 <= 12'h8d2;
        src11 <= 12'h16e;
        src12 <= 12'hf6e;
        src13 <= 12'hf41;
        src14 <= 12'h478;
        src15 <= 12'h74d;
        src16 <= 12'hf80;
        src17 <= 12'hd47;
        src18 <= 12'h90f;
        src19 <= 12'h288;
        src20 <= 12'h819;
        src21 <= 12'h9cf;
        src22 <= 12'h50a;
        src23 <= 12'h32a;
        src24 <= 12'hc8d;
        src25 <= 12'h8eb;
        src26 <= 12'h112;
        src27 <= 12'h25a;
        src28 <= 12'h528;
        src29 <= 12'h59;
        src30 <= 12'hdb6;
        src31 <= 12'h544;
        src32 <= 12'hd45;
        src33 <= 12'h552;
        src34 <= 12'hc4d;
        src35 <= 12'h28c;
        src36 <= 12'hf52;
        src37 <= 12'h903;
        src38 <= 12'hb56;
        src39 <= 12'he9c;
        src40 <= 12'h4b;
        src41 <= 12'haef;
        src42 <= 12'hb3b;
        src43 <= 12'h67b;
        src44 <= 12'hf4d;
        src45 <= 12'h50d;
        src46 <= 12'hcb7;
        src47 <= 12'h68e;
        src48 <= 12'hb5b;
        src49 <= 12'hfc1;
        src50 <= 12'h5b2;
        src51 <= 12'h151;
        src52 <= 12'hd31;
        src53 <= 12'h4f2;
        src54 <= 12'hac9;
        src55 <= 12'h390;
        src56 <= 12'h1d4;
        src57 <= 12'h11a;
        src58 <= 12'h363;
        src59 <= 12'ha0d;
        src60 <= 12'hc61;
        src61 <= 12'h74a;
        src62 <= 12'hd0c;
        src63 <= 12'hb5a;
        src64 <= 12'h3c9;
        src65 <= 12'ha28;
        src66 <= 12'h969;
        src67 <= 12'h598;
        src68 <= 12'hc85;
        src69 <= 12'h70;
        src70 <= 12'h758;
        src71 <= 12'h747;
        src72 <= 12'hd49;
        src73 <= 12'hdc6;
        src74 <= 12'h202;
        src75 <= 12'h20e;
        src76 <= 12'ha84;
        src77 <= 12'hec9;
        src78 <= 12'h69b;
        src79 <= 12'h506;
        src80 <= 12'h3c6;
        src81 <= 12'h6b3;
        src82 <= 12'hc37;
        src83 <= 12'hfab;
        src84 <= 12'h2b1;
        src85 <= 12'h406;
        src86 <= 12'h35e;
        src87 <= 12'h33;
        src88 <= 12'h8be;
        src89 <= 12'h5ea;
        src90 <= 12'h9dc;
        src91 <= 12'ha03;
        src92 <= 12'hefe;
        src93 <= 12'hae1;
        src94 <= 12'hb75;
        src95 <= 12'h473;
        src96 <= 12'h21b;
        src97 <= 12'hb6a;
        src98 <= 12'h967;
        src99 <= 12'h94b;
        src100 <= 12'h2ec;
        src101 <= 12'h122;
        src102 <= 12'hd4e;
        src103 <= 12'hee6;
        src104 <= 12'he32;
        src105 <= 12'h27e;
        src106 <= 12'h5e9;
        src107 <= 12'h1de;
        src108 <= 12'hd1a;
        src109 <= 12'hc4f;
        src110 <= 12'hfce;
        src111 <= 12'he2f;
        src112 <= 12'h95f;
        src113 <= 12'h228;
        src114 <= 12'hb38;
        src115 <= 12'h662;
        src116 <= 12'hf2e;
        src117 <= 12'h33d;
        src118 <= 12'h8da;
        src119 <= 12'hb5f;
        src120 <= 12'hb7c;
        src121 <= 12'h698;
        src122 <= 12'h23;
        src123 <= 12'h3f;
        src124 <= 12'ha4;
        src125 <= 12'hfd8;
        src126 <= 12'h356;
        src127 <= 12'hce6;
        exp <= 19'h4093d;
        #1
        src0 <= 12'hc37;
        src1 <= 12'h2c7;
        src2 <= 12'h76e;
        src3 <= 12'h3b9;
        src4 <= 12'hbf4;
        src5 <= 12'h1d1;
        src6 <= 12'h6cf;
        src7 <= 12'h6d3;
        src8 <= 12'h7af;
        src9 <= 12'h9c5;
        src10 <= 12'h212;
        src11 <= 12'hb4b;
        src12 <= 12'hf1a;
        src13 <= 12'hd4f;
        src14 <= 12'hc32;
        src15 <= 12'h7b5;
        src16 <= 12'h2c;
        src17 <= 12'hd56;
        src18 <= 12'h960;
        src19 <= 12'h69a;
        src20 <= 12'hbe0;
        src21 <= 12'hd5f;
        src22 <= 12'he7d;
        src23 <= 12'h5fc;
        src24 <= 12'h1be;
        src25 <= 12'ha08;
        src26 <= 12'h514;
        src27 <= 12'h764;
        src28 <= 12'h3b;
        src29 <= 12'hc4f;
        src30 <= 12'hc7e;
        src31 <= 12'hf9e;
        src32 <= 12'ha0f;
        src33 <= 12'hb4b;
        src34 <= 12'h8cb;
        src35 <= 12'h610;
        src36 <= 12'h93d;
        src37 <= 12'h34a;
        src38 <= 12'ha91;
        src39 <= 12'h5a7;
        src40 <= 12'ha8a;
        src41 <= 12'h9c9;
        src42 <= 12'hb00;
        src43 <= 12'h337;
        src44 <= 12'hc7e;
        src45 <= 12'hfe2;
        src46 <= 12'ha84;
        src47 <= 12'h2ce;
        src48 <= 12'h554;
        src49 <= 12'hb89;
        src50 <= 12'h433;
        src51 <= 12'hbec;
        src52 <= 12'ha9d;
        src53 <= 12'h5a8;
        src54 <= 12'h956;
        src55 <= 12'h544;
        src56 <= 12'h5bf;
        src57 <= 12'h86d;
        src58 <= 12'h122;
        src59 <= 12'hd14;
        src60 <= 12'h47f;
        src61 <= 12'h1e2;
        src62 <= 12'h720;
        src63 <= 12'h2a9;
        src64 <= 12'he92;
        src65 <= 12'h56f;
        src66 <= 12'hb64;
        src67 <= 12'hd8f;
        src68 <= 12'hd73;
        src69 <= 12'h273;
        src70 <= 12'hc7e;
        src71 <= 12'h724;
        src72 <= 12'hed8;
        src73 <= 12'h611;
        src74 <= 12'h6b2;
        src75 <= 12'h712;
        src76 <= 12'hfc1;
        src77 <= 12'hc39;
        src78 <= 12'h11c;
        src79 <= 12'h144;
        src80 <= 12'hf53;
        src81 <= 12'h652;
        src82 <= 12'h5e7;
        src83 <= 12'he4e;
        src84 <= 12'hc58;
        src85 <= 12'h1c7;
        src86 <= 12'haf3;
        src87 <= 12'h70;
        src88 <= 12'h199;
        src89 <= 12'ha0d;
        src90 <= 12'hbb9;
        src91 <= 12'h23a;
        src92 <= 12'h630;
        src93 <= 12'h5e7;
        src94 <= 12'h771;
        src95 <= 12'hca2;
        src96 <= 12'hddd;
        src97 <= 12'he4c;
        src98 <= 12'h2d0;
        src99 <= 12'h92c;
        src100 <= 12'he1;
        src101 <= 12'h63c;
        src102 <= 12'hd;
        src103 <= 12'h690;
        src104 <= 12'hf3a;
        src105 <= 12'h20;
        src106 <= 12'haad;
        src107 <= 12'h554;
        src108 <= 12'hd90;
        src109 <= 12'hb8e;
        src110 <= 12'hd29;
        src111 <= 12'h61;
        src112 <= 12'h649;
        src113 <= 12'hd3a;
        src114 <= 12'hab7;
        src115 <= 12'hc09;
        src116 <= 12'h1c4;
        src117 <= 12'h11;
        src118 <= 12'hd0b;
        src119 <= 12'h252;
        src120 <= 12'hdf0;
        src121 <= 12'hbf1;
        src122 <= 12'he3d;
        src123 <= 12'h797;
        src124 <= 12'hc0a;
        src125 <= 12'hcbe;
        src126 <= 12'h197;
        src127 <= 12'h1d7;
        exp <= 19'h41c40;
        #1
        src0 <= 12'h6fe;
        src1 <= 12'h2d1;
        src2 <= 12'he98;
        src3 <= 12'h39d;
        src4 <= 12'h3a4;
        src5 <= 12'h939;
        src6 <= 12'h3dd;
        src7 <= 12'h701;
        src8 <= 12'ha08;
        src9 <= 12'h9b2;
        src10 <= 12'h549;
        src11 <= 12'h33;
        src12 <= 12'he2c;
        src13 <= 12'h811;
        src14 <= 12'h86c;
        src15 <= 12'h277;
        src16 <= 12'hde1;
        src17 <= 12'hc54;
        src18 <= 12'h937;
        src19 <= 12'haf;
        src20 <= 12'hd81;
        src21 <= 12'h9e1;
        src22 <= 12'h40;
        src23 <= 12'ha25;
        src24 <= 12'h68d;
        src25 <= 12'hff3;
        src26 <= 12'h114;
        src27 <= 12'h464;
        src28 <= 12'h252;
        src29 <= 12'h7cc;
        src30 <= 12'h46f;
        src31 <= 12'hba;
        src32 <= 12'h17d;
        src33 <= 12'h248;
        src34 <= 12'hb70;
        src35 <= 12'h114;
        src36 <= 12'ha47;
        src37 <= 12'hac9;
        src38 <= 12'heed;
        src39 <= 12'h2e4;
        src40 <= 12'h151;
        src41 <= 12'hee4;
        src42 <= 12'h2ee;
        src43 <= 12'hee7;
        src44 <= 12'h5aa;
        src45 <= 12'h456;
        src46 <= 12'hb08;
        src47 <= 12'h3ba;
        src48 <= 12'h1c9;
        src49 <= 12'h998;
        src50 <= 12'h388;
        src51 <= 12'h440;
        src52 <= 12'h3eb;
        src53 <= 12'hcbf;
        src54 <= 12'hb4a;
        src55 <= 12'hdb5;
        src56 <= 12'ha6d;
        src57 <= 12'h2b9;
        src58 <= 12'he1e;
        src59 <= 12'hab1;
        src60 <= 12'h26b;
        src61 <= 12'hb96;
        src62 <= 12'h72e;
        src63 <= 12'h366;
        src64 <= 12'hade;
        src65 <= 12'h7c1;
        src66 <= 12'h718;
        src67 <= 12'h673;
        src68 <= 12'hd7f;
        src69 <= 12'h5c8;
        src70 <= 12'h3fb;
        src71 <= 12'h8da;
        src72 <= 12'h31e;
        src73 <= 12'hc01;
        src74 <= 12'h64d;
        src75 <= 12'h9d2;
        src76 <= 12'h310;
        src77 <= 12'h216;
        src78 <= 12'h240;
        src79 <= 12'h4e6;
        src80 <= 12'h831;
        src81 <= 12'h930;
        src82 <= 12'h6ff;
        src83 <= 12'h15a;
        src84 <= 12'he58;
        src85 <= 12'hbf1;
        src86 <= 12'he54;
        src87 <= 12'h434;
        src88 <= 12'h464;
        src89 <= 12'h9b;
        src90 <= 12'hd9;
        src91 <= 12'hff5;
        src92 <= 12'hdf1;
        src93 <= 12'he71;
        src94 <= 12'h9e2;
        src95 <= 12'h1;
        src96 <= 12'hbbe;
        src97 <= 12'hbe9;
        src98 <= 12'he45;
        src99 <= 12'hf3d;
        src100 <= 12'he33;
        src101 <= 12'hebd;
        src102 <= 12'h5e6;
        src103 <= 12'h5c2;
        src104 <= 12'haae;
        src105 <= 12'haa0;
        src106 <= 12'h235;
        src107 <= 12'hf58;
        src108 <= 12'hf42;
        src109 <= 12'hb45;
        src110 <= 12'h4c;
        src111 <= 12'h5a3;
        src112 <= 12'ha8c;
        src113 <= 12'hd83;
        src114 <= 12'h795;
        src115 <= 12'h1bf;
        src116 <= 12'ha7c;
        src117 <= 12'h926;
        src118 <= 12'h275;
        src119 <= 12'h821;
        src120 <= 12'h673;
        src121 <= 12'h43e;
        src122 <= 12'h8a4;
        src123 <= 12'h104;
        src124 <= 12'h603;
        src125 <= 12'hb2a;
        src126 <= 12'hd50;
        src127 <= 12'h489;
        exp <= 19'h3d701;
        #1
        src0 <= 12'hfe1;
        src1 <= 12'ha;
        src2 <= 12'h68d;
        src3 <= 12'h192;
        src4 <= 12'ha7d;
        src5 <= 12'hdd4;
        src6 <= 12'he77;
        src7 <= 12'ha02;
        src8 <= 12'h4ad;
        src9 <= 12'h730;
        src10 <= 12'h1de;
        src11 <= 12'h936;
        src12 <= 12'h7a;
        src13 <= 12'hde;
        src14 <= 12'he0e;
        src15 <= 12'hbe5;
        src16 <= 12'h208;
        src17 <= 12'h6c9;
        src18 <= 12'h2b4;
        src19 <= 12'h94c;
        src20 <= 12'h5c2;
        src21 <= 12'h20d;
        src22 <= 12'h6f2;
        src23 <= 12'hd79;
        src24 <= 12'h6a7;
        src25 <= 12'h7c0;
        src26 <= 12'h895;
        src27 <= 12'h58f;
        src28 <= 12'hee7;
        src29 <= 12'h812;
        src30 <= 12'h4c9;
        src31 <= 12'hf73;
        src32 <= 12'h50;
        src33 <= 12'h96a;
        src34 <= 12'h6f3;
        src35 <= 12'ha92;
        src36 <= 12'hcdf;
        src37 <= 12'hddc;
        src38 <= 12'hb01;
        src39 <= 12'h5d3;
        src40 <= 12'h496;
        src41 <= 12'h1b3;
        src42 <= 12'h18d;
        src43 <= 12'hddd;
        src44 <= 12'h8bf;
        src45 <= 12'haa;
        src46 <= 12'h7ad;
        src47 <= 12'h1fb;
        src48 <= 12'hf64;
        src49 <= 12'h1c3;
        src50 <= 12'h7b5;
        src51 <= 12'hf5e;
        src52 <= 12'h7fd;
        src53 <= 12'he36;
        src54 <= 12'ha92;
        src55 <= 12'h9e;
        src56 <= 12'hb9e;
        src57 <= 12'h844;
        src58 <= 12'h51e;
        src59 <= 12'h895;
        src60 <= 12'h80c;
        src61 <= 12'h344;
        src62 <= 12'h303;
        src63 <= 12'h8a6;
        src64 <= 12'hcf8;
        src65 <= 12'h877;
        src66 <= 12'hc7f;
        src67 <= 12'h5f5;
        src68 <= 12'h9af;
        src69 <= 12'h489;
        src70 <= 12'hb40;
        src71 <= 12'h3a2;
        src72 <= 12'hc72;
        src73 <= 12'ha5b;
        src74 <= 12'he02;
        src75 <= 12'h60d;
        src76 <= 12'hf24;
        src77 <= 12'h999;
        src78 <= 12'h237;
        src79 <= 12'h980;
        src80 <= 12'hb2d;
        src81 <= 12'he34;
        src82 <= 12'hb70;
        src83 <= 12'h872;
        src84 <= 12'h7ee;
        src85 <= 12'h290;
        src86 <= 12'heb7;
        src87 <= 12'h4ca;
        src88 <= 12'hcc5;
        src89 <= 12'hab;
        src90 <= 12'h975;
        src91 <= 12'hd6;
        src92 <= 12'h734;
        src93 <= 12'hb30;
        src94 <= 12'h143;
        src95 <= 12'hfaf;
        src96 <= 12'hb1e;
        src97 <= 12'h149;
        src98 <= 12'h7d2;
        src99 <= 12'hf0e;
        src100 <= 12'h8de;
        src101 <= 12'he64;
        src102 <= 12'ha12;
        src103 <= 12'h88d;
        src104 <= 12'h88d;
        src105 <= 12'h8c9;
        src106 <= 12'h6f0;
        src107 <= 12'h7ef;
        src108 <= 12'h616;
        src109 <= 12'h14f;
        src110 <= 12'h382;
        src111 <= 12'h20;
        src112 <= 12'hbff;
        src113 <= 12'h175;
        src114 <= 12'h19a;
        src115 <= 12'h44;
        src116 <= 12'h3aa;
        src117 <= 12'h71e;
        src118 <= 12'h696;
        src119 <= 12'h80;
        src120 <= 12'h843;
        src121 <= 12'hbfe;
        src122 <= 12'hfdc;
        src123 <= 12'h501;
        src124 <= 12'h24f;
        src125 <= 12'he2d;
        src126 <= 12'hbb0;
        src127 <= 12'hd07;
        exp <= 19'h3ec1d;
        #1
        src0 <= 12'hb1;
        src1 <= 12'h237;
        src2 <= 12'hccc;
        src3 <= 12'h695;
        src4 <= 12'hb13;
        src5 <= 12'haaf;
        src6 <= 12'hd10;
        src7 <= 12'h45c;
        src8 <= 12'he62;
        src9 <= 12'h272;
        src10 <= 12'h958;
        src11 <= 12'h9d7;
        src12 <= 12'hbc1;
        src13 <= 12'h181;
        src14 <= 12'h612;
        src15 <= 12'ha49;
        src16 <= 12'ha15;
        src17 <= 12'h42b;
        src18 <= 12'h318;
        src19 <= 12'hab1;
        src20 <= 12'h81c;
        src21 <= 12'hfcf;
        src22 <= 12'h10;
        src23 <= 12'h1c0;
        src24 <= 12'h1e2;
        src25 <= 12'h6f8;
        src26 <= 12'h2e;
        src27 <= 12'h74b;
        src28 <= 12'h219;
        src29 <= 12'hbb7;
        src30 <= 12'h76a;
        src31 <= 12'h6d1;
        src32 <= 12'h5b1;
        src33 <= 12'h95;
        src34 <= 12'hd14;
        src35 <= 12'hcdf;
        src36 <= 12'h601;
        src37 <= 12'h7d0;
        src38 <= 12'h9a5;
        src39 <= 12'h4b;
        src40 <= 12'hd52;
        src41 <= 12'hdc4;
        src42 <= 12'hb75;
        src43 <= 12'h8de;
        src44 <= 12'h5a0;
        src45 <= 12'h34d;
        src46 <= 12'h3ff;
        src47 <= 12'ha5e;
        src48 <= 12'h59c;
        src49 <= 12'h8fa;
        src50 <= 12'haa9;
        src51 <= 12'h472;
        src52 <= 12'hcea;
        src53 <= 12'h30e;
        src54 <= 12'hd63;
        src55 <= 12'h88d;
        src56 <= 12'hb78;
        src57 <= 12'h636;
        src58 <= 12'h7ff;
        src59 <= 12'hf42;
        src60 <= 12'h939;
        src61 <= 12'hf4;
        src62 <= 12'h43f;
        src63 <= 12'he22;
        src64 <= 12'h6ad;
        src65 <= 12'hbd5;
        src66 <= 12'h43;
        src67 <= 12'hfc0;
        src68 <= 12'hab3;
        src69 <= 12'h7a0;
        src70 <= 12'hf68;
        src71 <= 12'h615;
        src72 <= 12'hce;
        src73 <= 12'hb21;
        src74 <= 12'h204;
        src75 <= 12'h6c2;
        src76 <= 12'hb20;
        src77 <= 12'h3ae;
        src78 <= 12'h43c;
        src79 <= 12'hb4e;
        src80 <= 12'h23e;
        src81 <= 12'he69;
        src82 <= 12'hd98;
        src83 <= 12'he09;
        src84 <= 12'h7cd;
        src85 <= 12'h5e0;
        src86 <= 12'h467;
        src87 <= 12'hc92;
        src88 <= 12'hd4b;
        src89 <= 12'hc67;
        src90 <= 12'h7cb;
        src91 <= 12'h97c;
        src92 <= 12'ha49;
        src93 <= 12'h94c;
        src94 <= 12'h884;
        src95 <= 12'h18d;
        src96 <= 12'h1be;
        src97 <= 12'h72f;
        src98 <= 12'h1;
        src99 <= 12'h25b;
        src100 <= 12'hffc;
        src101 <= 12'h560;
        src102 <= 12'he23;
        src103 <= 12'hf0;
        src104 <= 12'h86a;
        src105 <= 12'hd04;
        src106 <= 12'h4e;
        src107 <= 12'h235;
        src108 <= 12'h401;
        src109 <= 12'hce5;
        src110 <= 12'h348;
        src111 <= 12'h761;
        src112 <= 12'h189;
        src113 <= 12'h93a;
        src114 <= 12'h8ae;
        src115 <= 12'ha34;
        src116 <= 12'h248;
        src117 <= 12'hb73;
        src118 <= 12'hb96;
        src119 <= 12'h6d7;
        src120 <= 12'h95e;
        src121 <= 12'he42;
        src122 <= 12'h59d;
        src123 <= 12'h6af;
        src124 <= 12'h766;
        src125 <= 12'h57a;
        src126 <= 12'h5c1;
        src127 <= 12'h478;
        exp <= 19'h3d5f5;
        #1
        src0 <= 12'haa;
        src1 <= 12'he26;
        src2 <= 12'h887;
        src3 <= 12'hc55;
        src4 <= 12'h143;
        src5 <= 12'h70e;
        src6 <= 12'h8d;
        src7 <= 12'h587;
        src8 <= 12'hbfc;
        src9 <= 12'h805;
        src10 <= 12'hc23;
        src11 <= 12'hdf6;
        src12 <= 12'hd15;
        src13 <= 12'h7f;
        src14 <= 12'h9e7;
        src15 <= 12'h73d;
        src16 <= 12'hb9b;
        src17 <= 12'hb4c;
        src18 <= 12'he9d;
        src19 <= 12'h347;
        src20 <= 12'hce6;
        src21 <= 12'h27;
        src22 <= 12'h594;
        src23 <= 12'ha05;
        src24 <= 12'h8c9;
        src25 <= 12'hc81;
        src26 <= 12'he91;
        src27 <= 12'ha6f;
        src28 <= 12'hd7c;
        src29 <= 12'h72;
        src30 <= 12'h838;
        src31 <= 12'h2d8;
        src32 <= 12'h4f5;
        src33 <= 12'h31c;
        src34 <= 12'h3bc;
        src35 <= 12'h5a3;
        src36 <= 12'h772;
        src37 <= 12'h3b0;
        src38 <= 12'h8ef;
        src39 <= 12'h7a4;
        src40 <= 12'h23d;
        src41 <= 12'h17a;
        src42 <= 12'hb9c;
        src43 <= 12'h640;
        src44 <= 12'h3b2;
        src45 <= 12'h3c6;
        src46 <= 12'he2c;
        src47 <= 12'hc82;
        src48 <= 12'h7b2;
        src49 <= 12'h88f;
        src50 <= 12'h7c4;
        src51 <= 12'h3f8;
        src52 <= 12'h2ff;
        src53 <= 12'h6b4;
        src54 <= 12'h581;
        src55 <= 12'h618;
        src56 <= 12'hb2e;
        src57 <= 12'h68;
        src58 <= 12'h98b;
        src59 <= 12'h28d;
        src60 <= 12'h5da;
        src61 <= 12'h975;
        src62 <= 12'hcd2;
        src63 <= 12'h48f;
        src64 <= 12'ha9b;
        src65 <= 12'hef;
        src66 <= 12'hfb0;
        src67 <= 12'h782;
        src68 <= 12'he68;
        src69 <= 12'haa2;
        src70 <= 12'h36f;
        src71 <= 12'h6c9;
        src72 <= 12'h841;
        src73 <= 12'h1fc;
        src74 <= 12'h765;
        src75 <= 12'hd47;
        src76 <= 12'hd0a;
        src77 <= 12'ha45;
        src78 <= 12'h5aa;
        src79 <= 12'h749;
        src80 <= 12'h24c;
        src81 <= 12'h345;
        src82 <= 12'h9be;
        src83 <= 12'haf8;
        src84 <= 12'hc0c;
        src85 <= 12'h4ce;
        src86 <= 12'h5e8;
        src87 <= 12'hde9;
        src88 <= 12'hf3d;
        src89 <= 12'had1;
        src90 <= 12'h7a2;
        src91 <= 12'hc54;
        src92 <= 12'h6e7;
        src93 <= 12'he25;
        src94 <= 12'hfcc;
        src95 <= 12'hc65;
        src96 <= 12'h492;
        src97 <= 12'heb1;
        src98 <= 12'hc8e;
        src99 <= 12'hc99;
        src100 <= 12'hb23;
        src101 <= 12'h5e4;
        src102 <= 12'hc;
        src103 <= 12'hf79;
        src104 <= 12'h947;
        src105 <= 12'hce5;
        src106 <= 12'heb0;
        src107 <= 12'h32e;
        src108 <= 12'hbb2;
        src109 <= 12'h78b;
        src110 <= 12'hd0f;
        src111 <= 12'hbea;
        src112 <= 12'h4da;
        src113 <= 12'ha98;
        src114 <= 12'h64d;
        src115 <= 12'h610;
        src116 <= 12'h1;
        src117 <= 12'h1b;
        src118 <= 12'hae3;
        src119 <= 12'hf59;
        src120 <= 12'h908;
        src121 <= 12'hb4c;
        src122 <= 12'he3d;
        src123 <= 12'hde6;
        src124 <= 12'he02;
        src125 <= 12'h49;
        src126 <= 12'hcde;
        src127 <= 12'h5f8;
        exp <= 19'h42a72;
        #1
        src0 <= 12'hf0f;
        src1 <= 12'h758;
        src2 <= 12'hc1a;
        src3 <= 12'he83;
        src4 <= 12'h15c;
        src5 <= 12'h860;
        src6 <= 12'h3bf;
        src7 <= 12'h489;
        src8 <= 12'h8e7;
        src9 <= 12'h39;
        src10 <= 12'h7f4;
        src11 <= 12'h2b9;
        src12 <= 12'h7b2;
        src13 <= 12'ha90;
        src14 <= 12'hdd3;
        src15 <= 12'h73a;
        src16 <= 12'hacc;
        src17 <= 12'h898;
        src18 <= 12'h26;
        src19 <= 12'hfe9;
        src20 <= 12'h5ee;
        src21 <= 12'hbd2;
        src22 <= 12'he7;
        src23 <= 12'hb7c;
        src24 <= 12'hb56;
        src25 <= 12'h71f;
        src26 <= 12'he68;
        src27 <= 12'h8a5;
        src28 <= 12'haaf;
        src29 <= 12'h632;
        src30 <= 12'h5e7;
        src31 <= 12'h117;
        src32 <= 12'h998;
        src33 <= 12'h8b;
        src34 <= 12'hdfa;
        src35 <= 12'h627;
        src36 <= 12'h8f6;
        src37 <= 12'h398;
        src38 <= 12'h50f;
        src39 <= 12'hbed;
        src40 <= 12'h682;
        src41 <= 12'h549;
        src42 <= 12'h2de;
        src43 <= 12'h8e;
        src44 <= 12'hb12;
        src45 <= 12'h4a8;
        src46 <= 12'hf4b;
        src47 <= 12'h75d;
        src48 <= 12'h27d;
        src49 <= 12'h954;
        src50 <= 12'h8a;
        src51 <= 12'hef8;
        src52 <= 12'h9bf;
        src53 <= 12'ha59;
        src54 <= 12'hd14;
        src55 <= 12'hf99;
        src56 <= 12'h6c3;
        src57 <= 12'hb3f;
        src58 <= 12'hfd3;
        src59 <= 12'hfdc;
        src60 <= 12'h4db;
        src61 <= 12'h5c2;
        src62 <= 12'hf83;
        src63 <= 12'ha3e;
        src64 <= 12'h148;
        src65 <= 12'h92f;
        src66 <= 12'h624;
        src67 <= 12'h406;
        src68 <= 12'h4ae;
        src69 <= 12'hb5b;
        src70 <= 12'h5da;
        src71 <= 12'hc68;
        src72 <= 12'h46d;
        src73 <= 12'h3a7;
        src74 <= 12'h95;
        src75 <= 12'h6b5;
        src76 <= 12'h61c;
        src77 <= 12'h5c6;
        src78 <= 12'h23b;
        src79 <= 12'ha45;
        src80 <= 12'h479;
        src81 <= 12'he3;
        src82 <= 12'hd93;
        src83 <= 12'h300;
        src84 <= 12'hf75;
        src85 <= 12'h4f3;
        src86 <= 12'hd7b;
        src87 <= 12'hcfc;
        src88 <= 12'h824;
        src89 <= 12'hebe;
        src90 <= 12'hd24;
        src91 <= 12'hd6d;
        src92 <= 12'h36a;
        src93 <= 12'h4a5;
        src94 <= 12'h959;
        src95 <= 12'h480;
        src96 <= 12'he66;
        src97 <= 12'h454;
        src98 <= 12'h8de;
        src99 <= 12'ha1e;
        src100 <= 12'h780;
        src101 <= 12'h64;
        src102 <= 12'he5f;
        src103 <= 12'hedf;
        src104 <= 12'h671;
        src105 <= 12'h24;
        src106 <= 12'h84c;
        src107 <= 12'hd92;
        src108 <= 12'hc13;
        src109 <= 12'h9ae;
        src110 <= 12'h7b2;
        src111 <= 12'hcc3;
        src112 <= 12'he73;
        src113 <= 12'h60d;
        src114 <= 12'h21a;
        src115 <= 12'h6b7;
        src116 <= 12'h9b8;
        src117 <= 12'h38f;
        src118 <= 12'he92;
        src119 <= 12'h3a0;
        src120 <= 12'hd2c;
        src121 <= 12'hc49;
        src122 <= 12'h78b;
        src123 <= 12'hc8f;
        src124 <= 12'h77;
        src125 <= 12'hfe5;
        src126 <= 12'h21d;
        src127 <= 12'h96e;
        exp <= 19'h4173f;
        #1
        src0 <= 12'h1da;
        src1 <= 12'hf09;
        src2 <= 12'h7f9;
        src3 <= 12'h393;
        src4 <= 12'h441;
        src5 <= 12'hf06;
        src6 <= 12'h18d;
        src7 <= 12'h1ee;
        src8 <= 12'haa6;
        src9 <= 12'he74;
        src10 <= 12'habe;
        src11 <= 12'h30e;
        src12 <= 12'he44;
        src13 <= 12'hf9a;
        src14 <= 12'hb2e;
        src15 <= 12'hd46;
        src16 <= 12'h5cf;
        src17 <= 12'h6f2;
        src18 <= 12'h752;
        src19 <= 12'h85a;
        src20 <= 12'hc9c;
        src21 <= 12'h645;
        src22 <= 12'he76;
        src23 <= 12'h81d;
        src24 <= 12'hfdd;
        src25 <= 12'h15;
        src26 <= 12'ha53;
        src27 <= 12'hb5a;
        src28 <= 12'ha81;
        src29 <= 12'h9d7;
        src30 <= 12'ha31;
        src31 <= 12'h976;
        src32 <= 12'hf8;
        src33 <= 12'h8e3;
        src34 <= 12'hf32;
        src35 <= 12'h1b1;
        src36 <= 12'h5e4;
        src37 <= 12'hef2;
        src38 <= 12'h3e6;
        src39 <= 12'h814;
        src40 <= 12'hec8;
        src41 <= 12'h111;
        src42 <= 12'hdc8;
        src43 <= 12'h9a7;
        src44 <= 12'h5d;
        src45 <= 12'hecc;
        src46 <= 12'h80c;
        src47 <= 12'h901;
        src48 <= 12'ha5b;
        src49 <= 12'hcf8;
        src50 <= 12'h43c;
        src51 <= 12'h348;
        src52 <= 12'hb00;
        src53 <= 12'h3cf;
        src54 <= 12'h263;
        src55 <= 12'h53f;
        src56 <= 12'h6eb;
        src57 <= 12'hc85;
        src58 <= 12'h8b5;
        src59 <= 12'h3e7;
        src60 <= 12'h5de;
        src61 <= 12'h1f3;
        src62 <= 12'ha9e;
        src63 <= 12'hbe6;
        src64 <= 12'hecd;
        src65 <= 12'hc87;
        src66 <= 12'hbb8;
        src67 <= 12'h226;
        src68 <= 12'h889;
        src69 <= 12'hca7;
        src70 <= 12'hc80;
        src71 <= 12'h89b;
        src72 <= 12'hc5c;
        src73 <= 12'hcfc;
        src74 <= 12'hfca;
        src75 <= 12'h808;
        src76 <= 12'ha0;
        src77 <= 12'h134;
        src78 <= 12'h99d;
        src79 <= 12'hb70;
        src80 <= 12'h7ff;
        src81 <= 12'h4bb;
        src82 <= 12'h988;
        src83 <= 12'hb87;
        src84 <= 12'hc78;
        src85 <= 12'h9ed;
        src86 <= 12'hb1d;
        src87 <= 12'h4a1;
        src88 <= 12'h8ee;
        src89 <= 12'hc25;
        src90 <= 12'h2f4;
        src91 <= 12'h17c;
        src92 <= 12'h14a;
        src93 <= 12'hdc2;
        src94 <= 12'hdbc;
        src95 <= 12'h293;
        src96 <= 12'h8d5;
        src97 <= 12'h34f;
        src98 <= 12'h736;
        src99 <= 12'h50f;
        src100 <= 12'h9a8;
        src101 <= 12'h9e1;
        src102 <= 12'hd8;
        src103 <= 12'hfff;
        src104 <= 12'h1c1;
        src105 <= 12'h663;
        src106 <= 12'h4e7;
        src107 <= 12'hb76;
        src108 <= 12'hffc;
        src109 <= 12'hdc;
        src110 <= 12'h88c;
        src111 <= 12'h23b;
        src112 <= 12'h84d;
        src113 <= 12'h398;
        src114 <= 12'hf7c;
        src115 <= 12'h49d;
        src116 <= 12'hecf;
        src117 <= 12'hb98;
        src118 <= 12'h741;
        src119 <= 12'hc7c;
        src120 <= 12'he58;
        src121 <= 12'h99f;
        src122 <= 12'hfd0;
        src123 <= 12'h752;
        src124 <= 12'h1dc;
        src125 <= 12'h2ff;
        src126 <= 12'h26d;
        src127 <= 12'hb40;
        exp <= 19'h4379b;
        #1
        src0 <= 12'h2db;
        src1 <= 12'h57a;
        src2 <= 12'h95c;
        src3 <= 12'hb53;
        src4 <= 12'hb12;
        src5 <= 12'hb99;
        src6 <= 12'h4a;
        src7 <= 12'hfa;
        src8 <= 12'h850;
        src9 <= 12'h127;
        src10 <= 12'h314;
        src11 <= 12'h81c;
        src12 <= 12'h7e9;
        src13 <= 12'h3de;
        src14 <= 12'h1c4;
        src15 <= 12'h154;
        src16 <= 12'haa4;
        src17 <= 12'hc9d;
        src18 <= 12'h321;
        src19 <= 12'h311;
        src20 <= 12'h264;
        src21 <= 12'ha63;
        src22 <= 12'h3d3;
        src23 <= 12'h96e;
        src24 <= 12'hf97;
        src25 <= 12'h98;
        src26 <= 12'hfea;
        src27 <= 12'hb12;
        src28 <= 12'h1d4;
        src29 <= 12'h2fc;
        src30 <= 12'h73b;
        src31 <= 12'ha2c;
        src32 <= 12'hb7d;
        src33 <= 12'hd19;
        src34 <= 12'he65;
        src35 <= 12'he1;
        src36 <= 12'h14;
        src37 <= 12'hc63;
        src38 <= 12'h7bd;
        src39 <= 12'h6e;
        src40 <= 12'hfe9;
        src41 <= 12'h8b7;
        src42 <= 12'h7da;
        src43 <= 12'h9c5;
        src44 <= 12'h84;
        src45 <= 12'h5eb;
        src46 <= 12'h42e;
        src47 <= 12'ha7b;
        src48 <= 12'h6ba;
        src49 <= 12'h2ce;
        src50 <= 12'h6a;
        src51 <= 12'haa9;
        src52 <= 12'h226;
        src53 <= 12'h314;
        src54 <= 12'h81c;
        src55 <= 12'h356;
        src56 <= 12'ha30;
        src57 <= 12'hc51;
        src58 <= 12'h682;
        src59 <= 12'h738;
        src60 <= 12'hf92;
        src61 <= 12'h12a;
        src62 <= 12'h396;
        src63 <= 12'hdd1;
        src64 <= 12'h58e;
        src65 <= 12'he8b;
        src66 <= 12'hbac;
        src67 <= 12'hac8;
        src68 <= 12'head;
        src69 <= 12'h46;
        src70 <= 12'h635;
        src71 <= 12'hd7a;
        src72 <= 12'hc43;
        src73 <= 12'h1de;
        src74 <= 12'hd8c;
        src75 <= 12'h7c;
        src76 <= 12'hcea;
        src77 <= 12'haee;
        src78 <= 12'hbd1;
        src79 <= 12'hb3d;
        src80 <= 12'h3a;
        src81 <= 12'h5c6;
        src82 <= 12'h4d3;
        src83 <= 12'hb6;
        src84 <= 12'h6c2;
        src85 <= 12'hd1d;
        src86 <= 12'h365;
        src87 <= 12'h690;
        src88 <= 12'hbbd;
        src89 <= 12'h1f6;
        src90 <= 12'h528;
        src91 <= 12'hc97;
        src92 <= 12'h7ba;
        src93 <= 12'h34b;
        src94 <= 12'h41a;
        src95 <= 12'hf8a;
        src96 <= 12'h8aa;
        src97 <= 12'hc79;
        src98 <= 12'h5d0;
        src99 <= 12'hbf2;
        src100 <= 12'he4d;
        src101 <= 12'h4cf;
        src102 <= 12'h854;
        src103 <= 12'h36;
        src104 <= 12'h9e0;
        src105 <= 12'h75d;
        src106 <= 12'h461;
        src107 <= 12'hb06;
        src108 <= 12'h4fa;
        src109 <= 12'h85c;
        src110 <= 12'h6f1;
        src111 <= 12'heb8;
        src112 <= 12'ha96;
        src113 <= 12'h966;
        src114 <= 12'h445;
        src115 <= 12'h212;
        src116 <= 12'h2b6;
        src117 <= 12'h167;
        src118 <= 12'hbe5;
        src119 <= 12'h6e6;
        src120 <= 12'h18d;
        src121 <= 12'h9ce;
        src122 <= 12'hfe8;
        src123 <= 12'h25a;
        src124 <= 12'h37c;
        src125 <= 12'hd1e;
        src126 <= 12'h58e;
        src127 <= 12'h4c5;
        exp <= 19'h3a879;
        #1
        src0 <= 12'ha3c;
        src1 <= 12'hd51;
        src2 <= 12'hb37;
        src3 <= 12'h600;
        src4 <= 12'h242;
        src5 <= 12'hf7c;
        src6 <= 12'h40;
        src7 <= 12'h4a2;
        src8 <= 12'h91b;
        src9 <= 12'h74c;
        src10 <= 12'h8d1;
        src11 <= 12'h754;
        src12 <= 12'h798;
        src13 <= 12'hf98;
        src14 <= 12'h78d;
        src15 <= 12'h6a2;
        src16 <= 12'hda3;
        src17 <= 12'h7d0;
        src18 <= 12'h62f;
        src19 <= 12'h9e7;
        src20 <= 12'h5c;
        src21 <= 12'hdf2;
        src22 <= 12'hc7b;
        src23 <= 12'ha92;
        src24 <= 12'h5e5;
        src25 <= 12'ha44;
        src26 <= 12'h585;
        src27 <= 12'h353;
        src28 <= 12'h288;
        src29 <= 12'h59d;
        src30 <= 12'h14b;
        src31 <= 12'ha81;
        src32 <= 12'ha48;
        src33 <= 12'h658;
        src34 <= 12'h846;
        src35 <= 12'h5d7;
        src36 <= 12'h201;
        src37 <= 12'h54b;
        src38 <= 12'h33e;
        src39 <= 12'h63f;
        src40 <= 12'hb5a;
        src41 <= 12'h971;
        src42 <= 12'h69e;
        src43 <= 12'hd2c;
        src44 <= 12'h1d;
        src45 <= 12'h4c6;
        src46 <= 12'hfa3;
        src47 <= 12'h216;
        src48 <= 12'h1f9;
        src49 <= 12'h201;
        src50 <= 12'h40d;
        src51 <= 12'h9cd;
        src52 <= 12'h47a;
        src53 <= 12'hdcc;
        src54 <= 12'hb19;
        src55 <= 12'h802;
        src56 <= 12'h37c;
        src57 <= 12'h3a0;
        src58 <= 12'hab1;
        src59 <= 12'h696;
        src60 <= 12'h776;
        src61 <= 12'h3f6;
        src62 <= 12'h31c;
        src63 <= 12'hb56;
        src64 <= 12'h206;
        src65 <= 12'h15;
        src66 <= 12'ha72;
        src67 <= 12'h100;
        src68 <= 12'hb85;
        src69 <= 12'h6f1;
        src70 <= 12'h500;
        src71 <= 12'ha46;
        src72 <= 12'hae3;
        src73 <= 12'h2af;
        src74 <= 12'haa7;
        src75 <= 12'h7b5;
        src76 <= 12'hf6b;
        src77 <= 12'ha25;
        src78 <= 12'h733;
        src79 <= 12'h5f3;
        src80 <= 12'hd30;
        src81 <= 12'h2a5;
        src82 <= 12'hfe4;
        src83 <= 12'h16b;
        src84 <= 12'h8d;
        src85 <= 12'h228;
        src86 <= 12'h895;
        src87 <= 12'h234;
        src88 <= 12'h5eb;
        src89 <= 12'h967;
        src90 <= 12'hd49;
        src91 <= 12'h443;
        src92 <= 12'h622;
        src93 <= 12'h8bb;
        src94 <= 12'h3b7;
        src95 <= 12'h93d;
        src96 <= 12'hb2a;
        src97 <= 12'h159;
        src98 <= 12'hd2a;
        src99 <= 12'h646;
        src100 <= 12'h8f1;
        src101 <= 12'hf29;
        src102 <= 12'h4a1;
        src103 <= 12'h52e;
        src104 <= 12'he2b;
        src105 <= 12'h5c0;
        src106 <= 12'h98f;
        src107 <= 12'hb66;
        src108 <= 12'he2c;
        src109 <= 12'h2b;
        src110 <= 12'h780;
        src111 <= 12'h107;
        src112 <= 12'h406;
        src113 <= 12'hb0e;
        src114 <= 12'heb1;
        src115 <= 12'h51e;
        src116 <= 12'h8a1;
        src117 <= 12'h757;
        src118 <= 12'h1c3;
        src119 <= 12'hd84;
        src120 <= 12'h60b;
        src121 <= 12'h6cd;
        src122 <= 12'h528;
        src123 <= 12'h61b;
        src124 <= 12'hf5a;
        src125 <= 12'h628;
        src126 <= 12'h92;
        src127 <= 12'hb37;
        exp <= 19'h3b3b2;
        #1
        src0 <= 12'hdb0;
        src1 <= 12'ha44;
        src2 <= 12'h92b;
        src3 <= 12'h8d4;
        src4 <= 12'h997;
        src5 <= 12'h60f;
        src6 <= 12'h7ac;
        src7 <= 12'h6a0;
        src8 <= 12'h770;
        src9 <= 12'ha9f;
        src10 <= 12'h552;
        src11 <= 12'h5f1;
        src12 <= 12'hc01;
        src13 <= 12'h1a6;
        src14 <= 12'h7e;
        src15 <= 12'h90d;
        src16 <= 12'h2c2;
        src17 <= 12'h6ab;
        src18 <= 12'hbdc;
        src19 <= 12'h28d;
        src20 <= 12'h98b;
        src21 <= 12'hed1;
        src22 <= 12'hdfc;
        src23 <= 12'hb88;
        src24 <= 12'h1be;
        src25 <= 12'ha24;
        src26 <= 12'he38;
        src27 <= 12'hd36;
        src28 <= 12'h9ad;
        src29 <= 12'hb13;
        src30 <= 12'h421;
        src31 <= 12'hf28;
        src32 <= 12'hd31;
        src33 <= 12'h1fc;
        src34 <= 12'h7eb;
        src35 <= 12'he27;
        src36 <= 12'h858;
        src37 <= 12'h1c2;
        src38 <= 12'heea;
        src39 <= 12'h3d7;
        src40 <= 12'h49f;
        src41 <= 12'ha0d;
        src42 <= 12'hf5c;
        src43 <= 12'h4b3;
        src44 <= 12'haf9;
        src45 <= 12'hdbe;
        src46 <= 12'hda1;
        src47 <= 12'h3cd;
        src48 <= 12'hdf4;
        src49 <= 12'he6e;
        src50 <= 12'hdc6;
        src51 <= 12'h9f;
        src52 <= 12'h788;
        src53 <= 12'hb22;
        src54 <= 12'h9c6;
        src55 <= 12'hb1e;
        src56 <= 12'h264;
        src57 <= 12'h501;
        src58 <= 12'hd6c;
        src59 <= 12'h7aa;
        src60 <= 12'hbd;
        src61 <= 12'ha1;
        src62 <= 12'hf38;
        src63 <= 12'h6c3;
        src64 <= 12'hf02;
        src65 <= 12'hf08;
        src66 <= 12'hd3a;
        src67 <= 12'h53c;
        src68 <= 12'hdfb;
        src69 <= 12'hc9e;
        src70 <= 12'h8f3;
        src71 <= 12'h79a;
        src72 <= 12'ha74;
        src73 <= 12'h3a4;
        src74 <= 12'h62d;
        src75 <= 12'h353;
        src76 <= 12'heec;
        src77 <= 12'ha51;
        src78 <= 12'h21b;
        src79 <= 12'h9c1;
        src80 <= 12'hb67;
        src81 <= 12'hfd4;
        src82 <= 12'h4b6;
        src83 <= 12'h508;
        src84 <= 12'h88d;
        src85 <= 12'h71d;
        src86 <= 12'hecb;
        src87 <= 12'h95e;
        src88 <= 12'h932;
        src89 <= 12'h282;
        src90 <= 12'h38e;
        src91 <= 12'h314;
        src92 <= 12'hb62;
        src93 <= 12'h720;
        src94 <= 12'h5a7;
        src95 <= 12'hcfd;
        src96 <= 12'hbd1;
        src97 <= 12'h5a6;
        src98 <= 12'h85d;
        src99 <= 12'h567;
        src100 <= 12'hd13;
        src101 <= 12'h6e;
        src102 <= 12'h824;
        src103 <= 12'h4e4;
        src104 <= 12'h286;
        src105 <= 12'h500;
        src106 <= 12'he46;
        src107 <= 12'hdb7;
        src108 <= 12'hf42;
        src109 <= 12'h42;
        src110 <= 12'hebb;
        src111 <= 12'h835;
        src112 <= 12'h654;
        src113 <= 12'h73;
        src114 <= 12'hc69;
        src115 <= 12'hff3;
        src116 <= 12'h8da;
        src117 <= 12'h17f;
        src118 <= 12'hc27;
        src119 <= 12'hd96;
        src120 <= 12'h1cb;
        src121 <= 12'hdf6;
        src122 <= 12'h286;
        src123 <= 12'hfbf;
        src124 <= 12'h555;
        src125 <= 12'hea5;
        src126 <= 12'h784;
        src127 <= 12'hc08;
        exp <= 19'h45bba;
        #1
        src0 <= 12'h349;
        src1 <= 12'hffa;
        src2 <= 12'h5ce;
        src3 <= 12'h4b2;
        src4 <= 12'hd59;
        src5 <= 12'h497;
        src6 <= 12'hfa0;
        src7 <= 12'heec;
        src8 <= 12'h482;
        src9 <= 12'hc19;
        src10 <= 12'h5e2;
        src11 <= 12'he25;
        src12 <= 12'h92f;
        src13 <= 12'hf0;
        src14 <= 12'h817;
        src15 <= 12'h751;
        src16 <= 12'h945;
        src17 <= 12'h24c;
        src18 <= 12'h62f;
        src19 <= 12'hb74;
        src20 <= 12'h683;
        src21 <= 12'hf10;
        src22 <= 12'hbf;
        src23 <= 12'h3bf;
        src24 <= 12'hf07;
        src25 <= 12'hecf;
        src26 <= 12'h7c2;
        src27 <= 12'h316;
        src28 <= 12'heb0;
        src29 <= 12'h5e0;
        src30 <= 12'ha9c;
        src31 <= 12'he95;
        src32 <= 12'hb6d;
        src33 <= 12'hf79;
        src34 <= 12'hf4f;
        src35 <= 12'h811;
        src36 <= 12'h36d;
        src37 <= 12'h78;
        src38 <= 12'h3f4;
        src39 <= 12'ha29;
        src40 <= 12'h2b2;
        src41 <= 12'h3fd;
        src42 <= 12'hf50;
        src43 <= 12'h303;
        src44 <= 12'h278;
        src45 <= 12'h96f;
        src46 <= 12'h22d;
        src47 <= 12'h5b6;
        src48 <= 12'h85d;
        src49 <= 12'ha15;
        src50 <= 12'h870;
        src51 <= 12'h9a;
        src52 <= 12'h26a;
        src53 <= 12'hc79;
        src54 <= 12'h617;
        src55 <= 12'h51d;
        src56 <= 12'h826;
        src57 <= 12'h890;
        src58 <= 12'hcc1;
        src59 <= 12'h44f;
        src60 <= 12'hb9;
        src61 <= 12'h7de;
        src62 <= 12'hcb2;
        src63 <= 12'hb14;
        src64 <= 12'h5c7;
        src65 <= 12'h6ef;
        src66 <= 12'hb4d;
        src67 <= 12'hb7;
        src68 <= 12'h1d0;
        src69 <= 12'h7bf;
        src70 <= 12'h1df;
        src71 <= 12'h83f;
        src72 <= 12'h2;
        src73 <= 12'h81a;
        src74 <= 12'he82;
        src75 <= 12'h878;
        src76 <= 12'h3c0;
        src77 <= 12'h191;
        src78 <= 12'h4cf;
        src79 <= 12'h25e;
        src80 <= 12'h120;
        src81 <= 12'h6e5;
        src82 <= 12'h74d;
        src83 <= 12'h683;
        src84 <= 12'h4da;
        src85 <= 12'h4c;
        src86 <= 12'h9d5;
        src87 <= 12'h867;
        src88 <= 12'h94a;
        src89 <= 12'ha08;
        src90 <= 12'h77e;
        src91 <= 12'hf4b;
        src92 <= 12'he15;
        src93 <= 12'h3e4;
        src94 <= 12'h43b;
        src95 <= 12'h89f;
        src96 <= 12'he64;
        src97 <= 12'hf78;
        src98 <= 12'h3e1;
        src99 <= 12'h2fc;
        src100 <= 12'hbda;
        src101 <= 12'heb8;
        src102 <= 12'hdd;
        src103 <= 12'h215;
        src104 <= 12'hb09;
        src105 <= 12'h1a5;
        src106 <= 12'h165;
        src107 <= 12'hccb;
        src108 <= 12'hc82;
        src109 <= 12'hf1e;
        src110 <= 12'h2d2;
        src111 <= 12'hdd4;
        src112 <= 12'h9ed;
        src113 <= 12'he0c;
        src114 <= 12'h31e;
        src115 <= 12'ha3e;
        src116 <= 12'h481;
        src117 <= 12'h816;
        src118 <= 12'h7d9;
        src119 <= 12'h80b;
        src120 <= 12'h943;
        src121 <= 12'h7bf;
        src122 <= 12'h6d1;
        src123 <= 12'h78a;
        src124 <= 12'h30c;
        src125 <= 12'h904;
        src126 <= 12'h958;
        src127 <= 12'h317;
        exp <= 19'h3d413;
        #1
        src0 <= 12'h600;
        src1 <= 12'h135;
        src2 <= 12'h779;
        src3 <= 12'h6c1;
        src4 <= 12'h78d;
        src5 <= 12'h1f7;
        src6 <= 12'hc25;
        src7 <= 12'h630;
        src8 <= 12'hf;
        src9 <= 12'h9f7;
        src10 <= 12'h51c;
        src11 <= 12'hc9f;
        src12 <= 12'h8a0;
        src13 <= 12'h798;
        src14 <= 12'hca1;
        src15 <= 12'h77b;
        src16 <= 12'h706;
        src17 <= 12'hd78;
        src18 <= 12'hc7b;
        src19 <= 12'h455;
        src20 <= 12'h36c;
        src21 <= 12'hc33;
        src22 <= 12'haf9;
        src23 <= 12'hf60;
        src24 <= 12'h2fa;
        src25 <= 12'h711;
        src26 <= 12'h400;
        src27 <= 12'hef7;
        src28 <= 12'hf2e;
        src29 <= 12'hcc8;
        src30 <= 12'h811;
        src31 <= 12'h524;
        src32 <= 12'hd2c;
        src33 <= 12'h68e;
        src34 <= 12'haef;
        src35 <= 12'hd03;
        src36 <= 12'h876;
        src37 <= 12'h9ad;
        src38 <= 12'h721;
        src39 <= 12'h334;
        src40 <= 12'h2ed;
        src41 <= 12'he89;
        src42 <= 12'hc31;
        src43 <= 12'hff3;
        src44 <= 12'hcbf;
        src45 <= 12'hd19;
        src46 <= 12'hf88;
        src47 <= 12'hfe3;
        src48 <= 12'h283;
        src49 <= 12'h526;
        src50 <= 12'hf57;
        src51 <= 12'hdc1;
        src52 <= 12'h2fd;
        src53 <= 12'hf96;
        src54 <= 12'h5cf;
        src55 <= 12'hca8;
        src56 <= 12'hf64;
        src57 <= 12'h436;
        src58 <= 12'hbab;
        src59 <= 12'ha85;
        src60 <= 12'hc97;
        src61 <= 12'h391;
        src62 <= 12'hbec;
        src63 <= 12'h2ab;
        src64 <= 12'h8c2;
        src65 <= 12'h848;
        src66 <= 12'h32b;
        src67 <= 12'h465;
        src68 <= 12'h282;
        src69 <= 12'he1c;
        src70 <= 12'h283;
        src71 <= 12'h278;
        src72 <= 12'hbdc;
        src73 <= 12'h725;
        src74 <= 12'h75;
        src75 <= 12'hbb6;
        src76 <= 12'h83a;
        src77 <= 12'h21b;
        src78 <= 12'h20;
        src79 <= 12'hd81;
        src80 <= 12'hde5;
        src81 <= 12'h662;
        src82 <= 12'he3e;
        src83 <= 12'h57;
        src84 <= 12'hfc5;
        src85 <= 12'hfba;
        src86 <= 12'h3fd;
        src87 <= 12'h4d1;
        src88 <= 12'hcf9;
        src89 <= 12'h29d;
        src90 <= 12'hb80;
        src91 <= 12'h1dc;
        src92 <= 12'he71;
        src93 <= 12'hf94;
        src94 <= 12'hfad;
        src95 <= 12'head;
        src96 <= 12'h9d0;
        src97 <= 12'hb82;
        src98 <= 12'hbb5;
        src99 <= 12'he31;
        src100 <= 12'hee;
        src101 <= 12'hb19;
        src102 <= 12'hb5b;
        src103 <= 12'ha3c;
        src104 <= 12'h638;
        src105 <= 12'h1c2;
        src106 <= 12'h169;
        src107 <= 12'h6e0;
        src108 <= 12'ha9;
        src109 <= 12'hb91;
        src110 <= 12'he4f;
        src111 <= 12'hbe6;
        src112 <= 12'hfb2;
        src113 <= 12'h63d;
        src114 <= 12'hfb8;
        src115 <= 12'h7f9;
        src116 <= 12'hfb3;
        src117 <= 12'hc70;
        src118 <= 12'h333;
        src119 <= 12'h7a9;
        src120 <= 12'hd49;
        src121 <= 12'h1d3;
        src122 <= 12'hb53;
        src123 <= 12'hb6;
        src124 <= 12'h985;
        src125 <= 12'h141;
        src126 <= 12'hc3d;
        src127 <= 12'h54a;
        exp <= 19'h4658d;
        #1
        src0 <= 12'hc28;
        src1 <= 12'h178;
        src2 <= 12'h877;
        src3 <= 12'hcb8;
        src4 <= 12'hae5;
        src5 <= 12'hf79;
        src6 <= 12'h78a;
        src7 <= 12'hbfa;
        src8 <= 12'h108;
        src9 <= 12'hc0c;
        src10 <= 12'h9f6;
        src11 <= 12'h879;
        src12 <= 12'h6ab;
        src13 <= 12'h4ca;
        src14 <= 12'haf0;
        src15 <= 12'hf13;
        src16 <= 12'h389;
        src17 <= 12'h288;
        src18 <= 12'h6c4;
        src19 <= 12'h66f;
        src20 <= 12'hd00;
        src21 <= 12'h688;
        src22 <= 12'h474;
        src23 <= 12'h52;
        src24 <= 12'hb8b;
        src25 <= 12'h7ef;
        src26 <= 12'hca2;
        src27 <= 12'h636;
        src28 <= 12'h268;
        src29 <= 12'h408;
        src30 <= 12'h1d4;
        src31 <= 12'he65;
        src32 <= 12'had4;
        src33 <= 12'h974;
        src34 <= 12'hd34;
        src35 <= 12'hb04;
        src36 <= 12'h994;
        src37 <= 12'h7ff;
        src38 <= 12'h16f;
        src39 <= 12'hc22;
        src40 <= 12'h4a3;
        src41 <= 12'h612;
        src42 <= 12'hc38;
        src43 <= 12'h2d;
        src44 <= 12'h9a3;
        src45 <= 12'h411;
        src46 <= 12'h213;
        src47 <= 12'hda6;
        src48 <= 12'h194;
        src49 <= 12'h86b;
        src50 <= 12'hc33;
        src51 <= 12'h44a;
        src52 <= 12'hf55;
        src53 <= 12'h59b;
        src54 <= 12'hd1;
        src55 <= 12'hb98;
        src56 <= 12'h17e;
        src57 <= 12'h6b7;
        src58 <= 12'hb2f;
        src59 <= 12'h7b4;
        src60 <= 12'h6f5;
        src61 <= 12'h38d;
        src62 <= 12'hb99;
        src63 <= 12'ha2;
        src64 <= 12'h329;
        src65 <= 12'he;
        src66 <= 12'h37e;
        src67 <= 12'h884;
        src68 <= 12'he9f;
        src69 <= 12'h80f;
        src70 <= 12'h445;
        src71 <= 12'h6a7;
        src72 <= 12'h607;
        src73 <= 12'hcbc;
        src74 <= 12'h31c;
        src75 <= 12'h9d9;
        src76 <= 12'h119;
        src77 <= 12'ha7b;
        src78 <= 12'hca0;
        src79 <= 12'heea;
        src80 <= 12'h8af;
        src81 <= 12'hba3;
        src82 <= 12'hbc5;
        src83 <= 12'h4f5;
        src84 <= 12'hf08;
        src85 <= 12'h730;
        src86 <= 12'h2d5;
        src87 <= 12'h59f;
        src88 <= 12'h4a5;
        src89 <= 12'hdea;
        src90 <= 12'hc3f;
        src91 <= 12'h955;
        src92 <= 12'h6d;
        src93 <= 12'h56f;
        src94 <= 12'h8aa;
        src95 <= 12'hf09;
        src96 <= 12'h821;
        src97 <= 12'h65;
        src98 <= 12'hd2e;
        src99 <= 12'hacc;
        src100 <= 12'hf75;
        src101 <= 12'hee0;
        src102 <= 12'h130;
        src103 <= 12'h343;
        src104 <= 12'hd9;
        src105 <= 12'h896;
        src106 <= 12'hf2f;
        src107 <= 12'hfb3;
        src108 <= 12'h52c;
        src109 <= 12'hbda;
        src110 <= 12'h43d;
        src111 <= 12'h431;
        src112 <= 12'hff7;
        src113 <= 12'ha2f;
        src114 <= 12'h439;
        src115 <= 12'hd5c;
        src116 <= 12'hd6a;
        src117 <= 12'h47a;
        src118 <= 12'h5c4;
        src119 <= 12'h310;
        src120 <= 12'hf69;
        src121 <= 12'h438;
        src122 <= 12'he83;
        src123 <= 12'h42a;
        src124 <= 12'h9c0;
        src125 <= 12'h340;
        src126 <= 12'hd21;
        src127 <= 12'h47f;
        exp <= 19'h3fd8f;
        #1
        src0 <= 12'h605;
        src1 <= 12'h29a;
        src2 <= 12'h5dc;
        src3 <= 12'ha09;
        src4 <= 12'hd9d;
        src5 <= 12'h300;
        src6 <= 12'hb77;
        src7 <= 12'h9e9;
        src8 <= 12'h465;
        src9 <= 12'h916;
        src10 <= 12'h197;
        src11 <= 12'hc03;
        src12 <= 12'h1d3;
        src13 <= 12'h708;
        src14 <= 12'h983;
        src15 <= 12'hc47;
        src16 <= 12'h96b;
        src17 <= 12'hac7;
        src18 <= 12'hc14;
        src19 <= 12'hac3;
        src20 <= 12'h554;
        src21 <= 12'h571;
        src22 <= 12'ha26;
        src23 <= 12'h44;
        src24 <= 12'hbc4;
        src25 <= 12'hf35;
        src26 <= 12'hfe8;
        src27 <= 12'hcec;
        src28 <= 12'h57b;
        src29 <= 12'hfe5;
        src30 <= 12'h9b;
        src31 <= 12'h6d5;
        src32 <= 12'hc0b;
        src33 <= 12'ha9d;
        src34 <= 12'h298;
        src35 <= 12'h844;
        src36 <= 12'h931;
        src37 <= 12'h1f0;
        src38 <= 12'h538;
        src39 <= 12'h3e3;
        src40 <= 12'hdb0;
        src41 <= 12'ha7;
        src42 <= 12'h9f3;
        src43 <= 12'h907;
        src44 <= 12'h98a;
        src45 <= 12'h1f7;
        src46 <= 12'ha04;
        src47 <= 12'hf30;
        src48 <= 12'ha8f;
        src49 <= 12'h717;
        src50 <= 12'h7b6;
        src51 <= 12'h18d;
        src52 <= 12'h377;
        src53 <= 12'h63f;
        src54 <= 12'hea6;
        src55 <= 12'hdcd;
        src56 <= 12'h382;
        src57 <= 12'h742;
        src58 <= 12'h214;
        src59 <= 12'hf90;
        src60 <= 12'hb10;
        src61 <= 12'h186;
        src62 <= 12'h3ee;
        src63 <= 12'h11e;
        src64 <= 12'hb47;
        src65 <= 12'ha47;
        src66 <= 12'h90c;
        src67 <= 12'hdc;
        src68 <= 12'h91b;
        src69 <= 12'h342;
        src70 <= 12'h52;
        src71 <= 12'he0d;
        src72 <= 12'ha27;
        src73 <= 12'ha9b;
        src74 <= 12'h3b9;
        src75 <= 12'h6f6;
        src76 <= 12'h902;
        src77 <= 12'h26f;
        src78 <= 12'h3c7;
        src79 <= 12'h4fe;
        src80 <= 12'h482;
        src81 <= 12'hc2;
        src82 <= 12'hb26;
        src83 <= 12'h8b2;
        src84 <= 12'h4ce;
        src85 <= 12'h30e;
        src86 <= 12'h1ae;
        src87 <= 12'h8ad;
        src88 <= 12'hc18;
        src89 <= 12'hffe;
        src90 <= 12'h33e;
        src91 <= 12'hb2e;
        src92 <= 12'h1f5;
        src93 <= 12'hf83;
        src94 <= 12'h7aa;
        src95 <= 12'hc5;
        src96 <= 12'h945;
        src97 <= 12'hffe;
        src98 <= 12'h380;
        src99 <= 12'hd6a;
        src100 <= 12'h728;
        src101 <= 12'hb01;
        src102 <= 12'h3e5;
        src103 <= 12'he94;
        src104 <= 12'h407;
        src105 <= 12'hc4c;
        src106 <= 12'hcd6;
        src107 <= 12'h18e;
        src108 <= 12'h37c;
        src109 <= 12'h6e3;
        src110 <= 12'hf14;
        src111 <= 12'h832;
        src112 <= 12'h67c;
        src113 <= 12'h15b;
        src114 <= 12'hb03;
        src115 <= 12'h765;
        src116 <= 12'he12;
        src117 <= 12'h88;
        src118 <= 12'h644;
        src119 <= 12'h23a;
        src120 <= 12'h6b4;
        src121 <= 12'he7d;
        src122 <= 12'hd20;
        src123 <= 12'h66e;
        src124 <= 12'h112;
        src125 <= 12'h77c;
        src126 <= 12'h1a0;
        src127 <= 12'h8d2;
        exp <= 19'h3d1c8;
        #1
        src0 <= 12'hf01;
        src1 <= 12'h213;
        src2 <= 12'hf70;
        src3 <= 12'ha93;
        src4 <= 12'hebe;
        src5 <= 12'h715;
        src6 <= 12'h86e;
        src7 <= 12'h26d;
        src8 <= 12'h54e;
        src9 <= 12'h910;
        src10 <= 12'hbe5;
        src11 <= 12'hf49;
        src12 <= 12'h6b4;
        src13 <= 12'hd0f;
        src14 <= 12'h58d;
        src15 <= 12'h933;
        src16 <= 12'hf53;
        src17 <= 12'h4d2;
        src18 <= 12'h62a;
        src19 <= 12'h814;
        src20 <= 12'he23;
        src21 <= 12'h964;
        src22 <= 12'h36b;
        src23 <= 12'h4ff;
        src24 <= 12'hc38;
        src25 <= 12'h1a8;
        src26 <= 12'he80;
        src27 <= 12'hb03;
        src28 <= 12'h1c8;
        src29 <= 12'h1c4;
        src30 <= 12'hedb;
        src31 <= 12'hb2f;
        src32 <= 12'h971;
        src33 <= 12'hbb0;
        src34 <= 12'hd2b;
        src35 <= 12'h903;
        src36 <= 12'hbd4;
        src37 <= 12'hc4e;
        src38 <= 12'hf88;
        src39 <= 12'h7c5;
        src40 <= 12'h85d;
        src41 <= 12'h846;
        src42 <= 12'hf05;
        src43 <= 12'h5fe;
        src44 <= 12'h418;
        src45 <= 12'hbf1;
        src46 <= 12'h45c;
        src47 <= 12'h4a5;
        src48 <= 12'hf73;
        src49 <= 12'h5b0;
        src50 <= 12'ha4e;
        src51 <= 12'h856;
        src52 <= 12'h839;
        src53 <= 12'he3;
        src54 <= 12'h324;
        src55 <= 12'hb38;
        src56 <= 12'hab0;
        src57 <= 12'hb02;
        src58 <= 12'h167;
        src59 <= 12'h8;
        src60 <= 12'hba3;
        src61 <= 12'h2e4;
        src62 <= 12'hdad;
        src63 <= 12'h126;
        src64 <= 12'h7a8;
        src65 <= 12'hc45;
        src66 <= 12'h9e3;
        src67 <= 12'h2b1;
        src68 <= 12'h5af;
        src69 <= 12'h1a5;
        src70 <= 12'h1a0;
        src71 <= 12'h725;
        src72 <= 12'h6ab;
        src73 <= 12'hc2;
        src74 <= 12'h45;
        src75 <= 12'he83;
        src76 <= 12'h34b;
        src77 <= 12'h1cb;
        src78 <= 12'h4e7;
        src79 <= 12'h935;
        src80 <= 12'h570;
        src81 <= 12'hb84;
        src82 <= 12'h1f2;
        src83 <= 12'ha67;
        src84 <= 12'hcd;
        src85 <= 12'h442;
        src86 <= 12'hcd;
        src87 <= 12'hee6;
        src88 <= 12'h258;
        src89 <= 12'h4e2;
        src90 <= 12'h313;
        src91 <= 12'hfb5;
        src92 <= 12'h913;
        src93 <= 12'hd31;
        src94 <= 12'h8c;
        src95 <= 12'h68a;
        src96 <= 12'h625;
        src97 <= 12'h337;
        src98 <= 12'hf9d;
        src99 <= 12'h815;
        src100 <= 12'hecd;
        src101 <= 12'hc53;
        src102 <= 12'hd3b;
        src103 <= 12'h9cf;
        src104 <= 12'h156;
        src105 <= 12'ha5e;
        src106 <= 12'h17f;
        src107 <= 12'hc7c;
        src108 <= 12'h1af;
        src109 <= 12'h68;
        src110 <= 12'hf8e;
        src111 <= 12'hcb4;
        src112 <= 12'h8ed;
        src113 <= 12'he7a;
        src114 <= 12'h7fb;
        src115 <= 12'h431;
        src116 <= 12'h7da;
        src117 <= 12'had5;
        src118 <= 12'h769;
        src119 <= 12'h30d;
        src120 <= 12'h77b;
        src121 <= 12'h20e;
        src122 <= 12'he02;
        src123 <= 12'h96f;
        src124 <= 12'hb81;
        src125 <= 12'h9bd;
        src126 <= 12'h2cb;
        src127 <= 12'hca5;
        exp <= 19'h40155;
        #1
        src0 <= 12'h893;
        src1 <= 12'h5e8;
        src2 <= 12'h839;
        src3 <= 12'h7e3;
        src4 <= 12'h8e4;
        src5 <= 12'h6ee;
        src6 <= 12'h351;
        src7 <= 12'h403;
        src8 <= 12'h4b2;
        src9 <= 12'h864;
        src10 <= 12'h7aa;
        src11 <= 12'hd4;
        src12 <= 12'h9eb;
        src13 <= 12'hf66;
        src14 <= 12'h12f;
        src15 <= 12'he11;
        src16 <= 12'h45e;
        src17 <= 12'h499;
        src18 <= 12'hc36;
        src19 <= 12'hde9;
        src20 <= 12'ha28;
        src21 <= 12'h750;
        src22 <= 12'h491;
        src23 <= 12'heac;
        src24 <= 12'hf9c;
        src25 <= 12'hb84;
        src26 <= 12'h8e7;
        src27 <= 12'he40;
        src28 <= 12'h624;
        src29 <= 12'h65c;
        src30 <= 12'h8b5;
        src31 <= 12'hf43;
        src32 <= 12'h40a;
        src33 <= 12'hd6a;
        src34 <= 12'h91b;
        src35 <= 12'ha17;
        src36 <= 12'h336;
        src37 <= 12'h786;
        src38 <= 12'ha81;
        src39 <= 12'h7bc;
        src40 <= 12'hcca;
        src41 <= 12'he17;
        src42 <= 12'haf4;
        src43 <= 12'ha8b;
        src44 <= 12'h57b;
        src45 <= 12'hf35;
        src46 <= 12'h96;
        src47 <= 12'hfe8;
        src48 <= 12'h73d;
        src49 <= 12'h218;
        src50 <= 12'h2b;
        src51 <= 12'h959;
        src52 <= 12'h844;
        src53 <= 12'he57;
        src54 <= 12'h6a2;
        src55 <= 12'h1b8;
        src56 <= 12'h156;
        src57 <= 12'h810;
        src58 <= 12'hd1e;
        src59 <= 12'h330;
        src60 <= 12'hc8;
        src61 <= 12'h8c0;
        src62 <= 12'h3c9;
        src63 <= 12'h724;
        src64 <= 12'hb9f;
        src65 <= 12'h32b;
        src66 <= 12'h819;
        src67 <= 12'h9b;
        src68 <= 12'h693;
        src69 <= 12'h930;
        src70 <= 12'he3c;
        src71 <= 12'hda6;
        src72 <= 12'h863;
        src73 <= 12'hbb2;
        src74 <= 12'hcec;
        src75 <= 12'h62e;
        src76 <= 12'h769;
        src77 <= 12'h83b;
        src78 <= 12'h59;
        src79 <= 12'h1fb;
        src80 <= 12'h1f3;
        src81 <= 12'h768;
        src82 <= 12'h9dc;
        src83 <= 12'h72;
        src84 <= 12'h5dc;
        src85 <= 12'h557;
        src86 <= 12'h47f;
        src87 <= 12'ha0f;
        src88 <= 12'h24e;
        src89 <= 12'hc60;
        src90 <= 12'h981;
        src91 <= 12'h725;
        src92 <= 12'h3fb;
        src93 <= 12'h262;
        src94 <= 12'h298;
        src95 <= 12'hf3e;
        src96 <= 12'hce3;
        src97 <= 12'h68b;
        src98 <= 12'h25f;
        src99 <= 12'h2b9;
        src100 <= 12'h585;
        src101 <= 12'h698;
        src102 <= 12'h8cc;
        src103 <= 12'he31;
        src104 <= 12'h784;
        src105 <= 12'hf10;
        src106 <= 12'h19a;
        src107 <= 12'hcfd;
        src108 <= 12'h89e;
        src109 <= 12'h1ad;
        src110 <= 12'hca7;
        src111 <= 12'hbde;
        src112 <= 12'hfd6;
        src113 <= 12'h82b;
        src114 <= 12'h2e6;
        src115 <= 12'h3e9;
        src116 <= 12'h954;
        src117 <= 12'h9e;
        src118 <= 12'h8e7;
        src119 <= 12'hc9a;
        src120 <= 12'hab9;
        src121 <= 12'hf2e;
        src122 <= 12'he3f;
        src123 <= 12'h20f;
        src124 <= 12'h2dd;
        src125 <= 12'hfd3;
        src126 <= 12'haa5;
        src127 <= 12'h50a;
        exp <= 19'h3f93d;
        #1
        src0 <= 12'hb60;
        src1 <= 12'h40c;
        src2 <= 12'heea;
        src3 <= 12'h124;
        src4 <= 12'h658;
        src5 <= 12'h564;
        src6 <= 12'h336;
        src7 <= 12'h7c;
        src8 <= 12'h2f8;
        src9 <= 12'ha80;
        src10 <= 12'h191;
        src11 <= 12'h19c;
        src12 <= 12'h564;
        src13 <= 12'h7f4;
        src14 <= 12'h3fd;
        src15 <= 12'h377;
        src16 <= 12'h716;
        src17 <= 12'hbf5;
        src18 <= 12'hef9;
        src19 <= 12'h5ff;
        src20 <= 12'h1ff;
        src21 <= 12'h5b4;
        src22 <= 12'h63e;
        src23 <= 12'h6f2;
        src24 <= 12'h9bc;
        src25 <= 12'h1f7;
        src26 <= 12'hb36;
        src27 <= 12'heaa;
        src28 <= 12'h2cf;
        src29 <= 12'h7b0;
        src30 <= 12'h6d0;
        src31 <= 12'h37;
        src32 <= 12'hefe;
        src33 <= 12'h32a;
        src34 <= 12'h36d;
        src35 <= 12'habf;
        src36 <= 12'h8c3;
        src37 <= 12'h24a;
        src38 <= 12'he05;
        src39 <= 12'h4ff;
        src40 <= 12'h28d;
        src41 <= 12'hc72;
        src42 <= 12'he25;
        src43 <= 12'h82a;
        src44 <= 12'h4c0;
        src45 <= 12'hf8c;
        src46 <= 12'h164;
        src47 <= 12'h300;
        src48 <= 12'h8d7;
        src49 <= 12'h432;
        src50 <= 12'h276;
        src51 <= 12'hd0a;
        src52 <= 12'heb2;
        src53 <= 12'hf81;
        src54 <= 12'h4db;
        src55 <= 12'heff;
        src56 <= 12'h209;
        src57 <= 12'h5e0;
        src58 <= 12'he5c;
        src59 <= 12'h875;
        src60 <= 12'h56f;
        src61 <= 12'h30;
        src62 <= 12'hf7;
        src63 <= 12'hf00;
        src64 <= 12'h5f4;
        src65 <= 12'h138;
        src66 <= 12'hdb6;
        src67 <= 12'he16;
        src68 <= 12'h896;
        src69 <= 12'h6f8;
        src70 <= 12'h48d;
        src71 <= 12'ha56;
        src72 <= 12'h76e;
        src73 <= 12'h4eb;
        src74 <= 12'h7e;
        src75 <= 12'hd29;
        src76 <= 12'h5f3;
        src77 <= 12'hd89;
        src78 <= 12'h310;
        src79 <= 12'hee;
        src80 <= 12'h99a;
        src81 <= 12'haf6;
        src82 <= 12'h422;
        src83 <= 12'h17;
        src84 <= 12'h857;
        src85 <= 12'hf66;
        src86 <= 12'hafc;
        src87 <= 12'h48d;
        src88 <= 12'hc36;
        src89 <= 12'hfcb;
        src90 <= 12'h749;
        src91 <= 12'heca;
        src92 <= 12'hbef;
        src93 <= 12'h91d;
        src94 <= 12'h3d7;
        src95 <= 12'hb67;
        src96 <= 12'h64;
        src97 <= 12'hfb0;
        src98 <= 12'hb81;
        src99 <= 12'h336;
        src100 <= 12'h75e;
        src101 <= 12'ha84;
        src102 <= 12'h469;
        src103 <= 12'hfae;
        src104 <= 12'h3a6;
        src105 <= 12'heef;
        src106 <= 12'h8e;
        src107 <= 12'h6b;
        src108 <= 12'h7d4;
        src109 <= 12'h68d;
        src110 <= 12'hc2a;
        src111 <= 12'hd8a;
        src112 <= 12'h338;
        src113 <= 12'h2e0;
        src114 <= 12'h32d;
        src115 <= 12'h672;
        src116 <= 12'ha2c;
        src117 <= 12'h648;
        src118 <= 12'habd;
        src119 <= 12'h14c;
        src120 <= 12'h92f;
        src121 <= 12'hfbf;
        src122 <= 12'h94b;
        src123 <= 12'h906;
        src124 <= 12'h861;
        src125 <= 12'h8b8;
        src126 <= 12'hd55;
        src127 <= 12'ha32;
        exp <= 19'h3d16b;
        #1
        src0 <= 12'hb71;
        src1 <= 12'h863;
        src2 <= 12'h1d4;
        src3 <= 12'h6a6;
        src4 <= 12'h9b8;
        src5 <= 12'h610;
        src6 <= 12'h6e0;
        src7 <= 12'haa3;
        src8 <= 12'h2c7;
        src9 <= 12'he1d;
        src10 <= 12'hbc;
        src11 <= 12'h44d;
        src12 <= 12'haa4;
        src13 <= 12'h4b9;
        src14 <= 12'hbe5;
        src15 <= 12'hce6;
        src16 <= 12'he62;
        src17 <= 12'h893;
        src18 <= 12'h325;
        src19 <= 12'hff6;
        src20 <= 12'h968;
        src21 <= 12'haa;
        src22 <= 12'h1f6;
        src23 <= 12'h537;
        src24 <= 12'h71c;
        src25 <= 12'hc0b;
        src26 <= 12'h3cb;
        src27 <= 12'hdd2;
        src28 <= 12'h73c;
        src29 <= 12'hfc;
        src30 <= 12'h5d8;
        src31 <= 12'h589;
        src32 <= 12'hee9;
        src33 <= 12'h976;
        src34 <= 12'ha5e;
        src35 <= 12'hf35;
        src36 <= 12'h942;
        src37 <= 12'h3d9;
        src38 <= 12'h1ef;
        src39 <= 12'hbb6;
        src40 <= 12'h1dd;
        src41 <= 12'hef9;
        src42 <= 12'hac5;
        src43 <= 12'hd02;
        src44 <= 12'h983;
        src45 <= 12'hebe;
        src46 <= 12'he02;
        src47 <= 12'hd94;
        src48 <= 12'h737;
        src49 <= 12'hdd3;
        src50 <= 12'hb3a;
        src51 <= 12'ha35;
        src52 <= 12'h6e5;
        src53 <= 12'h5e7;
        src54 <= 12'haac;
        src55 <= 12'h231;
        src56 <= 12'h625;
        src57 <= 12'he8;
        src58 <= 12'h24;
        src59 <= 12'h617;
        src60 <= 12'hb62;
        src61 <= 12'hc1b;
        src62 <= 12'h1c2;
        src63 <= 12'hc01;
        src64 <= 12'h7c1;
        src65 <= 12'he0d;
        src66 <= 12'h1;
        src67 <= 12'h6e6;
        src68 <= 12'h9d5;
        src69 <= 12'h39d;
        src70 <= 12'ha93;
        src71 <= 12'h82b;
        src72 <= 12'h837;
        src73 <= 12'hd52;
        src74 <= 12'h9f5;
        src75 <= 12'h372;
        src76 <= 12'h803;
        src77 <= 12'h6c7;
        src78 <= 12'h3fa;
        src79 <= 12'h49a;
        src80 <= 12'h2d3;
        src81 <= 12'h118;
        src82 <= 12'hed1;
        src83 <= 12'h297;
        src84 <= 12'h1ef;
        src85 <= 12'hc0e;
        src86 <= 12'hc88;
        src87 <= 12'h605;
        src88 <= 12'hb0b;
        src89 <= 12'h3a9;
        src90 <= 12'h98c;
        src91 <= 12'hb30;
        src92 <= 12'h7ed;
        src93 <= 12'hd17;
        src94 <= 12'h2df;
        src95 <= 12'he9f;
        src96 <= 12'h755;
        src97 <= 12'hde5;
        src98 <= 12'h24e;
        src99 <= 12'h18c;
        src100 <= 12'h2d1;
        src101 <= 12'h3d4;
        src102 <= 12'hd9d;
        src103 <= 12'hcd3;
        src104 <= 12'hfd4;
        src105 <= 12'h828;
        src106 <= 12'hbb4;
        src107 <= 12'h8d3;
        src108 <= 12'hd60;
        src109 <= 12'h791;
        src110 <= 12'hdc5;
        src111 <= 12'h726;
        src112 <= 12'h181;
        src113 <= 12'he26;
        src114 <= 12'hde4;
        src115 <= 12'h67b;
        src116 <= 12'h599;
        src117 <= 12'heb0;
        src118 <= 12'hef5;
        src119 <= 12'h21b;
        src120 <= 12'h927;
        src121 <= 12'hdfe;
        src122 <= 12'h59e;
        src123 <= 12'h348;
        src124 <= 12'h2d4;
        src125 <= 12'h4ed;
        src126 <= 12'hc51;
        src127 <= 12'h8bd;
        exp <= 19'h41ced;
        #1
        src0 <= 12'hada;
        src1 <= 12'h3a;
        src2 <= 12'h26f;
        src3 <= 12'h2f6;
        src4 <= 12'h5d;
        src5 <= 12'hce7;
        src6 <= 12'h2b2;
        src7 <= 12'h42c;
        src8 <= 12'hea7;
        src9 <= 12'h49b;
        src10 <= 12'he1f;
        src11 <= 12'h26b;
        src12 <= 12'h75c;
        src13 <= 12'h89a;
        src14 <= 12'h255;
        src15 <= 12'h669;
        src16 <= 12'h6cf;
        src17 <= 12'h8c;
        src18 <= 12'h91d;
        src19 <= 12'hbc9;
        src20 <= 12'h9cc;
        src21 <= 12'haa7;
        src22 <= 12'haca;
        src23 <= 12'ha47;
        src24 <= 12'h635;
        src25 <= 12'hc8e;
        src26 <= 12'h5cd;
        src27 <= 12'hbea;
        src28 <= 12'h3c;
        src29 <= 12'h806;
        src30 <= 12'h9a5;
        src31 <= 12'h3e6;
        src32 <= 12'ha53;
        src33 <= 12'h70c;
        src34 <= 12'hac6;
        src35 <= 12'h898;
        src36 <= 12'hb04;
        src37 <= 12'hbe1;
        src38 <= 12'hc1d;
        src39 <= 12'h6f3;
        src40 <= 12'h4b9;
        src41 <= 12'h55a;
        src42 <= 12'h8bc;
        src43 <= 12'hc85;
        src44 <= 12'h327;
        src45 <= 12'hf3f;
        src46 <= 12'hf2b;
        src47 <= 12'h57f;
        src48 <= 12'hf47;
        src49 <= 12'h725;
        src50 <= 12'h4b5;
        src51 <= 12'hbad;
        src52 <= 12'hc6c;
        src53 <= 12'hadf;
        src54 <= 12'hc20;
        src55 <= 12'h629;
        src56 <= 12'h485;
        src57 <= 12'h404;
        src58 <= 12'hf83;
        src59 <= 12'h7e6;
        src60 <= 12'hd57;
        src61 <= 12'h89f;
        src62 <= 12'h950;
        src63 <= 12'h643;
        src64 <= 12'h3da;
        src65 <= 12'hc6;
        src66 <= 12'h99e;
        src67 <= 12'h6d2;
        src68 <= 12'h6b7;
        src69 <= 12'h97c;
        src70 <= 12'hf4a;
        src71 <= 12'h358;
        src72 <= 12'h3de;
        src73 <= 12'hf95;
        src74 <= 12'h245;
        src75 <= 12'he4b;
        src76 <= 12'h364;
        src77 <= 12'hf49;
        src78 <= 12'h507;
        src79 <= 12'h318;
        src80 <= 12'h8ca;
        src81 <= 12'haec;
        src82 <= 12'h529;
        src83 <= 12'h228;
        src84 <= 12'h533;
        src85 <= 12'h6a2;
        src86 <= 12'haab;
        src87 <= 12'h811;
        src88 <= 12'hcd1;
        src89 <= 12'hb29;
        src90 <= 12'h8be;
        src91 <= 12'h980;
        src92 <= 12'hc1;
        src93 <= 12'hc10;
        src94 <= 12'h9e9;
        src95 <= 12'h442;
        src96 <= 12'hf35;
        src97 <= 12'h12c;
        src98 <= 12'h6ad;
        src99 <= 12'hcf5;
        src100 <= 12'hd37;
        src101 <= 12'h6a6;
        src102 <= 12'h5f;
        src103 <= 12'hcae;
        src104 <= 12'h7e6;
        src105 <= 12'hf1c;
        src106 <= 12'h21b;
        src107 <= 12'ha1a;
        src108 <= 12'h861;
        src109 <= 12'hcf;
        src110 <= 12'hac8;
        src111 <= 12'ha86;
        src112 <= 12'h826;
        src113 <= 12'h512;
        src114 <= 12'h694;
        src115 <= 12'h8b;
        src116 <= 12'h21;
        src117 <= 12'ha51;
        src118 <= 12'h79c;
        src119 <= 12'h367;
        src120 <= 12'h666;
        src121 <= 12'hee;
        src122 <= 12'h638;
        src123 <= 12'hc32;
        src124 <= 12'h1b3;
        src125 <= 12'h870;
        src126 <= 12'h874;
        src127 <= 12'h18e;
        exp <= 19'h3dfeb;
        #1
        src0 <= 12'h739;
        src1 <= 12'hf39;
        src2 <= 12'hd2d;
        src3 <= 12'heb0;
        src4 <= 12'h759;
        src5 <= 12'h27b;
        src6 <= 12'h3f3;
        src7 <= 12'hcd9;
        src8 <= 12'hde1;
        src9 <= 12'h49;
        src10 <= 12'h477;
        src11 <= 12'hd7d;
        src12 <= 12'h713;
        src13 <= 12'he8a;
        src14 <= 12'hbb;
        src15 <= 12'h535;
        src16 <= 12'h444;
        src17 <= 12'he55;
        src18 <= 12'h42d;
        src19 <= 12'ha8f;
        src20 <= 12'h75;
        src21 <= 12'h57;
        src22 <= 12'hf92;
        src23 <= 12'h43;
        src24 <= 12'h313;
        src25 <= 12'hcd6;
        src26 <= 12'h3ee;
        src27 <= 12'h631;
        src28 <= 12'h52a;
        src29 <= 12'h5ed;
        src30 <= 12'h81a;
        src31 <= 12'hcd8;
        src32 <= 12'h97c;
        src33 <= 12'h9b6;
        src34 <= 12'h11f;
        src35 <= 12'h618;
        src36 <= 12'hed;
        src37 <= 12'ha71;
        src38 <= 12'h4fd;
        src39 <= 12'h886;
        src40 <= 12'h23f;
        src41 <= 12'hab0;
        src42 <= 12'h604;
        src43 <= 12'h6c8;
        src44 <= 12'hf5b;
        src45 <= 12'ha30;
        src46 <= 12'hccb;
        src47 <= 12'h896;
        src48 <= 12'hb5;
        src49 <= 12'h8a3;
        src50 <= 12'h6e7;
        src51 <= 12'h620;
        src52 <= 12'h6ff;
        src53 <= 12'h80d;
        src54 <= 12'hafa;
        src55 <= 12'ha86;
        src56 <= 12'hfb8;
        src57 <= 12'ha9b;
        src58 <= 12'h16c;
        src59 <= 12'hcef;
        src60 <= 12'h56;
        src61 <= 12'heb4;
        src62 <= 12'h2ad;
        src63 <= 12'h986;
        src64 <= 12'h736;
        src65 <= 12'hf54;
        src66 <= 12'h641;
        src67 <= 12'h302;
        src68 <= 12'h451;
        src69 <= 12'h804;
        src70 <= 12'h86b;
        src71 <= 12'h9e4;
        src72 <= 12'hd09;
        src73 <= 12'h7bc;
        src74 <= 12'h409;
        src75 <= 12'hf;
        src76 <= 12'h8c9;
        src77 <= 12'h4a5;
        src78 <= 12'h65d;
        src79 <= 12'h9ce;
        src80 <= 12'h97f;
        src81 <= 12'hdd0;
        src82 <= 12'hdc3;
        src83 <= 12'hbb6;
        src84 <= 12'h51;
        src85 <= 12'h19;
        src86 <= 12'hb10;
        src87 <= 12'hb7;
        src88 <= 12'hf74;
        src89 <= 12'hac9;
        src90 <= 12'hd75;
        src91 <= 12'ha38;
        src92 <= 12'hc2b;
        src93 <= 12'h42e;
        src94 <= 12'h1b;
        src95 <= 12'hf15;
        src96 <= 12'h73b;
        src97 <= 12'hae6;
        src98 <= 12'habb;
        src99 <= 12'hdfe;
        src100 <= 12'h811;
        src101 <= 12'h68e;
        src102 <= 12'h3cb;
        src103 <= 12'hf9c;
        src104 <= 12'hb93;
        src105 <= 12'h652;
        src106 <= 12'h44a;
        src107 <= 12'hd4c;
        src108 <= 12'h65c;
        src109 <= 12'h3ed;
        src110 <= 12'h5e3;
        src111 <= 12'ha4a;
        src112 <= 12'hcd7;
        src113 <= 12'h898;
        src114 <= 12'he64;
        src115 <= 12'haa0;
        src116 <= 12'ha1d;
        src117 <= 12'h206;
        src118 <= 12'h5a;
        src119 <= 12'h528;
        src120 <= 12'h7e7;
        src121 <= 12'h5b8;
        src122 <= 12'h86;
        src123 <= 12'h232;
        src124 <= 12'he9f;
        src125 <= 12'h303;
        src126 <= 12'h5cc;
        src127 <= 12'h97e;
        exp <= 19'h3eee7;
        #1
        src0 <= 12'h17;
        src1 <= 12'h71d;
        src2 <= 12'h934;
        src3 <= 12'hb6b;
        src4 <= 12'h261;
        src5 <= 12'h260;
        src6 <= 12'hfec;
        src7 <= 12'h285;
        src8 <= 12'h90d;
        src9 <= 12'hed9;
        src10 <= 12'h164;
        src11 <= 12'h996;
        src12 <= 12'h476;
        src13 <= 12'hb78;
        src14 <= 12'hd82;
        src15 <= 12'h44a;
        src16 <= 12'hefd;
        src17 <= 12'h19d;
        src18 <= 12'h2e1;
        src19 <= 12'hdb1;
        src20 <= 12'hb3;
        src21 <= 12'h20e;
        src22 <= 12'h4b4;
        src23 <= 12'hc71;
        src24 <= 12'h5e8;
        src25 <= 12'he1f;
        src26 <= 12'h122;
        src27 <= 12'h53f;
        src28 <= 12'hd7c;
        src29 <= 12'h45d;
        src30 <= 12'h807;
        src31 <= 12'h418;
        src32 <= 12'hb75;
        src33 <= 12'h503;
        src34 <= 12'hdcf;
        src35 <= 12'h19;
        src36 <= 12'hf66;
        src37 <= 12'h4fb;
        src38 <= 12'h61;
        src39 <= 12'h1aa;
        src40 <= 12'h380;
        src41 <= 12'h1d3;
        src42 <= 12'h104;
        src43 <= 12'h361;
        src44 <= 12'h687;
        src45 <= 12'h478;
        src46 <= 12'h2a8;
        src47 <= 12'hbd3;
        src48 <= 12'hb9;
        src49 <= 12'hd53;
        src50 <= 12'he6f;
        src51 <= 12'hc;
        src52 <= 12'h5b6;
        src53 <= 12'hea0;
        src54 <= 12'h78;
        src55 <= 12'hf0e;
        src56 <= 12'h59b;
        src57 <= 12'ha05;
        src58 <= 12'hc9a;
        src59 <= 12'hec6;
        src60 <= 12'h8f;
        src61 <= 12'hdcf;
        src62 <= 12'h95c;
        src63 <= 12'hcc9;
        src64 <= 12'hc51;
        src65 <= 12'h4b9;
        src66 <= 12'h619;
        src67 <= 12'h1c5;
        src68 <= 12'hab7;
        src69 <= 12'h375;
        src70 <= 12'hcdd;
        src71 <= 12'ha24;
        src72 <= 12'h5d9;
        src73 <= 12'h5b1;
        src74 <= 12'hc0a;
        src75 <= 12'h826;
        src76 <= 12'he3c;
        src77 <= 12'h8d3;
        src78 <= 12'hb98;
        src79 <= 12'ha5a;
        src80 <= 12'h56d;
        src81 <= 12'h101;
        src82 <= 12'hc78;
        src83 <= 12'h564;
        src84 <= 12'h7;
        src85 <= 12'hfe2;
        src86 <= 12'hcc9;
        src87 <= 12'h48f;
        src88 <= 12'h6e0;
        src89 <= 12'hf6e;
        src90 <= 12'he78;
        src91 <= 12'h8af;
        src92 <= 12'h2b;
        src93 <= 12'h11d;
        src94 <= 12'h6b3;
        src95 <= 12'h6b3;
        src96 <= 12'h4e5;
        src97 <= 12'hff9;
        src98 <= 12'h1a7;
        src99 <= 12'hb33;
        src100 <= 12'hd95;
        src101 <= 12'h855;
        src102 <= 12'h80f;
        src103 <= 12'he55;
        src104 <= 12'heee;
        src105 <= 12'h147;
        src106 <= 12'hf9a;
        src107 <= 12'hd42;
        src108 <= 12'hc81;
        src109 <= 12'h7a7;
        src110 <= 12'hf18;
        src111 <= 12'hbf0;
        src112 <= 12'hc9e;
        src113 <= 12'h78e;
        src114 <= 12'h681;
        src115 <= 12'h772;
        src116 <= 12'h29d;
        src117 <= 12'h1a6;
        src118 <= 12'h719;
        src119 <= 12'hd94;
        src120 <= 12'h543;
        src121 <= 12'h25b;
        src122 <= 12'h394;
        src123 <= 12'hf26;
        src124 <= 12'hd52;
        src125 <= 12'h4e0;
        src126 <= 12'h6be;
        src127 <= 12'h8b2;
        exp <= 19'h3eec3;
        #1
        src0 <= 12'h3d1;
        src1 <= 12'hbe0;
        src2 <= 12'he3;
        src3 <= 12'hb;
        src4 <= 12'h8e;
        src5 <= 12'h56b;
        src6 <= 12'hf3c;
        src7 <= 12'hda;
        src8 <= 12'h835;
        src9 <= 12'h1f;
        src10 <= 12'h364;
        src11 <= 12'h79a;
        src12 <= 12'h570;
        src13 <= 12'hc8b;
        src14 <= 12'h1b9;
        src15 <= 12'h1bb;
        src16 <= 12'h613;
        src17 <= 12'h653;
        src18 <= 12'h5f5;
        src19 <= 12'h3b0;
        src20 <= 12'hfe2;
        src21 <= 12'h55b;
        src22 <= 12'h376;
        src23 <= 12'h6d1;
        src24 <= 12'hf97;
        src25 <= 12'h497;
        src26 <= 12'hcfc;
        src27 <= 12'h74c;
        src28 <= 12'hef5;
        src29 <= 12'h3b4;
        src30 <= 12'hda7;
        src31 <= 12'h1a5;
        src32 <= 12'h320;
        src33 <= 12'he3a;
        src34 <= 12'hddb;
        src35 <= 12'h2c1;
        src36 <= 12'h794;
        src37 <= 12'h7dd;
        src38 <= 12'hc1e;
        src39 <= 12'he9f;
        src40 <= 12'h27;
        src41 <= 12'h69e;
        src42 <= 12'he00;
        src43 <= 12'h6c8;
        src44 <= 12'h708;
        src45 <= 12'hc33;
        src46 <= 12'h42b;
        src47 <= 12'h895;
        src48 <= 12'h9e5;
        src49 <= 12'h763;
        src50 <= 12'h8d;
        src51 <= 12'h393;
        src52 <= 12'hcbb;
        src53 <= 12'hd87;
        src54 <= 12'hf8b;
        src55 <= 12'h360;
        src56 <= 12'hdb1;
        src57 <= 12'ha70;
        src58 <= 12'h537;
        src59 <= 12'h644;
        src60 <= 12'hae0;
        src61 <= 12'hb1d;
        src62 <= 12'h5cf;
        src63 <= 12'hdec;
        src64 <= 12'hfcd;
        src65 <= 12'hce7;
        src66 <= 12'h968;
        src67 <= 12'h272;
        src68 <= 12'hee3;
        src69 <= 12'hf27;
        src70 <= 12'h5c9;
        src71 <= 12'hb79;
        src72 <= 12'hb54;
        src73 <= 12'h452;
        src74 <= 12'hc33;
        src75 <= 12'hb7;
        src76 <= 12'hf55;
        src77 <= 12'h214;
        src78 <= 12'h8f8;
        src79 <= 12'h694;
        src80 <= 12'h311;
        src81 <= 12'h188;
        src82 <= 12'hf2b;
        src83 <= 12'h67e;
        src84 <= 12'h2a1;
        src85 <= 12'h6b9;
        src86 <= 12'hb21;
        src87 <= 12'heb;
        src88 <= 12'h1ab;
        src89 <= 12'h8bc;
        src90 <= 12'h83c;
        src91 <= 12'hbb0;
        src92 <= 12'h8d7;
        src93 <= 12'h65e;
        src94 <= 12'h1b6;
        src95 <= 12'h44d;
        src96 <= 12'h1ac;
        src97 <= 12'h498;
        src98 <= 12'h525;
        src99 <= 12'h38f;
        src100 <= 12'h349;
        src101 <= 12'hfbc;
        src102 <= 12'hab0;
        src103 <= 12'h52a;
        src104 <= 12'h77b;
        src105 <= 12'hcc7;
        src106 <= 12'hca5;
        src107 <= 12'h19c;
        src108 <= 12'h4a3;
        src109 <= 12'h133;
        src110 <= 12'hd87;
        src111 <= 12'h281;
        src112 <= 12'hbb8;
        src113 <= 12'h7f;
        src114 <= 12'h580;
        src115 <= 12'hbaa;
        src116 <= 12'h630;
        src117 <= 12'h521;
        src118 <= 12'h2f1;
        src119 <= 12'he1d;
        src120 <= 12'he90;
        src121 <= 12'ha16;
        src122 <= 12'he4d;
        src123 <= 12'he04;
        src124 <= 12'h580;
        src125 <= 12'hd71;
        src126 <= 12'h215;
        src127 <= 12'h8e7;
        exp <= 19'h3d66c;
        #1
        src0 <= 12'h27a;
        src1 <= 12'h679;
        src2 <= 12'hf01;
        src3 <= 12'h249;
        src4 <= 12'h489;
        src5 <= 12'hcb4;
        src6 <= 12'hebf;
        src7 <= 12'ha17;
        src8 <= 12'hf92;
        src9 <= 12'heab;
        src10 <= 12'hb49;
        src11 <= 12'h5e;
        src12 <= 12'h368;
        src13 <= 12'hbc3;
        src14 <= 12'h35c;
        src15 <= 12'h36b;
        src16 <= 12'h7e9;
        src17 <= 12'h91f;
        src18 <= 12'h7e7;
        src19 <= 12'h118;
        src20 <= 12'h2dc;
        src21 <= 12'h939;
        src22 <= 12'h213;
        src23 <= 12'hcfa;
        src24 <= 12'h1a9;
        src25 <= 12'h63f;
        src26 <= 12'hd6c;
        src27 <= 12'h812;
        src28 <= 12'h189;
        src29 <= 12'hb92;
        src30 <= 12'h655;
        src31 <= 12'he0e;
        src32 <= 12'hfbd;
        src33 <= 12'h4b7;
        src34 <= 12'h8d8;
        src35 <= 12'h536;
        src36 <= 12'h618;
        src37 <= 12'ha2e;
        src38 <= 12'h621;
        src39 <= 12'h7ca;
        src40 <= 12'h411;
        src41 <= 12'h42;
        src42 <= 12'h26c;
        src43 <= 12'ha67;
        src44 <= 12'h6cf;
        src45 <= 12'h8b9;
        src46 <= 12'h956;
        src47 <= 12'hfc5;
        src48 <= 12'hea;
        src49 <= 12'ha5b;
        src50 <= 12'h58e;
        src51 <= 12'h32a;
        src52 <= 12'h9fc;
        src53 <= 12'hbf0;
        src54 <= 12'h6ea;
        src55 <= 12'h865;
        src56 <= 12'h869;
        src57 <= 12'he7c;
        src58 <= 12'hb14;
        src59 <= 12'h667;
        src60 <= 12'h80c;
        src61 <= 12'he53;
        src62 <= 12'hb2a;
        src63 <= 12'h948;
        src64 <= 12'hf34;
        src65 <= 12'hac8;
        src66 <= 12'hfe8;
        src67 <= 12'h5b8;
        src68 <= 12'h844;
        src69 <= 12'hbc0;
        src70 <= 12'h1ee;
        src71 <= 12'h332;
        src72 <= 12'hec9;
        src73 <= 12'h56d;
        src74 <= 12'hc99;
        src75 <= 12'hb02;
        src76 <= 12'hae5;
        src77 <= 12'hee0;
        src78 <= 12'h257;
        src79 <= 12'h7db;
        src80 <= 12'hbc0;
        src81 <= 12'h295;
        src82 <= 12'h96c;
        src83 <= 12'ha60;
        src84 <= 12'heaf;
        src85 <= 12'h945;
        src86 <= 12'h328;
        src87 <= 12'h97f;
        src88 <= 12'h9e9;
        src89 <= 12'ha2d;
        src90 <= 12'hd04;
        src91 <= 12'h692;
        src92 <= 12'h777;
        src93 <= 12'h5e1;
        src94 <= 12'he4b;
        src95 <= 12'h859;
        src96 <= 12'h8ad;
        src97 <= 12'h7eb;
        src98 <= 12'h66d;
        src99 <= 12'h907;
        src100 <= 12'hcf0;
        src101 <= 12'h605;
        src102 <= 12'hdc;
        src103 <= 12'hd51;
        src104 <= 12'h823;
        src105 <= 12'h7f5;
        src106 <= 12'h821;
        src107 <= 12'h374;
        src108 <= 12'hdda;
        src109 <= 12'h98a;
        src110 <= 12'hf41;
        src111 <= 12'h4a8;
        src112 <= 12'h564;
        src113 <= 12'h2fc;
        src114 <= 12'he73;
        src115 <= 12'hb83;
        src116 <= 12'hb31;
        src117 <= 12'h194;
        src118 <= 12'ha60;
        src119 <= 12'haf8;
        src120 <= 12'h740;
        src121 <= 12'h987;
        src122 <= 12'h13;
        src123 <= 12'ha70;
        src124 <= 12'h584;
        src125 <= 12'ha46;
        src126 <= 12'hb9b;
        src127 <= 12'h595;
        exp <= 19'h432e3;
        #1
        src0 <= 12'h51b;
        src1 <= 12'h300;
        src2 <= 12'hafc;
        src3 <= 12'hf4;
        src4 <= 12'h3e6;
        src5 <= 12'hd4f;
        src6 <= 12'h20e;
        src7 <= 12'habd;
        src8 <= 12'h552;
        src9 <= 12'h767;
        src10 <= 12'h6f5;
        src11 <= 12'hbab;
        src12 <= 12'hcc1;
        src13 <= 12'ha60;
        src14 <= 12'haed;
        src15 <= 12'h7df;
        src16 <= 12'hfed;
        src17 <= 12'h207;
        src18 <= 12'he6a;
        src19 <= 12'hb26;
        src20 <= 12'h322;
        src21 <= 12'he85;
        src22 <= 12'h172;
        src23 <= 12'hbec;
        src24 <= 12'hb0;
        src25 <= 12'h2b2;
        src26 <= 12'he3e;
        src27 <= 12'h3e0;
        src28 <= 12'hb42;
        src29 <= 12'hc25;
        src30 <= 12'he61;
        src31 <= 12'h186;
        src32 <= 12'h304;
        src33 <= 12'h5d3;
        src34 <= 12'h58b;
        src35 <= 12'h649;
        src36 <= 12'hcf5;
        src37 <= 12'hbf;
        src38 <= 12'he40;
        src39 <= 12'h73e;
        src40 <= 12'hd38;
        src41 <= 12'h7e;
        src42 <= 12'hc5;
        src43 <= 12'h3;
        src44 <= 12'hc73;
        src45 <= 12'h310;
        src46 <= 12'hd6b;
        src47 <= 12'h706;
        src48 <= 12'hdc0;
        src49 <= 12'hb96;
        src50 <= 12'hc0f;
        src51 <= 12'h338;
        src52 <= 12'h282;
        src53 <= 12'hdb;
        src54 <= 12'h5dc;
        src55 <= 12'hb9c;
        src56 <= 12'ha57;
        src57 <= 12'h560;
        src58 <= 12'h474;
        src59 <= 12'hbff;
        src60 <= 12'h1d2;
        src61 <= 12'h85;
        src62 <= 12'h6f7;
        src63 <= 12'h9b3;
        src64 <= 12'h9e6;
        src65 <= 12'h514;
        src66 <= 12'h27f;
        src67 <= 12'h10e;
        src68 <= 12'h594;
        src69 <= 12'hba1;
        src70 <= 12'h444;
        src71 <= 12'h4b0;
        src72 <= 12'hc87;
        src73 <= 12'h48c;
        src74 <= 12'h8b1;
        src75 <= 12'h1e5;
        src76 <= 12'h812;
        src77 <= 12'h195;
        src78 <= 12'h710;
        src79 <= 12'hdc9;
        src80 <= 12'h4db;
        src81 <= 12'had6;
        src82 <= 12'hca6;
        src83 <= 12'h6f2;
        src84 <= 12'h72;
        src85 <= 12'h782;
        src86 <= 12'hdcc;
        src87 <= 12'h5f2;
        src88 <= 12'h4ae;
        src89 <= 12'h5d9;
        src90 <= 12'hef1;
        src91 <= 12'h5a0;
        src92 <= 12'hee0;
        src93 <= 12'h6d9;
        src94 <= 12'h93f;
        src95 <= 12'hd9;
        src96 <= 12'h48e;
        src97 <= 12'hf73;
        src98 <= 12'h592;
        src99 <= 12'h64d;
        src100 <= 12'h2d1;
        src101 <= 12'h634;
        src102 <= 12'h13f;
        src103 <= 12'h6a8;
        src104 <= 12'h28c;
        src105 <= 12'h460;
        src106 <= 12'h2;
        src107 <= 12'hcac;
        src108 <= 12'h970;
        src109 <= 12'h758;
        src110 <= 12'h62a;
        src111 <= 12'h56;
        src112 <= 12'hc06;
        src113 <= 12'hbdb;
        src114 <= 12'h169;
        src115 <= 12'h246;
        src116 <= 12'h6ea;
        src117 <= 12'h75f;
        src118 <= 12'h306;
        src119 <= 12'h96c;
        src120 <= 12'ha56;
        src121 <= 12'h60a;
        src122 <= 12'hc90;
        src123 <= 12'h44e;
        src124 <= 12'h631;
        src125 <= 12'h982;
        src126 <= 12'hb2d;
        src127 <= 12'hac8;
        exp <= 19'h39b30;
        #1
        src0 <= 12'h957;
        src1 <= 12'hf77;
        src2 <= 12'hb4e;
        src3 <= 12'h7da;
        src4 <= 12'h575;
        src5 <= 12'ha6e;
        src6 <= 12'h9bb;
        src7 <= 12'h248;
        src8 <= 12'hcd;
        src9 <= 12'h60d;
        src10 <= 12'h9a5;
        src11 <= 12'h9c4;
        src12 <= 12'he51;
        src13 <= 12'haf9;
        src14 <= 12'hd63;
        src15 <= 12'h478;
        src16 <= 12'h7f1;
        src17 <= 12'hac1;
        src18 <= 12'h724;
        src19 <= 12'h5dd;
        src20 <= 12'h1fd;
        src21 <= 12'hba0;
        src22 <= 12'hd64;
        src23 <= 12'hb30;
        src24 <= 12'h8dd;
        src25 <= 12'h4b2;
        src26 <= 12'h431;
        src27 <= 12'hb31;
        src28 <= 12'he23;
        src29 <= 12'h78f;
        src30 <= 12'h159;
        src31 <= 12'hb9b;
        src32 <= 12'h2f1;
        src33 <= 12'ha8d;
        src34 <= 12'h7ea;
        src35 <= 12'h4de;
        src36 <= 12'hcde;
        src37 <= 12'h761;
        src38 <= 12'h187;
        src39 <= 12'h1fd;
        src40 <= 12'he10;
        src41 <= 12'h97e;
        src42 <= 12'h2c3;
        src43 <= 12'h77f;
        src44 <= 12'h211;
        src45 <= 12'h5b0;
        src46 <= 12'h802;
        src47 <= 12'h86f;
        src48 <= 12'he2;
        src49 <= 12'hf0;
        src50 <= 12'ha09;
        src51 <= 12'h915;
        src52 <= 12'hccb;
        src53 <= 12'hd46;
        src54 <= 12'hab3;
        src55 <= 12'hcd4;
        src56 <= 12'hd01;
        src57 <= 12'h531;
        src58 <= 12'h902;
        src59 <= 12'haea;
        src60 <= 12'h1a3;
        src61 <= 12'hb14;
        src62 <= 12'ha29;
        src63 <= 12'h3eb;
        src64 <= 12'h26;
        src65 <= 12'hc1f;
        src66 <= 12'h7bf;
        src67 <= 12'hb29;
        src68 <= 12'h764;
        src69 <= 12'h830;
        src70 <= 12'h4;
        src71 <= 12'hbf2;
        src72 <= 12'ha3e;
        src73 <= 12'h322;
        src74 <= 12'h923;
        src75 <= 12'hb89;
        src76 <= 12'hafd;
        src77 <= 12'ha74;
        src78 <= 12'h126;
        src79 <= 12'h34a;
        src80 <= 12'h15e;
        src81 <= 12'h90a;
        src82 <= 12'hab8;
        src83 <= 12'h87c;
        src84 <= 12'h87a;
        src85 <= 12'h4fe;
        src86 <= 12'h499;
        src87 <= 12'h51e;
        src88 <= 12'h4b6;
        src89 <= 12'h3eb;
        src90 <= 12'hba3;
        src91 <= 12'hd66;
        src92 <= 12'h408;
        src93 <= 12'h36d;
        src94 <= 12'h349;
        src95 <= 12'hce8;
        src96 <= 12'hca3;
        src97 <= 12'hf16;
        src98 <= 12'heb2;
        src99 <= 12'h590;
        src100 <= 12'h67c;
        src101 <= 12'h4fe;
        src102 <= 12'h62c;
        src103 <= 12'h1bd;
        src104 <= 12'h589;
        src105 <= 12'h9f3;
        src106 <= 12'h58e;
        src107 <= 12'hc6d;
        src108 <= 12'hd0a;
        src109 <= 12'hda;
        src110 <= 12'h33c;
        src111 <= 12'h15f;
        src112 <= 12'h711;
        src113 <= 12'h7f3;
        src114 <= 12'h137;
        src115 <= 12'h19f;
        src116 <= 12'h142;
        src117 <= 12'hf04;
        src118 <= 12'hba7;
        src119 <= 12'ha01;
        src120 <= 12'hac6;
        src121 <= 12'hdf4;
        src122 <= 12'he0;
        src123 <= 12'h939;
        src124 <= 12'hdb5;
        src125 <= 12'he80;
        src126 <= 12'h9d0;
        src127 <= 12'h993;
        exp <= 19'h3ec81;
        #1
        src0 <= 12'h546;
        src1 <= 12'h39;
        src2 <= 12'ha14;
        src3 <= 12'hf18;
        src4 <= 12'h902;
        src5 <= 12'h611;
        src6 <= 12'h8a7;
        src7 <= 12'h294;
        src8 <= 12'h2de;
        src9 <= 12'h195;
        src10 <= 12'hfd1;
        src11 <= 12'h162;
        src12 <= 12'h358;
        src13 <= 12'h523;
        src14 <= 12'h770;
        src15 <= 12'h36e;
        src16 <= 12'h6df;
        src17 <= 12'h119;
        src18 <= 12'h255;
        src19 <= 12'h903;
        src20 <= 12'hfc2;
        src21 <= 12'h267;
        src22 <= 12'ha41;
        src23 <= 12'h71e;
        src24 <= 12'h1b4;
        src25 <= 12'h33b;
        src26 <= 12'hca2;
        src27 <= 12'haed;
        src28 <= 12'hfde;
        src29 <= 12'he50;
        src30 <= 12'h57d;
        src31 <= 12'h43d;
        src32 <= 12'hfe3;
        src33 <= 12'hf8c;
        src34 <= 12'hd1;
        src35 <= 12'h728;
        src36 <= 12'h414;
        src37 <= 12'h8d2;
        src38 <= 12'h3e7;
        src39 <= 12'h18b;
        src40 <= 12'hd58;
        src41 <= 12'h153;
        src42 <= 12'h6fc;
        src43 <= 12'hc3;
        src44 <= 12'hed4;
        src45 <= 12'haa3;
        src46 <= 12'he14;
        src47 <= 12'h8;
        src48 <= 12'haa7;
        src49 <= 12'h854;
        src50 <= 12'h6fd;
        src51 <= 12'hb41;
        src52 <= 12'h426;
        src53 <= 12'he87;
        src54 <= 12'h80e;
        src55 <= 12'h83c;
        src56 <= 12'ha55;
        src57 <= 12'h706;
        src58 <= 12'hf6d;
        src59 <= 12'h9e7;
        src60 <= 12'h589;
        src61 <= 12'hbea;
        src62 <= 12'hc63;
        src63 <= 12'h92e;
        src64 <= 12'h200;
        src65 <= 12'ha2d;
        src66 <= 12'h55f;
        src67 <= 12'hf91;
        src68 <= 12'he31;
        src69 <= 12'h82d;
        src70 <= 12'ha1f;
        src71 <= 12'h715;
        src72 <= 12'hf2e;
        src73 <= 12'hf59;
        src74 <= 12'h867;
        src75 <= 12'h1c3;
        src76 <= 12'h9cf;
        src77 <= 12'hec0;
        src78 <= 12'h761;
        src79 <= 12'h82;
        src80 <= 12'h477;
        src81 <= 12'hd9c;
        src82 <= 12'h952;
        src83 <= 12'h762;
        src84 <= 12'h572;
        src85 <= 12'h53d;
        src86 <= 12'h1c3;
        src87 <= 12'he7;
        src88 <= 12'h746;
        src89 <= 12'hb97;
        src90 <= 12'hb27;
        src91 <= 12'h546;
        src92 <= 12'h83d;
        src93 <= 12'h90c;
        src94 <= 12'hef7;
        src95 <= 12'hffb;
        src96 <= 12'h5e3;
        src97 <= 12'hb1e;
        src98 <= 12'h28;
        src99 <= 12'h10b;
        src100 <= 12'hd85;
        src101 <= 12'h8ef;
        src102 <= 12'h4f;
        src103 <= 12'h248;
        src104 <= 12'h56;
        src105 <= 12'hc60;
        src106 <= 12'h7fa;
        src107 <= 12'h8a0;
        src108 <= 12'hda0;
        src109 <= 12'hfcd;
        src110 <= 12'h62b;
        src111 <= 12'h488;
        src112 <= 12'h8bf;
        src113 <= 12'h104;
        src114 <= 12'h75d;
        src115 <= 12'h371;
        src116 <= 12'heaa;
        src117 <= 12'h478;
        src118 <= 12'h9f8;
        src119 <= 12'h499;
        src120 <= 12'hbdb;
        src121 <= 12'h5de;
        src122 <= 12'h325;
        src123 <= 12'hb2a;
        src124 <= 12'h12b;
        src125 <= 12'hdb2;
        src126 <= 12'h5dd;
        src127 <= 12'h530;
        exp <= 19'h3e532;
        #1
        src0 <= 12'h1c9;
        src1 <= 12'he3;
        src2 <= 12'h196;
        src3 <= 12'h663;
        src4 <= 12'h548;
        src5 <= 12'ha2a;
        src6 <= 12'h6d3;
        src7 <= 12'hdb0;
        src8 <= 12'hfc3;
        src9 <= 12'h4a6;
        src10 <= 12'h95;
        src11 <= 12'h5c5;
        src12 <= 12'haed;
        src13 <= 12'h966;
        src14 <= 12'hf2b;
        src15 <= 12'hf50;
        src16 <= 12'hebf;
        src17 <= 12'h6c0;
        src18 <= 12'hc1e;
        src19 <= 12'h7a2;
        src20 <= 12'h187;
        src21 <= 12'h987;
        src22 <= 12'h657;
        src23 <= 12'hea2;
        src24 <= 12'hee9;
        src25 <= 12'h2bd;
        src26 <= 12'he46;
        src27 <= 12'hb8e;
        src28 <= 12'h616;
        src29 <= 12'h581;
        src30 <= 12'h3c;
        src31 <= 12'h446;
        src32 <= 12'h1d6;
        src33 <= 12'he7a;
        src34 <= 12'h9bd;
        src35 <= 12'hf12;
        src36 <= 12'h188;
        src37 <= 12'h4b;
        src38 <= 12'h77a;
        src39 <= 12'haf1;
        src40 <= 12'h86d;
        src41 <= 12'h667;
        src42 <= 12'h9fa;
        src43 <= 12'hc2d;
        src44 <= 12'hbeb;
        src45 <= 12'hbd8;
        src46 <= 12'h24;
        src47 <= 12'hc4c;
        src48 <= 12'h853;
        src49 <= 12'h387;
        src50 <= 12'hb;
        src51 <= 12'h38c;
        src52 <= 12'h5ef;
        src53 <= 12'h9aa;
        src54 <= 12'hcc6;
        src55 <= 12'h11a;
        src56 <= 12'hd70;
        src57 <= 12'hc9f;
        src58 <= 12'hb26;
        src59 <= 12'h846;
        src60 <= 12'hc0;
        src61 <= 12'h215;
        src62 <= 12'hf26;
        src63 <= 12'h7e3;
        src64 <= 12'h809;
        src65 <= 12'hc8;
        src66 <= 12'h777;
        src67 <= 12'h989;
        src68 <= 12'h4a7;
        src69 <= 12'h412;
        src70 <= 12'h8f2;
        src71 <= 12'h5ce;
        src72 <= 12'hbf6;
        src73 <= 12'h186;
        src74 <= 12'hc5b;
        src75 <= 12'hf18;
        src76 <= 12'hb29;
        src77 <= 12'hcc;
        src78 <= 12'h27b;
        src79 <= 12'hf0c;
        src80 <= 12'h488;
        src81 <= 12'hde6;
        src82 <= 12'hce2;
        src83 <= 12'h707;
        src84 <= 12'he3d;
        src85 <= 12'hd0b;
        src86 <= 12'h7df;
        src87 <= 12'h579;
        src88 <= 12'h4e3;
        src89 <= 12'h301;
        src90 <= 12'h51c;
        src91 <= 12'h458;
        src92 <= 12'h832;
        src93 <= 12'h655;
        src94 <= 12'hc31;
        src95 <= 12'h863;
        src96 <= 12'h85f;
        src97 <= 12'h653;
        src98 <= 12'h839;
        src99 <= 12'ha61;
        src100 <= 12'h582;
        src101 <= 12'h995;
        src102 <= 12'hc3f;
        src103 <= 12'h94f;
        src104 <= 12'h51c;
        src105 <= 12'h65a;
        src106 <= 12'h1f8;
        src107 <= 12'h478;
        src108 <= 12'ha4d;
        src109 <= 12'he24;
        src110 <= 12'h9fa;
        src111 <= 12'hefb;
        src112 <= 12'hff;
        src113 <= 12'h259;
        src114 <= 12'h5c8;
        src115 <= 12'h76b;
        src116 <= 12'h14e;
        src117 <= 12'hcff;
        src118 <= 12'ha40;
        src119 <= 12'hb8c;
        src120 <= 12'had2;
        src121 <= 12'h2f;
        src122 <= 12'hc71;
        src123 <= 12'h580;
        src124 <= 12'h24;
        src125 <= 12'he22;
        src126 <= 12'h3c4;
        src127 <= 12'h644;
        exp <= 19'h3ea12;
        #1
        src0 <= 12'hb3;
        src1 <= 12'hc38;
        src2 <= 12'hc19;
        src3 <= 12'h81e;
        src4 <= 12'hd16;
        src5 <= 12'hcbc;
        src6 <= 12'h169;
        src7 <= 12'he22;
        src8 <= 12'h345;
        src9 <= 12'h277;
        src10 <= 12'h22f;
        src11 <= 12'h15f;
        src12 <= 12'hdfe;
        src13 <= 12'h7e5;
        src14 <= 12'h8ef;
        src15 <= 12'h8e5;
        src16 <= 12'h613;
        src17 <= 12'h602;
        src18 <= 12'h3e6;
        src19 <= 12'h86c;
        src20 <= 12'h831;
        src21 <= 12'h4ae;
        src22 <= 12'h822;
        src23 <= 12'h603;
        src24 <= 12'h3f1;
        src25 <= 12'h5b2;
        src26 <= 12'h8ce;
        src27 <= 12'h60e;
        src28 <= 12'ha80;
        src29 <= 12'hee;
        src30 <= 12'he69;
        src31 <= 12'h628;
        src32 <= 12'ha51;
        src33 <= 12'h857;
        src34 <= 12'ha58;
        src35 <= 12'h435;
        src36 <= 12'h497;
        src37 <= 12'h823;
        src38 <= 12'h26b;
        src39 <= 12'ha11;
        src40 <= 12'hfb0;
        src41 <= 12'h860;
        src42 <= 12'hd00;
        src43 <= 12'h28;
        src44 <= 12'hee;
        src45 <= 12'h376;
        src46 <= 12'h331;
        src47 <= 12'hb74;
        src48 <= 12'h160;
        src49 <= 12'h485;
        src50 <= 12'h1a5;
        src51 <= 12'h43;
        src52 <= 12'h597;
        src53 <= 12'h495;
        src54 <= 12'h25d;
        src55 <= 12'hae6;
        src56 <= 12'h512;
        src57 <= 12'ha63;
        src58 <= 12'hd06;
        src59 <= 12'h3fb;
        src60 <= 12'h189;
        src61 <= 12'h197;
        src62 <= 12'hafa;
        src63 <= 12'hab0;
        src64 <= 12'h429;
        src65 <= 12'h758;
        src66 <= 12'h66c;
        src67 <= 12'h60;
        src68 <= 12'hefc;
        src69 <= 12'h5f0;
        src70 <= 12'h6c7;
        src71 <= 12'h127;
        src72 <= 12'h6b2;
        src73 <= 12'hab2;
        src74 <= 12'h10e;
        src75 <= 12'hcc4;
        src76 <= 12'had5;
        src77 <= 12'h9db;
        src78 <= 12'h393;
        src79 <= 12'h329;
        src80 <= 12'h407;
        src81 <= 12'h3cb;
        src82 <= 12'h757;
        src83 <= 12'h521;
        src84 <= 12'h6f3;
        src85 <= 12'hec7;
        src86 <= 12'haea;
        src87 <= 12'hbb5;
        src88 <= 12'hf24;
        src89 <= 12'hd53;
        src90 <= 12'h148;
        src91 <= 12'hdb0;
        src92 <= 12'h9ee;
        src93 <= 12'hd45;
        src94 <= 12'h816;
        src95 <= 12'h65c;
        src96 <= 12'h24d;
        src97 <= 12'h9a7;
        src98 <= 12'h50c;
        src99 <= 12'h30a;
        src100 <= 12'hb73;
        src101 <= 12'h805;
        src102 <= 12'h3a4;
        src103 <= 12'h9d1;
        src104 <= 12'h9f9;
        src105 <= 12'h104;
        src106 <= 12'h7;
        src107 <= 12'hf9b;
        src108 <= 12'h220;
        src109 <= 12'h51b;
        src110 <= 12'h4f7;
        src111 <= 12'h40a;
        src112 <= 12'hc5d;
        src113 <= 12'hbb6;
        src114 <= 12'hecc;
        src115 <= 12'ha75;
        src116 <= 12'h97;
        src117 <= 12'ha9f;
        src118 <= 12'h17;
        src119 <= 12'ha8c;
        src120 <= 12'h98c;
        src121 <= 12'h70f;
        src122 <= 12'h2c7;
        src123 <= 12'h176;
        src124 <= 12'hd35;
        src125 <= 12'h2b1;
        src126 <= 12'h3f6;
        src127 <= 12'h222;
        exp <= 19'h37fe6;
        #1
        src0 <= 12'hf5c;
        src1 <= 12'h3d9;
        src2 <= 12'h3cb;
        src3 <= 12'ha4;
        src4 <= 12'hac1;
        src5 <= 12'h3e0;
        src6 <= 12'h257;
        src7 <= 12'h60b;
        src8 <= 12'h616;
        src9 <= 12'hbe9;
        src10 <= 12'he2f;
        src11 <= 12'h2cd;
        src12 <= 12'h119;
        src13 <= 12'hc3b;
        src14 <= 12'h117;
        src15 <= 12'h607;
        src16 <= 12'h7e;
        src17 <= 12'h746;
        src18 <= 12'h31d;
        src19 <= 12'h75b;
        src20 <= 12'he0a;
        src21 <= 12'h1da;
        src22 <= 12'ha6c;
        src23 <= 12'habb;
        src24 <= 12'h3d1;
        src25 <= 12'h5f7;
        src26 <= 12'he5b;
        src27 <= 12'hc68;
        src28 <= 12'h8fc;
        src29 <= 12'h351;
        src30 <= 12'h892;
        src31 <= 12'h7d2;
        src32 <= 12'h445;
        src33 <= 12'h18a;
        src34 <= 12'h25f;
        src35 <= 12'h36e;
        src36 <= 12'h4a7;
        src37 <= 12'h1fb;
        src38 <= 12'h40f;
        src39 <= 12'h866;
        src40 <= 12'hdb3;
        src41 <= 12'h4f2;
        src42 <= 12'hd8d;
        src43 <= 12'ha6e;
        src44 <= 12'hb8f;
        src45 <= 12'h70a;
        src46 <= 12'h492;
        src47 <= 12'h251;
        src48 <= 12'h921;
        src49 <= 12'haf6;
        src50 <= 12'h219;
        src51 <= 12'h609;
        src52 <= 12'h2d8;
        src53 <= 12'h3fa;
        src54 <= 12'hef2;
        src55 <= 12'hf43;
        src56 <= 12'hf10;
        src57 <= 12'h8ca;
        src58 <= 12'h608;
        src59 <= 12'h18a;
        src60 <= 12'h705;
        src61 <= 12'h685;
        src62 <= 12'h3fd;
        src63 <= 12'hae6;
        src64 <= 12'hc17;
        src65 <= 12'hf2d;
        src66 <= 12'hd82;
        src67 <= 12'h2bb;
        src68 <= 12'hb8;
        src69 <= 12'h260;
        src70 <= 12'hf3f;
        src71 <= 12'hb61;
        src72 <= 12'h1e8;
        src73 <= 12'h49;
        src74 <= 12'hbd8;
        src75 <= 12'h9fa;
        src76 <= 12'h35d;
        src77 <= 12'h482;
        src78 <= 12'h785;
        src79 <= 12'h9d7;
        src80 <= 12'he98;
        src81 <= 12'h4c9;
        src82 <= 12'h9fa;
        src83 <= 12'h6d2;
        src84 <= 12'hbc8;
        src85 <= 12'h848;
        src86 <= 12'h387;
        src87 <= 12'h5ca;
        src88 <= 12'h33c;
        src89 <= 12'h23;
        src90 <= 12'h70d;
        src91 <= 12'h833;
        src92 <= 12'h774;
        src93 <= 12'hb2d;
        src94 <= 12'hf55;
        src95 <= 12'hb94;
        src96 <= 12'h2c5;
        src97 <= 12'h891;
        src98 <= 12'h17c;
        src99 <= 12'ha48;
        src100 <= 12'h427;
        src101 <= 12'h37d;
        src102 <= 12'h1f5;
        src103 <= 12'h278;
        src104 <= 12'h492;
        src105 <= 12'h6b6;
        src106 <= 12'h427;
        src107 <= 12'h96d;
        src108 <= 12'h965;
        src109 <= 12'had0;
        src110 <= 12'hcb4;
        src111 <= 12'h98b;
        src112 <= 12'hf04;
        src113 <= 12'h9c8;
        src114 <= 12'h796;
        src115 <= 12'hc5b;
        src116 <= 12'had1;
        src117 <= 12'h2ea;
        src118 <= 12'hebf;
        src119 <= 12'h6c7;
        src120 <= 12'h38d;
        src121 <= 12'h9b7;
        src122 <= 12'h943;
        src123 <= 12'hfbd;
        src124 <= 12'hc19;
        src125 <= 12'h929;
        src126 <= 12'h1a2;
        src127 <= 12'hba5;
        exp <= 19'h3b9f3;
        #1
        src0 <= 12'hbcf;
        src1 <= 12'h54;
        src2 <= 12'h5ce;
        src3 <= 12'h856;
        src4 <= 12'hfbd;
        src5 <= 12'h2f3;
        src6 <= 12'h477;
        src7 <= 12'hcb5;
        src8 <= 12'h4ca;
        src9 <= 12'hcd4;
        src10 <= 12'h4a;
        src11 <= 12'he6d;
        src12 <= 12'h7d7;
        src13 <= 12'ha1b;
        src14 <= 12'h67e;
        src15 <= 12'h324;
        src16 <= 12'hd2a;
        src17 <= 12'hf66;
        src18 <= 12'h8e;
        src19 <= 12'h555;
        src20 <= 12'h24f;
        src21 <= 12'h474;
        src22 <= 12'hf38;
        src23 <= 12'h9f7;
        src24 <= 12'h6d7;
        src25 <= 12'h36d;
        src26 <= 12'hf31;
        src27 <= 12'h52;
        src28 <= 12'h552;
        src29 <= 12'hdd6;
        src30 <= 12'h3f0;
        src31 <= 12'h4ee;
        src32 <= 12'h5ca;
        src33 <= 12'h296;
        src34 <= 12'hf82;
        src35 <= 12'h7b5;
        src36 <= 12'h790;
        src37 <= 12'h8cd;
        src38 <= 12'hc63;
        src39 <= 12'h3ec;
        src40 <= 12'h62e;
        src41 <= 12'h43b;
        src42 <= 12'h37;
        src43 <= 12'hdd7;
        src44 <= 12'h366;
        src45 <= 12'h9d9;
        src46 <= 12'h6e6;
        src47 <= 12'hd9f;
        src48 <= 12'h118;
        src49 <= 12'hfe0;
        src50 <= 12'hb47;
        src51 <= 12'h2cc;
        src52 <= 12'h8f7;
        src53 <= 12'h1e4;
        src54 <= 12'h74c;
        src55 <= 12'hee0;
        src56 <= 12'h234;
        src57 <= 12'hee1;
        src58 <= 12'h0;
        src59 <= 12'h264;
        src60 <= 12'hab3;
        src61 <= 12'h97a;
        src62 <= 12'hcf5;
        src63 <= 12'hf2b;
        src64 <= 12'h194;
        src65 <= 12'hfe8;
        src66 <= 12'h225;
        src67 <= 12'h7a0;
        src68 <= 12'haa7;
        src69 <= 12'h239;
        src70 <= 12'h6ee;
        src71 <= 12'hba;
        src72 <= 12'h613;
        src73 <= 12'h7c5;
        src74 <= 12'had3;
        src75 <= 12'ha88;
        src76 <= 12'hff1;
        src77 <= 12'hd0c;
        src78 <= 12'h912;
        src79 <= 12'h1ce;
        src80 <= 12'h828;
        src81 <= 12'h335;
        src82 <= 12'h23f;
        src83 <= 12'h80d;
        src84 <= 12'h444;
        src85 <= 12'h15a;
        src86 <= 12'hb5a;
        src87 <= 12'hfe5;
        src88 <= 12'haae;
        src89 <= 12'h671;
        src90 <= 12'hecf;
        src91 <= 12'h9ca;
        src92 <= 12'h8cc;
        src93 <= 12'h183;
        src94 <= 12'h6fd;
        src95 <= 12'h958;
        src96 <= 12'hbcf;
        src97 <= 12'h5a7;
        src98 <= 12'hd45;
        src99 <= 12'h507;
        src100 <= 12'hdd5;
        src101 <= 12'h5a5;
        src102 <= 12'ha00;
        src103 <= 12'h908;
        src104 <= 12'h68c;
        src105 <= 12'h771;
        src106 <= 12'h2ec;
        src107 <= 12'hb10;
        src108 <= 12'h346;
        src109 <= 12'h18e;
        src110 <= 12'hf6a;
        src111 <= 12'h70f;
        src112 <= 12'h55e;
        src113 <= 12'hc36;
        src114 <= 12'h133;
        src115 <= 12'h87;
        src116 <= 12'h771;
        src117 <= 12'h1f9;
        src118 <= 12'hba3;
        src119 <= 12'h4c5;
        src120 <= 12'hfd3;
        src121 <= 12'hda0;
        src122 <= 12'h80b;
        src123 <= 12'h855;
        src124 <= 12'h193;
        src125 <= 12'hcb3;
        src126 <= 12'h273;
        src127 <= 12'hfe5;
        exp <= 19'h3e36a;
        #1
        src0 <= 12'hcc4;
        src1 <= 12'h3a7;
        src2 <= 12'h468;
        src3 <= 12'h135;
        src4 <= 12'hf43;
        src5 <= 12'ha0c;
        src6 <= 12'h4e;
        src7 <= 12'h718;
        src8 <= 12'hac9;
        src9 <= 12'hfbd;
        src10 <= 12'hd4a;
        src11 <= 12'h55b;
        src12 <= 12'h8c6;
        src13 <= 12'h32f;
        src14 <= 12'h3d5;
        src15 <= 12'h892;
        src16 <= 12'h176;
        src17 <= 12'h726;
        src18 <= 12'h14f;
        src19 <= 12'h9c1;
        src20 <= 12'h477;
        src21 <= 12'hd44;
        src22 <= 12'hc41;
        src23 <= 12'hed7;
        src24 <= 12'ha93;
        src25 <= 12'hb2c;
        src26 <= 12'hcd9;
        src27 <= 12'hf93;
        src28 <= 12'h8dd;
        src29 <= 12'hdf6;
        src30 <= 12'h6f0;
        src31 <= 12'hf41;
        src32 <= 12'h3ac;
        src33 <= 12'hda7;
        src34 <= 12'h8fc;
        src35 <= 12'hac6;
        src36 <= 12'hfe9;
        src37 <= 12'he87;
        src38 <= 12'h316;
        src39 <= 12'hc24;
        src40 <= 12'h7f;
        src41 <= 12'h6b6;
        src42 <= 12'hfc8;
        src43 <= 12'hee3;
        src44 <= 12'he71;
        src45 <= 12'h216;
        src46 <= 12'h5b;
        src47 <= 12'hd09;
        src48 <= 12'he01;
        src49 <= 12'h6b;
        src50 <= 12'hf6b;
        src51 <= 12'h1e6;
        src52 <= 12'hdc3;
        src53 <= 12'h317;
        src54 <= 12'h1ca;
        src55 <= 12'h407;
        src56 <= 12'h378;
        src57 <= 12'hee7;
        src58 <= 12'ha3;
        src59 <= 12'h70f;
        src60 <= 12'h66b;
        src61 <= 12'haaa;
        src62 <= 12'hb9f;
        src63 <= 12'h56a;
        src64 <= 12'h4c3;
        src65 <= 12'hfb6;
        src66 <= 12'hb0a;
        src67 <= 12'h964;
        src68 <= 12'h3be;
        src69 <= 12'hc0b;
        src70 <= 12'h8aa;
        src71 <= 12'h20a;
        src72 <= 12'hd8;
        src73 <= 12'h4cc;
        src74 <= 12'ha76;
        src75 <= 12'hdcb;
        src76 <= 12'h5cd;
        src77 <= 12'hae3;
        src78 <= 12'h81c;
        src79 <= 12'h968;
        src80 <= 12'h523;
        src81 <= 12'hf20;
        src82 <= 12'he3a;
        src83 <= 12'h8;
        src84 <= 12'h4e4;
        src85 <= 12'h6a5;
        src86 <= 12'h4a7;
        src87 <= 12'hf1;
        src88 <= 12'h97;
        src89 <= 12'hd43;
        src90 <= 12'h284;
        src91 <= 12'ha38;
        src92 <= 12'ha35;
        src93 <= 12'hc1e;
        src94 <= 12'ha7c;
        src95 <= 12'hc53;
        src96 <= 12'h6b3;
        src97 <= 12'h7dd;
        src98 <= 12'h1c8;
        src99 <= 12'h8ce;
        src100 <= 12'hcb5;
        src101 <= 12'h43c;
        src102 <= 12'hee9;
        src103 <= 12'ha57;
        src104 <= 12'ha9b;
        src105 <= 12'h51b;
        src106 <= 12'hf08;
        src107 <= 12'hae2;
        src108 <= 12'h901;
        src109 <= 12'hc23;
        src110 <= 12'ha25;
        src111 <= 12'h246;
        src112 <= 12'hfc5;
        src113 <= 12'hbc4;
        src114 <= 12'hb08;
        src115 <= 12'hd95;
        src116 <= 12'h8d1;
        src117 <= 12'hf1a;
        src118 <= 12'hd24;
        src119 <= 12'hc34;
        src120 <= 12'h991;
        src121 <= 12'h5f;
        src122 <= 12'ha4c;
        src123 <= 12'h665;
        src124 <= 12'h4c2;
        src125 <= 12'hf07;
        src126 <= 12'hc07;
        src127 <= 12'h444;
        exp <= 19'h45692;
        #1
        src0 <= 12'h9d4;
        src1 <= 12'h836;
        src2 <= 12'h5e5;
        src3 <= 12'h885;
        src4 <= 12'h8f0;
        src5 <= 12'h447;
        src6 <= 12'h72d;
        src7 <= 12'hc36;
        src8 <= 12'hf05;
        src9 <= 12'h15a;
        src10 <= 12'h493;
        src11 <= 12'hb49;
        src12 <= 12'hd7d;
        src13 <= 12'h6ea;
        src14 <= 12'h66d;
        src15 <= 12'hb81;
        src16 <= 12'h546;
        src17 <= 12'heb6;
        src18 <= 12'hd71;
        src19 <= 12'hde2;
        src20 <= 12'hb62;
        src21 <= 12'h379;
        src22 <= 12'h30d;
        src23 <= 12'hbf7;
        src24 <= 12'h740;
        src25 <= 12'heeb;
        src26 <= 12'h66b;
        src27 <= 12'h63e;
        src28 <= 12'h19f;
        src29 <= 12'h6ef;
        src30 <= 12'h436;
        src31 <= 12'h326;
        src32 <= 12'h8e4;
        src33 <= 12'h92a;
        src34 <= 12'hf28;
        src35 <= 12'hb35;
        src36 <= 12'hc48;
        src37 <= 12'hb9a;
        src38 <= 12'hd32;
        src39 <= 12'hb12;
        src40 <= 12'hbb;
        src41 <= 12'hf00;
        src42 <= 12'h408;
        src43 <= 12'hf5f;
        src44 <= 12'h860;
        src45 <= 12'h262;
        src46 <= 12'h5da;
        src47 <= 12'h36a;
        src48 <= 12'hbb;
        src49 <= 12'h2c1;
        src50 <= 12'hc0;
        src51 <= 12'hb7e;
        src52 <= 12'h2;
        src53 <= 12'h5b1;
        src54 <= 12'h6cb;
        src55 <= 12'haba;
        src56 <= 12'h126;
        src57 <= 12'h19c;
        src58 <= 12'h358;
        src59 <= 12'h8a6;
        src60 <= 12'h4d3;
        src61 <= 12'hd0e;
        src62 <= 12'ha93;
        src63 <= 12'h734;
        src64 <= 12'h650;
        src65 <= 12'h252;
        src66 <= 12'h9d8;
        src67 <= 12'hc6;
        src68 <= 12'hba8;
        src69 <= 12'h8f4;
        src70 <= 12'h5f2;
        src71 <= 12'h1b6;
        src72 <= 12'h462;
        src73 <= 12'hc1;
        src74 <= 12'he61;
        src75 <= 12'h1e2;
        src76 <= 12'hd42;
        src77 <= 12'h66e;
        src78 <= 12'he22;
        src79 <= 12'he8b;
        src80 <= 12'hb2;
        src81 <= 12'h244;
        src82 <= 12'hfb7;
        src83 <= 12'h26e;
        src84 <= 12'hfa9;
        src85 <= 12'h2d0;
        src86 <= 12'h760;
        src87 <= 12'h967;
        src88 <= 12'hfd7;
        src89 <= 12'h776;
        src90 <= 12'ha32;
        src91 <= 12'h72c;
        src92 <= 12'h7f4;
        src93 <= 12'h95e;
        src94 <= 12'h231;
        src95 <= 12'hf89;
        src96 <= 12'h60d;
        src97 <= 12'hd21;
        src98 <= 12'h29d;
        src99 <= 12'hefe;
        src100 <= 12'h812;
        src101 <= 12'he50;
        src102 <= 12'hb78;
        src103 <= 12'hd15;
        src104 <= 12'hd5a;
        src105 <= 12'h59a;
        src106 <= 12'h4a5;
        src107 <= 12'h57c;
        src108 <= 12'hc2a;
        src109 <= 12'h68b;
        src110 <= 12'h81c;
        src111 <= 12'h87d;
        src112 <= 12'h689;
        src113 <= 12'hf92;
        src114 <= 12'hf37;
        src115 <= 12'hb49;
        src116 <= 12'hd2c;
        src117 <= 12'ha4e;
        src118 <= 12'h9fd;
        src119 <= 12'h825;
        src120 <= 12'h11d;
        src121 <= 12'hddc;
        src122 <= 12'he18;
        src123 <= 12'h641;
        src124 <= 12'h234;
        src125 <= 12'h8;
        src126 <= 12'h6d0;
        src127 <= 12'h850;
        exp <= 19'h410f6;
        #1
        src0 <= 12'hae0;
        src1 <= 12'h9d0;
        src2 <= 12'hd;
        src3 <= 12'he06;
        src4 <= 12'ha06;
        src5 <= 12'ha2e;
        src6 <= 12'h3ed;
        src7 <= 12'h3c4;
        src8 <= 12'hf34;
        src9 <= 12'h244;
        src10 <= 12'h53f;
        src11 <= 12'hca9;
        src12 <= 12'heda;
        src13 <= 12'h5de;
        src14 <= 12'h5a;
        src15 <= 12'h571;
        src16 <= 12'h9a;
        src17 <= 12'h134;
        src18 <= 12'hbcb;
        src19 <= 12'h6ef;
        src20 <= 12'hd2e;
        src21 <= 12'h6bf;
        src22 <= 12'h3b9;
        src23 <= 12'h970;
        src24 <= 12'hbff;
        src25 <= 12'h70;
        src26 <= 12'h8f1;
        src27 <= 12'h665;
        src28 <= 12'hb07;
        src29 <= 12'hf87;
        src30 <= 12'hcf0;
        src31 <= 12'h344;
        src32 <= 12'h468;
        src33 <= 12'h2b7;
        src34 <= 12'h903;
        src35 <= 12'h358;
        src36 <= 12'ha1b;
        src37 <= 12'hcd4;
        src38 <= 12'h164;
        src39 <= 12'h838;
        src40 <= 12'hd65;
        src41 <= 12'ha46;
        src42 <= 12'h5ad;
        src43 <= 12'h8fe;
        src44 <= 12'h120;
        src45 <= 12'h136;
        src46 <= 12'h4e0;
        src47 <= 12'h387;
        src48 <= 12'hf48;
        src49 <= 12'h643;
        src50 <= 12'h963;
        src51 <= 12'hbe0;
        src52 <= 12'h4dc;
        src53 <= 12'h1c1;
        src54 <= 12'h20b;
        src55 <= 12'hba2;
        src56 <= 12'he24;
        src57 <= 12'h97a;
        src58 <= 12'he23;
        src59 <= 12'he4f;
        src60 <= 12'h3e4;
        src61 <= 12'h244;
        src62 <= 12'h551;
        src63 <= 12'ha1d;
        src64 <= 12'hf1a;
        src65 <= 12'h371;
        src66 <= 12'h822;
        src67 <= 12'ha4b;
        src68 <= 12'h508;
        src69 <= 12'h347;
        src70 <= 12'ha35;
        src71 <= 12'h97a;
        src72 <= 12'h5ef;
        src73 <= 12'hd79;
        src74 <= 12'h3f6;
        src75 <= 12'h941;
        src76 <= 12'had1;
        src77 <= 12'h698;
        src78 <= 12'hb64;
        src79 <= 12'he35;
        src80 <= 12'h2df;
        src81 <= 12'h6f2;
        src82 <= 12'h322;
        src83 <= 12'h1fa;
        src84 <= 12'h29f;
        src85 <= 12'h5a5;
        src86 <= 12'h125;
        src87 <= 12'h3b1;
        src88 <= 12'h8ad;
        src89 <= 12'h6ca;
        src90 <= 12'hb69;
        src91 <= 12'haf7;
        src92 <= 12'h5e3;
        src93 <= 12'h5f4;
        src94 <= 12'h64a;
        src95 <= 12'h60a;
        src96 <= 12'hd70;
        src97 <= 12'h50;
        src98 <= 12'h4a0;
        src99 <= 12'hb8f;
        src100 <= 12'h1c6;
        src101 <= 12'h540;
        src102 <= 12'h362;
        src103 <= 12'hf57;
        src104 <= 12'hd51;
        src105 <= 12'hff1;
        src106 <= 12'hf96;
        src107 <= 12'h18e;
        src108 <= 12'h264;
        src109 <= 12'h787;
        src110 <= 12'h18e;
        src111 <= 12'h1bf;
        src112 <= 12'hcb7;
        src113 <= 12'hf66;
        src114 <= 12'h72c;
        src115 <= 12'h4c6;
        src116 <= 12'h668;
        src117 <= 12'h678;
        src118 <= 12'he34;
        src119 <= 12'ha7d;
        src120 <= 12'h87b;
        src121 <= 12'haec;
        src122 <= 12'hfc2;
        src123 <= 12'h477;
        src124 <= 12'h784;
        src125 <= 12'haba;
        src126 <= 12'h3a;
        src127 <= 12'h580;
        exp <= 19'h3cdaa;
        #1
        src0 <= 12'h6d0;
        src1 <= 12'h4e8;
        src2 <= 12'hf5;
        src3 <= 12'he05;
        src4 <= 12'h60d;
        src5 <= 12'h2b;
        src6 <= 12'h5ac;
        src7 <= 12'h7ad;
        src8 <= 12'h842;
        src9 <= 12'h63e;
        src10 <= 12'h6de;
        src11 <= 12'h49d;
        src12 <= 12'hed0;
        src13 <= 12'h6b3;
        src14 <= 12'h2ef;
        src15 <= 12'h980;
        src16 <= 12'hdc;
        src17 <= 12'hcb8;
        src18 <= 12'h70;
        src19 <= 12'haf8;
        src20 <= 12'h8a5;
        src21 <= 12'h12b;
        src22 <= 12'h59e;
        src23 <= 12'h1ab;
        src24 <= 12'heb0;
        src25 <= 12'h848;
        src26 <= 12'h1d5;
        src27 <= 12'h7a3;
        src28 <= 12'haaf;
        src29 <= 12'hf64;
        src30 <= 12'h538;
        src31 <= 12'h453;
        src32 <= 12'hc16;
        src33 <= 12'hc12;
        src34 <= 12'hc3;
        src35 <= 12'hfa2;
        src36 <= 12'hc36;
        src37 <= 12'h77b;
        src38 <= 12'hf67;
        src39 <= 12'h33c;
        src40 <= 12'hba9;
        src41 <= 12'hc45;
        src42 <= 12'h11f;
        src43 <= 12'hfc0;
        src44 <= 12'hf04;
        src45 <= 12'h55d;
        src46 <= 12'h64a;
        src47 <= 12'hc36;
        src48 <= 12'he76;
        src49 <= 12'h705;
        src50 <= 12'h57c;
        src51 <= 12'hc8;
        src52 <= 12'he7f;
        src53 <= 12'hd11;
        src54 <= 12'h332;
        src55 <= 12'he82;
        src56 <= 12'h80b;
        src57 <= 12'h739;
        src58 <= 12'h6e0;
        src59 <= 12'ha83;
        src60 <= 12'h9c5;
        src61 <= 12'habb;
        src62 <= 12'h61d;
        src63 <= 12'hb06;
        src64 <= 12'h824;
        src65 <= 12'hb1c;
        src66 <= 12'hbcf;
        src67 <= 12'h116;
        src68 <= 12'h9e6;
        src69 <= 12'h167;
        src70 <= 12'h48c;
        src71 <= 12'hc47;
        src72 <= 12'h2f5;
        src73 <= 12'h585;
        src74 <= 12'h87d;
        src75 <= 12'hdfc;
        src76 <= 12'h4c9;
        src77 <= 12'he9a;
        src78 <= 12'hd4b;
        src79 <= 12'hcfd;
        src80 <= 12'hba6;
        src81 <= 12'h8d5;
        src82 <= 12'hd3e;
        src83 <= 12'hf5c;
        src84 <= 12'h772;
        src85 <= 12'h8fb;
        src86 <= 12'h527;
        src87 <= 12'h51d;
        src88 <= 12'hf37;
        src89 <= 12'h9f6;
        src90 <= 12'hb66;
        src91 <= 12'h13;
        src92 <= 12'hf1;
        src93 <= 12'hf79;
        src94 <= 12'hd96;
        src95 <= 12'hd9;
        src96 <= 12'hf0d;
        src97 <= 12'h993;
        src98 <= 12'h3ff;
        src99 <= 12'h629;
        src100 <= 12'hd1e;
        src101 <= 12'h4ec;
        src102 <= 12'haae;
        src103 <= 12'hefd;
        src104 <= 12'h74a;
        src105 <= 12'h99d;
        src106 <= 12'h56e;
        src107 <= 12'hcb2;
        src108 <= 12'hf39;
        src109 <= 12'h6af;
        src110 <= 12'h201;
        src111 <= 12'h91f;
        src112 <= 12'h63f;
        src113 <= 12'hc71;
        src114 <= 12'h10f;
        src115 <= 12'h80a;
        src116 <= 12'hd6e;
        src117 <= 12'hec0;
        src118 <= 12'hbb2;
        src119 <= 12'h652;
        src120 <= 12'he32;
        src121 <= 12'ha27;
        src122 <= 12'h572;
        src123 <= 12'h966;
        src124 <= 12'h7f5;
        src125 <= 12'h933;
        src126 <= 12'hb81;
        src127 <= 12'h642;
        exp <= 19'h444fa;
        #1
        src0 <= 12'h4b9;
        src1 <= 12'h42c;
        src2 <= 12'h526;
        src3 <= 12'he5d;
        src4 <= 12'h4b9;
        src5 <= 12'h3c8;
        src6 <= 12'hd3d;
        src7 <= 12'h8a6;
        src8 <= 12'hb1e;
        src9 <= 12'h492;
        src10 <= 12'h365;
        src11 <= 12'h55f;
        src12 <= 12'hcfa;
        src13 <= 12'hb34;
        src14 <= 12'h2eb;
        src15 <= 12'h7;
        src16 <= 12'h20a;
        src17 <= 12'h3;
        src18 <= 12'h264;
        src19 <= 12'hda;
        src20 <= 12'h774;
        src21 <= 12'he42;
        src22 <= 12'hb87;
        src23 <= 12'h6d7;
        src24 <= 12'h5a5;
        src25 <= 12'hc20;
        src26 <= 12'h4c0;
        src27 <= 12'h23b;
        src28 <= 12'ha32;
        src29 <= 12'h6ba;
        src30 <= 12'hd64;
        src31 <= 12'h42d;
        src32 <= 12'hddd;
        src33 <= 12'hcff;
        src34 <= 12'h64a;
        src35 <= 12'h305;
        src36 <= 12'h648;
        src37 <= 12'ha65;
        src38 <= 12'h5d2;
        src39 <= 12'h151;
        src40 <= 12'hfd;
        src41 <= 12'hfa0;
        src42 <= 12'hee1;
        src43 <= 12'h89d;
        src44 <= 12'hbae;
        src45 <= 12'hdf;
        src46 <= 12'h739;
        src47 <= 12'hc39;
        src48 <= 12'hed4;
        src49 <= 12'hb2a;
        src50 <= 12'h546;
        src51 <= 12'h354;
        src52 <= 12'h793;
        src53 <= 12'h565;
        src54 <= 12'h96f;
        src55 <= 12'h6b1;
        src56 <= 12'h50e;
        src57 <= 12'h3e6;
        src58 <= 12'h938;
        src59 <= 12'h651;
        src60 <= 12'hc9d;
        src61 <= 12'hb18;
        src62 <= 12'h9f1;
        src63 <= 12'h6c9;
        src64 <= 12'h920;
        src65 <= 12'h8ad;
        src66 <= 12'h39b;
        src67 <= 12'hb7d;
        src68 <= 12'h74c;
        src69 <= 12'hbae;
        src70 <= 12'hdce;
        src71 <= 12'h3b7;
        src72 <= 12'hd7b;
        src73 <= 12'h7df;
        src74 <= 12'hd77;
        src75 <= 12'h1a3;
        src76 <= 12'hbf1;
        src77 <= 12'hda7;
        src78 <= 12'ha08;
        src79 <= 12'h65b;
        src80 <= 12'haa7;
        src81 <= 12'h23f;
        src82 <= 12'hfb9;
        src83 <= 12'he1f;
        src84 <= 12'h16f;
        src85 <= 12'hf35;
        src86 <= 12'h4ab;
        src87 <= 12'h14b;
        src88 <= 12'hea2;
        src89 <= 12'h2ab;
        src90 <= 12'h256;
        src91 <= 12'hc70;
        src92 <= 12'he52;
        src93 <= 12'h6ac;
        src94 <= 12'he9a;
        src95 <= 12'h8e3;
        src96 <= 12'h7ed;
        src97 <= 12'hbad;
        src98 <= 12'hbf6;
        src99 <= 12'h30e;
        src100 <= 12'hc5c;
        src101 <= 12'haab;
        src102 <= 12'ha9a;
        src103 <= 12'h6b6;
        src104 <= 12'h647;
        src105 <= 12'hb04;
        src106 <= 12'h50c;
        src107 <= 12'h9ef;
        src108 <= 12'h10a;
        src109 <= 12'h25b;
        src110 <= 12'h459;
        src111 <= 12'h100;
        src112 <= 12'h24f;
        src113 <= 12'h5a;
        src114 <= 12'hd2b;
        src115 <= 12'h9a9;
        src116 <= 12'h7a2;
        src117 <= 12'h944;
        src118 <= 12'h1ff;
        src119 <= 12'h821;
        src120 <= 12'h7fc;
        src121 <= 12'h729;
        src122 <= 12'h3ce;
        src123 <= 12'hccc;
        src124 <= 12'h287;
        src125 <= 12'h972;
        src126 <= 12'h74a;
        src127 <= 12'h57a;
        exp <= 19'h3de5e;
        #1
        src0 <= 12'h52d;
        src1 <= 12'hcd3;
        src2 <= 12'h43d;
        src3 <= 12'hfdd;
        src4 <= 12'h513;
        src5 <= 12'hc22;
        src6 <= 12'h835;
        src7 <= 12'h9a6;
        src8 <= 12'h406;
        src9 <= 12'hfbb;
        src10 <= 12'hfd7;
        src11 <= 12'he44;
        src12 <= 12'hb7;
        src13 <= 12'hcba;
        src14 <= 12'ha38;
        src15 <= 12'h6b0;
        src16 <= 12'h601;
        src17 <= 12'hcc0;
        src18 <= 12'h780;
        src19 <= 12'h6e7;
        src20 <= 12'h706;
        src21 <= 12'hc10;
        src22 <= 12'h872;
        src23 <= 12'h561;
        src24 <= 12'hf48;
        src25 <= 12'h874;
        src26 <= 12'h476;
        src27 <= 12'h3cc;
        src28 <= 12'h806;
        src29 <= 12'hc8d;
        src30 <= 12'h5d5;
        src31 <= 12'h4c7;
        src32 <= 12'h874;
        src33 <= 12'hdf1;
        src34 <= 12'hb5b;
        src35 <= 12'h539;
        src36 <= 12'h91f;
        src37 <= 12'h4f3;
        src38 <= 12'h927;
        src39 <= 12'h263;
        src40 <= 12'he3b;
        src41 <= 12'h6d7;
        src42 <= 12'h63f;
        src43 <= 12'h5ed;
        src44 <= 12'h30b;
        src45 <= 12'h7c6;
        src46 <= 12'ha65;
        src47 <= 12'h6d1;
        src48 <= 12'h928;
        src49 <= 12'h65e;
        src50 <= 12'h65a;
        src51 <= 12'h9dc;
        src52 <= 12'hb0e;
        src53 <= 12'h376;
        src54 <= 12'h651;
        src55 <= 12'h48d;
        src56 <= 12'ha5e;
        src57 <= 12'h6d3;
        src58 <= 12'h9af;
        src59 <= 12'hfc2;
        src60 <= 12'h9da;
        src61 <= 12'hbc5;
        src62 <= 12'h1a5;
        src63 <= 12'h316;
        src64 <= 12'h7db;
        src65 <= 12'h127;
        src66 <= 12'hb6;
        src67 <= 12'h1bf;
        src68 <= 12'hfd8;
        src69 <= 12'h12a;
        src70 <= 12'h8df;
        src71 <= 12'he6f;
        src72 <= 12'hf40;
        src73 <= 12'hf82;
        src74 <= 12'ha1d;
        src75 <= 12'heb9;
        src76 <= 12'hfcd;
        src77 <= 12'h284;
        src78 <= 12'h945;
        src79 <= 12'hf11;
        src80 <= 12'hc09;
        src81 <= 12'h992;
        src82 <= 12'h719;
        src83 <= 12'h59b;
        src84 <= 12'hf86;
        src85 <= 12'hcfd;
        src86 <= 12'h8c7;
        src87 <= 12'hb95;
        src88 <= 12'h1e;
        src89 <= 12'hd17;
        src90 <= 12'hc56;
        src91 <= 12'h189;
        src92 <= 12'h376;
        src93 <= 12'hba;
        src94 <= 12'he9e;
        src95 <= 12'h3d;
        src96 <= 12'hf83;
        src97 <= 12'h829;
        src98 <= 12'h613;
        src99 <= 12'ha47;
        src100 <= 12'h87c;
        src101 <= 12'hfb8;
        src102 <= 12'hf53;
        src103 <= 12'h854;
        src104 <= 12'he67;
        src105 <= 12'hd03;
        src106 <= 12'h69d;
        src107 <= 12'h5a2;
        src108 <= 12'h2c8;
        src109 <= 12'h9bd;
        src110 <= 12'h1b4;
        src111 <= 12'h3b5;
        src112 <= 12'h137;
        src113 <= 12'h14a;
        src114 <= 12'hea6;
        src115 <= 12'hbd8;
        src116 <= 12'hb69;
        src117 <= 12'h595;
        src118 <= 12'ha45;
        src119 <= 12'h54f;
        src120 <= 12'hc05;
        src121 <= 12'hcb7;
        src122 <= 12'hd5c;
        src123 <= 12'h1db;
        src124 <= 12'h6a6;
        src125 <= 12'h9b;
        src126 <= 12'h375;
        src127 <= 12'h104;
        exp <= 19'h4309a;
        #1
        src0 <= 12'h8d7;
        src1 <= 12'h21a;
        src2 <= 12'h328;
        src3 <= 12'ha81;
        src4 <= 12'h5ab;
        src5 <= 12'hdda;
        src6 <= 12'h7aa;
        src7 <= 12'h393;
        src8 <= 12'hfbc;
        src9 <= 12'hddd;
        src10 <= 12'h79e;
        src11 <= 12'hbd9;
        src12 <= 12'h65e;
        src13 <= 12'hc78;
        src14 <= 12'haba;
        src15 <= 12'h18a;
        src16 <= 12'h131;
        src17 <= 12'hcf4;
        src18 <= 12'hb04;
        src19 <= 12'hd74;
        src20 <= 12'h4f4;
        src21 <= 12'h907;
        src22 <= 12'h25f;
        src23 <= 12'hd80;
        src24 <= 12'h290;
        src25 <= 12'h582;
        src26 <= 12'hd83;
        src27 <= 12'hccc;
        src28 <= 12'h5eb;
        src29 <= 12'h62b;
        src30 <= 12'ha0e;
        src31 <= 12'h7d0;
        src32 <= 12'h4b1;
        src33 <= 12'had9;
        src34 <= 12'h9e5;
        src35 <= 12'h81d;
        src36 <= 12'h284;
        src37 <= 12'h18c;
        src38 <= 12'h3c6;
        src39 <= 12'hcb6;
        src40 <= 12'h674;
        src41 <= 12'h181;
        src42 <= 12'h29a;
        src43 <= 12'h88;
        src44 <= 12'h412;
        src45 <= 12'h66c;
        src46 <= 12'h5c2;
        src47 <= 12'h27e;
        src48 <= 12'h128;
        src49 <= 12'h225;
        src50 <= 12'h25;
        src51 <= 12'h592;
        src52 <= 12'hd77;
        src53 <= 12'hce9;
        src54 <= 12'hf9c;
        src55 <= 12'h794;
        src56 <= 12'hcb6;
        src57 <= 12'h2f1;
        src58 <= 12'hcc0;
        src59 <= 12'hc74;
        src60 <= 12'h37f;
        src61 <= 12'h83;
        src62 <= 12'h242;
        src63 <= 12'hee3;
        src64 <= 12'hdfd;
        src65 <= 12'h45c;
        src66 <= 12'h76c;
        src67 <= 12'ha9;
        src68 <= 12'hdc9;
        src69 <= 12'h647;
        src70 <= 12'h2b7;
        src71 <= 12'h4d9;
        src72 <= 12'he17;
        src73 <= 12'h665;
        src74 <= 12'h5a8;
        src75 <= 12'h9e5;
        src76 <= 12'h528;
        src77 <= 12'h4c7;
        src78 <= 12'hec8;
        src79 <= 12'hcd6;
        src80 <= 12'hd9;
        src81 <= 12'h80;
        src82 <= 12'h4d1;
        src83 <= 12'h10f;
        src84 <= 12'h5dd;
        src85 <= 12'h3cb;
        src86 <= 12'h7f;
        src87 <= 12'h892;
        src88 <= 12'h9b2;
        src89 <= 12'h738;
        src90 <= 12'h611;
        src91 <= 12'h189;
        src92 <= 12'hf42;
        src93 <= 12'he98;
        src94 <= 12'hcb1;
        src95 <= 12'hf11;
        src96 <= 12'h515;
        src97 <= 12'ha97;
        src98 <= 12'h145;
        src99 <= 12'h587;
        src100 <= 12'hc2d;
        src101 <= 12'h42f;
        src102 <= 12'h327;
        src103 <= 12'hb5d;
        src104 <= 12'h237;
        src105 <= 12'h73c;
        src106 <= 12'h71c;
        src107 <= 12'h55;
        src108 <= 12'hbb3;
        src109 <= 12'h149;
        src110 <= 12'h5d6;
        src111 <= 12'hbae;
        src112 <= 12'h890;
        src113 <= 12'h3f1;
        src114 <= 12'h852;
        src115 <= 12'h3e3;
        src116 <= 12'h45e;
        src117 <= 12'h78b;
        src118 <= 12'h98e;
        src119 <= 12'h190;
        src120 <= 12'hc0c;
        src121 <= 12'hece;
        src122 <= 12'h54c;
        src123 <= 12'hc1c;
        src124 <= 12'ha64;
        src125 <= 12'ha6d;
        src126 <= 12'h4ba;
        src127 <= 12'hc1b;
        exp <= 19'h3aaec;
        #1
        src0 <= 12'h833;
        src1 <= 12'h5a4;
        src2 <= 12'hea1;
        src3 <= 12'h15b;
        src4 <= 12'hb80;
        src5 <= 12'ha9c;
        src6 <= 12'hfc6;
        src7 <= 12'he4c;
        src8 <= 12'hc3d;
        src9 <= 12'h2f8;
        src10 <= 12'hbc;
        src11 <= 12'hfda;
        src12 <= 12'he85;
        src13 <= 12'hdca;
        src14 <= 12'h2b9;
        src15 <= 12'h63b;
        src16 <= 12'h8cd;
        src17 <= 12'h8db;
        src18 <= 12'h887;
        src19 <= 12'hf49;
        src20 <= 12'heb2;
        src21 <= 12'h200;
        src22 <= 12'h6c0;
        src23 <= 12'hb44;
        src24 <= 12'h1ad;
        src25 <= 12'h9ae;
        src26 <= 12'hc81;
        src27 <= 12'h771;
        src28 <= 12'h651;
        src29 <= 12'hd2e;
        src30 <= 12'h7a1;
        src31 <= 12'h360;
        src32 <= 12'h2a3;
        src33 <= 12'hbad;
        src34 <= 12'hde9;
        src35 <= 12'hd69;
        src36 <= 12'h6be;
        src37 <= 12'h823;
        src38 <= 12'hcf1;
        src39 <= 12'h786;
        src40 <= 12'h29e;
        src41 <= 12'hc2a;
        src42 <= 12'h8e1;
        src43 <= 12'h84c;
        src44 <= 12'hb16;
        src45 <= 12'h256;
        src46 <= 12'h4bd;
        src47 <= 12'hd69;
        src48 <= 12'haec;
        src49 <= 12'h7ee;
        src50 <= 12'hdf3;
        src51 <= 12'h4c;
        src52 <= 12'h31a;
        src53 <= 12'h831;
        src54 <= 12'hec;
        src55 <= 12'hd8f;
        src56 <= 12'ha45;
        src57 <= 12'h669;
        src58 <= 12'hef4;
        src59 <= 12'h57a;
        src60 <= 12'h53c;
        src61 <= 12'h1c3;
        src62 <= 12'h403;
        src63 <= 12'h411;
        src64 <= 12'he10;
        src65 <= 12'h8a4;
        src66 <= 12'h5ce;
        src67 <= 12'hb7;
        src68 <= 12'h639;
        src69 <= 12'h16e;
        src70 <= 12'h2df;
        src71 <= 12'h6a;
        src72 <= 12'h3;
        src73 <= 12'hde6;
        src74 <= 12'h1c1;
        src75 <= 12'h29;
        src76 <= 12'h32d;
        src77 <= 12'h67d;
        src78 <= 12'ha46;
        src79 <= 12'hee9;
        src80 <= 12'hf94;
        src81 <= 12'he52;
        src82 <= 12'ha3d;
        src83 <= 12'h8a1;
        src84 <= 12'hd2e;
        src85 <= 12'he59;
        src86 <= 12'hcc2;
        src87 <= 12'h37;
        src88 <= 12'h310;
        src89 <= 12'h3dd;
        src90 <= 12'he54;
        src91 <= 12'h775;
        src92 <= 12'h48d;
        src93 <= 12'h423;
        src94 <= 12'h2d;
        src95 <= 12'h300;
        src96 <= 12'h3d4;
        src97 <= 12'hbe8;
        src98 <= 12'ha95;
        src99 <= 12'h851;
        src100 <= 12'hf26;
        src101 <= 12'hc90;
        src102 <= 12'h149;
        src103 <= 12'h910;
        src104 <= 12'hfe8;
        src105 <= 12'h8a7;
        src106 <= 12'hc5d;
        src107 <= 12'h194;
        src108 <= 12'h765;
        src109 <= 12'he90;
        src110 <= 12'h53f;
        src111 <= 12'he10;
        src112 <= 12'hae;
        src113 <= 12'ha67;
        src114 <= 12'hf7d;
        src115 <= 12'hdb0;
        src116 <= 12'h79b;
        src117 <= 12'h78;
        src118 <= 12'hfa6;
        src119 <= 12'hb87;
        src120 <= 12'hfb5;
        src121 <= 12'h557;
        src122 <= 12'h9af;
        src123 <= 12'hc78;
        src124 <= 12'hf8d;
        src125 <= 12'h191;
        src126 <= 12'h794;
        src127 <= 12'h65e;
        exp <= 19'h4277f;
        #1
        src0 <= 12'hd92;
        src1 <= 12'h427;
        src2 <= 12'hf0f;
        src3 <= 12'hbc9;
        src4 <= 12'he75;
        src5 <= 12'h5e5;
        src6 <= 12'h676;
        src7 <= 12'hb4d;
        src8 <= 12'h1e2;
        src9 <= 12'h4;
        src10 <= 12'hee3;
        src11 <= 12'h4d8;
        src12 <= 12'h310;
        src13 <= 12'hc8a;
        src14 <= 12'h243;
        src15 <= 12'hbac;
        src16 <= 12'hc2e;
        src17 <= 12'h704;
        src18 <= 12'h34;
        src19 <= 12'h24b;
        src20 <= 12'h7ec;
        src21 <= 12'h8c4;
        src22 <= 12'h502;
        src23 <= 12'h248;
        src24 <= 12'h161;
        src25 <= 12'hbbf;
        src26 <= 12'h9e3;
        src27 <= 12'h888;
        src28 <= 12'h4b9;
        src29 <= 12'h9db;
        src30 <= 12'ha5f;
        src31 <= 12'h474;
        src32 <= 12'h77c;
        src33 <= 12'h74e;
        src34 <= 12'hfc0;
        src35 <= 12'hc6b;
        src36 <= 12'had8;
        src37 <= 12'h312;
        src38 <= 12'h858;
        src39 <= 12'hea1;
        src40 <= 12'h9b;
        src41 <= 12'hd79;
        src42 <= 12'hf80;
        src43 <= 12'h6e2;
        src44 <= 12'heef;
        src45 <= 12'hdf;
        src46 <= 12'ha7e;
        src47 <= 12'h38e;
        src48 <= 12'hed4;
        src49 <= 12'h812;
        src50 <= 12'hde5;
        src51 <= 12'ha12;
        src52 <= 12'h7d6;
        src53 <= 12'h185;
        src54 <= 12'h7d5;
        src55 <= 12'hd9f;
        src56 <= 12'h725;
        src57 <= 12'h841;
        src58 <= 12'hc7c;
        src59 <= 12'h131;
        src60 <= 12'h40e;
        src61 <= 12'hd97;
        src62 <= 12'hdb6;
        src63 <= 12'hfd1;
        src64 <= 12'h9ec;
        src65 <= 12'h4bb;
        src66 <= 12'h5bd;
        src67 <= 12'h73a;
        src68 <= 12'hd33;
        src69 <= 12'h54a;
        src70 <= 12'h764;
        src71 <= 12'hb6d;
        src72 <= 12'hc61;
        src73 <= 12'h2f1;
        src74 <= 12'hbd;
        src75 <= 12'h411;
        src76 <= 12'hf77;
        src77 <= 12'h94b;
        src78 <= 12'h30b;
        src79 <= 12'ha89;
        src80 <= 12'ha5b;
        src81 <= 12'h412;
        src82 <= 12'hfa4;
        src83 <= 12'ha83;
        src84 <= 12'h3aa;
        src85 <= 12'h1e5;
        src86 <= 12'hc64;
        src87 <= 12'h9d4;
        src88 <= 12'hc10;
        src89 <= 12'h477;
        src90 <= 12'haa0;
        src91 <= 12'h7c8;
        src92 <= 12'h120;
        src93 <= 12'h5de;
        src94 <= 12'ha67;
        src95 <= 12'h8e0;
        src96 <= 12'h390;
        src97 <= 12'h70e;
        src98 <= 12'h2d7;
        src99 <= 12'h3ae;
        src100 <= 12'ha9f;
        src101 <= 12'h20d;
        src102 <= 12'hd78;
        src103 <= 12'h3ad;
        src104 <= 12'he2b;
        src105 <= 12'h6fb;
        src106 <= 12'h6c5;
        src107 <= 12'h131;
        src108 <= 12'h5b0;
        src109 <= 12'h4b3;
        src110 <= 12'h9b5;
        src111 <= 12'h16;
        src112 <= 12'h122;
        src113 <= 12'h1dc;
        src114 <= 12'hd0d;
        src115 <= 12'h5cb;
        src116 <= 12'h9c0;
        src117 <= 12'hfb;
        src118 <= 12'h62b;
        src119 <= 12'h2cc;
        src120 <= 12'hdf0;
        src121 <= 12'hbf7;
        src122 <= 12'hb4;
        src123 <= 12'h636;
        src124 <= 12'h1ce;
        src125 <= 12'hfad;
        src126 <= 12'he33;
        src127 <= 12'ha85;
        exp <= 19'h3ee43;
        #1
        src0 <= 12'he04;
        src1 <= 12'h6fe;
        src2 <= 12'ha95;
        src3 <= 12'had4;
        src4 <= 12'h835;
        src5 <= 12'h628;
        src6 <= 12'h8aa;
        src7 <= 12'h593;
        src8 <= 12'h7d5;
        src9 <= 12'he68;
        src10 <= 12'hcc4;
        src11 <= 12'he9d;
        src12 <= 12'h3dc;
        src13 <= 12'hc;
        src14 <= 12'hbb6;
        src15 <= 12'h287;
        src16 <= 12'h72;
        src17 <= 12'h9f0;
        src18 <= 12'hb28;
        src19 <= 12'hf26;
        src20 <= 12'hcb6;
        src21 <= 12'hfcd;
        src22 <= 12'h18c;
        src23 <= 12'hcf7;
        src24 <= 12'hbb6;
        src25 <= 12'h1ae;
        src26 <= 12'hc9c;
        src27 <= 12'h1a8;
        src28 <= 12'hb1d;
        src29 <= 12'h2e9;
        src30 <= 12'hd01;
        src31 <= 12'h2e3;
        src32 <= 12'h164;
        src33 <= 12'h415;
        src34 <= 12'haaf;
        src35 <= 12'h92a;
        src36 <= 12'h109;
        src37 <= 12'ha9;
        src38 <= 12'h9b;
        src39 <= 12'h613;
        src40 <= 12'h8c3;
        src41 <= 12'h929;
        src42 <= 12'h2f7;
        src43 <= 12'h73e;
        src44 <= 12'hb03;
        src45 <= 12'hcb8;
        src46 <= 12'hb59;
        src47 <= 12'hffb;
        src48 <= 12'hc75;
        src49 <= 12'h9f8;
        src50 <= 12'h869;
        src51 <= 12'h21e;
        src52 <= 12'h8b2;
        src53 <= 12'h48a;
        src54 <= 12'h8e;
        src55 <= 12'h486;
        src56 <= 12'hc03;
        src57 <= 12'he58;
        src58 <= 12'h95d;
        src59 <= 12'he1e;
        src60 <= 12'haa7;
        src61 <= 12'he2b;
        src62 <= 12'he5f;
        src63 <= 12'h4a;
        src64 <= 12'h8a6;
        src65 <= 12'h17b;
        src66 <= 12'h103;
        src67 <= 12'h307;
        src68 <= 12'hf92;
        src69 <= 12'h42f;
        src70 <= 12'hccc;
        src71 <= 12'h6dc;
        src72 <= 12'hb9b;
        src73 <= 12'h86b;
        src74 <= 12'h342;
        src75 <= 12'h6be;
        src76 <= 12'hc58;
        src77 <= 12'hfba;
        src78 <= 12'h721;
        src79 <= 12'h4cb;
        src80 <= 12'hc;
        src81 <= 12'h7d7;
        src82 <= 12'h1ea;
        src83 <= 12'h5cd;
        src84 <= 12'h5eb;
        src85 <= 12'h9c2;
        src86 <= 12'h6ef;
        src87 <= 12'h3f9;
        src88 <= 12'hc54;
        src89 <= 12'h60c;
        src90 <= 12'h2a3;
        src91 <= 12'hfae;
        src92 <= 12'h88;
        src93 <= 12'hce;
        src94 <= 12'h480;
        src95 <= 12'h119;
        src96 <= 12'h89d;
        src97 <= 12'h9e2;
        src98 <= 12'he7e;
        src99 <= 12'he72;
        src100 <= 12'h5a3;
        src101 <= 12'h3ab;
        src102 <= 12'h6f4;
        src103 <= 12'h15a;
        src104 <= 12'h5e7;
        src105 <= 12'h557;
        src106 <= 12'he47;
        src107 <= 12'hca9;
        src108 <= 12'h64;
        src109 <= 12'h402;
        src110 <= 12'h88f;
        src111 <= 12'hfae;
        src112 <= 12'h2c8;
        src113 <= 12'h892;
        src114 <= 12'he2f;
        src115 <= 12'h348;
        src116 <= 12'hc7c;
        src117 <= 12'he95;
        src118 <= 12'hde4;
        src119 <= 12'hca8;
        src120 <= 12'hfeb;
        src121 <= 12'h105;
        src122 <= 12'hf25;
        src123 <= 12'h230;
        src124 <= 12'h277;
        src125 <= 12'h7e2;
        src126 <= 12'hb52;
        src127 <= 12'ha51;
        exp <= 19'h3fb79;
        #1
        src0 <= 12'hba3;
        src1 <= 12'hbc5;
        src2 <= 12'hb0;
        src3 <= 12'h8b2;
        src4 <= 12'hb17;
        src5 <= 12'hdfe;
        src6 <= 12'h72d;
        src7 <= 12'h957;
        src8 <= 12'h12f;
        src9 <= 12'h939;
        src10 <= 12'h9df;
        src11 <= 12'hfe;
        src12 <= 12'h644;
        src13 <= 12'h9ab;
        src14 <= 12'h566;
        src15 <= 12'hd90;
        src16 <= 12'ha38;
        src17 <= 12'h846;
        src18 <= 12'hbda;
        src19 <= 12'h47;
        src20 <= 12'h23d;
        src21 <= 12'hfd;
        src22 <= 12'hc0f;
        src23 <= 12'h660;
        src24 <= 12'h57e;
        src25 <= 12'hcb1;
        src26 <= 12'h623;
        src27 <= 12'hbfe;
        src28 <= 12'h420;
        src29 <= 12'hc30;
        src30 <= 12'h67b;
        src31 <= 12'h36f;
        src32 <= 12'h56d;
        src33 <= 12'h224;
        src34 <= 12'h699;
        src35 <= 12'hfa0;
        src36 <= 12'hf7c;
        src37 <= 12'h621;
        src38 <= 12'h333;
        src39 <= 12'hd8f;
        src40 <= 12'hf21;
        src41 <= 12'ha59;
        src42 <= 12'h414;
        src43 <= 12'hd6d;
        src44 <= 12'h353;
        src45 <= 12'h45;
        src46 <= 12'h9a9;
        src47 <= 12'h75e;
        src48 <= 12'h1e8;
        src49 <= 12'hca;
        src50 <= 12'h8ad;
        src51 <= 12'h36d;
        src52 <= 12'hfb8;
        src53 <= 12'h50c;
        src54 <= 12'hd9b;
        src55 <= 12'h855;
        src56 <= 12'h9af;
        src57 <= 12'ha33;
        src58 <= 12'h2a5;
        src59 <= 12'he03;
        src60 <= 12'h3af;
        src61 <= 12'hbf;
        src62 <= 12'hbc9;
        src63 <= 12'h5a3;
        src64 <= 12'h1dc;
        src65 <= 12'h75;
        src66 <= 12'h836;
        src67 <= 12'hf30;
        src68 <= 12'hf66;
        src69 <= 12'h874;
        src70 <= 12'h469;
        src71 <= 12'h94d;
        src72 <= 12'h9a1;
        src73 <= 12'he32;
        src74 <= 12'haf8;
        src75 <= 12'h5a4;
        src76 <= 12'hec;
        src77 <= 12'h707;
        src78 <= 12'h972;
        src79 <= 12'hf11;
        src80 <= 12'ha63;
        src81 <= 12'h7ac;
        src82 <= 12'he87;
        src83 <= 12'h7b8;
        src84 <= 12'h542;
        src85 <= 12'hf3b;
        src86 <= 12'h16c;
        src87 <= 12'hc1;
        src88 <= 12'h330;
        src89 <= 12'hea4;
        src90 <= 12'h12f;
        src91 <= 12'h240;
        src92 <= 12'hfd3;
        src93 <= 12'hb8c;
        src94 <= 12'h1e5;
        src95 <= 12'h6;
        src96 <= 12'hd34;
        src97 <= 12'hc2e;
        src98 <= 12'h5a8;
        src99 <= 12'hb38;
        src100 <= 12'h817;
        src101 <= 12'hd08;
        src102 <= 12'ha95;
        src103 <= 12'h95;
        src104 <= 12'h709;
        src105 <= 12'hf07;
        src106 <= 12'h22b;
        src107 <= 12'hc3a;
        src108 <= 12'h19f;
        src109 <= 12'h253;
        src110 <= 12'hb1;
        src111 <= 12'ha56;
        src112 <= 12'h22c;
        src113 <= 12'h121;
        src114 <= 12'ha48;
        src115 <= 12'h788;
        src116 <= 12'hf18;
        src117 <= 12'h997;
        src118 <= 12'h3c8;
        src119 <= 12'h564;
        src120 <= 12'hed5;
        src121 <= 12'hcc3;
        src122 <= 12'hb2f;
        src123 <= 12'hfc3;
        src124 <= 12'h1a8;
        src125 <= 12'hd;
        src126 <= 12'h95b;
        src127 <= 12'h34;
        exp <= 19'h3dd76;
        #1
        src0 <= 12'h405;
        src1 <= 12'h631;
        src2 <= 12'h40f;
        src3 <= 12'h3f2;
        src4 <= 12'h80e;
        src5 <= 12'h8c5;
        src6 <= 12'h15a;
        src7 <= 12'hb3c;
        src8 <= 12'hbf;
        src9 <= 12'h17f;
        src10 <= 12'he0d;
        src11 <= 12'hfb7;
        src12 <= 12'hbe0;
        src13 <= 12'h57b;
        src14 <= 12'h34f;
        src15 <= 12'hade;
        src16 <= 12'h75d;
        src17 <= 12'h454;
        src18 <= 12'h24a;
        src19 <= 12'h9f6;
        src20 <= 12'h9d8;
        src21 <= 12'h7ae;
        src22 <= 12'h553;
        src23 <= 12'h6d0;
        src24 <= 12'h52d;
        src25 <= 12'ha58;
        src26 <= 12'h8ea;
        src27 <= 12'h576;
        src28 <= 12'ha5b;
        src29 <= 12'h213;
        src30 <= 12'h155;
        src31 <= 12'h13b;
        src32 <= 12'h224;
        src33 <= 12'h33c;
        src34 <= 12'h1ee;
        src35 <= 12'hc48;
        src36 <= 12'h106;
        src37 <= 12'hade;
        src38 <= 12'h33a;
        src39 <= 12'h231;
        src40 <= 12'hc4b;
        src41 <= 12'h239;
        src42 <= 12'h5f0;
        src43 <= 12'h673;
        src44 <= 12'h529;
        src45 <= 12'hd69;
        src46 <= 12'h4f6;
        src47 <= 12'h823;
        src48 <= 12'h3bc;
        src49 <= 12'h8d6;
        src50 <= 12'he2d;
        src51 <= 12'h7bc;
        src52 <= 12'h201;
        src53 <= 12'h270;
        src54 <= 12'h599;
        src55 <= 12'h11;
        src56 <= 12'h78a;
        src57 <= 12'h76e;
        src58 <= 12'h537;
        src59 <= 12'h415;
        src60 <= 12'h984;
        src61 <= 12'ha1c;
        src62 <= 12'h9b0;
        src63 <= 12'hd48;
        src64 <= 12'hb53;
        src65 <= 12'hc0d;
        src66 <= 12'h271;
        src67 <= 12'hbdb;
        src68 <= 12'h1b7;
        src69 <= 12'hf12;
        src70 <= 12'hee;
        src71 <= 12'hcf0;
        src72 <= 12'haf2;
        src73 <= 12'h815;
        src74 <= 12'h6ba;
        src75 <= 12'h464;
        src76 <= 12'h65a;
        src77 <= 12'h6fe;
        src78 <= 12'h5fb;
        src79 <= 12'hde4;
        src80 <= 12'ha7f;
        src81 <= 12'hdbe;
        src82 <= 12'h8f2;
        src83 <= 12'h209;
        src84 <= 12'h52;
        src85 <= 12'h4ea;
        src86 <= 12'h84e;
        src87 <= 12'h2f4;
        src88 <= 12'h306;
        src89 <= 12'hee4;
        src90 <= 12'hd52;
        src91 <= 12'hb1d;
        src92 <= 12'h92f;
        src93 <= 12'he70;
        src94 <= 12'h44;
        src95 <= 12'h17e;
        src96 <= 12'hac6;
        src97 <= 12'hdc7;
        src98 <= 12'h6ee;
        src99 <= 12'h697;
        src100 <= 12'h395;
        src101 <= 12'he0d;
        src102 <= 12'h561;
        src103 <= 12'h19f;
        src104 <= 12'hba6;
        src105 <= 12'h6f9;
        src106 <= 12'h535;
        src107 <= 12'h5c7;
        src108 <= 12'hfa6;
        src109 <= 12'hd2a;
        src110 <= 12'h1a7;
        src111 <= 12'h4dd;
        src112 <= 12'hc56;
        src113 <= 12'h5d1;
        src114 <= 12'hdd3;
        src115 <= 12'h1a8;
        src116 <= 12'h8cd;
        src117 <= 12'hd03;
        src118 <= 12'hcb7;
        src119 <= 12'h477;
        src120 <= 12'h97f;
        src121 <= 12'h4af;
        src122 <= 12'hbfb;
        src123 <= 12'h6af;
        src124 <= 12'h2ee;
        src125 <= 12'h364;
        src126 <= 12'ha41;
        src127 <= 12'h73d;
        exp <= 19'h39c9a;
        #1
        src0 <= 12'h193;
        src1 <= 12'h9e4;
        src2 <= 12'h163;
        src3 <= 12'h9ee;
        src4 <= 12'h1fc;
        src5 <= 12'h88e;
        src6 <= 12'h668;
        src7 <= 12'h2f9;
        src8 <= 12'ha50;
        src9 <= 12'h160;
        src10 <= 12'h5bf;
        src11 <= 12'h31e;
        src12 <= 12'hdc0;
        src13 <= 12'hae4;
        src14 <= 12'h16c;
        src15 <= 12'hdee;
        src16 <= 12'h21b;
        src17 <= 12'hab3;
        src18 <= 12'h9bf;
        src19 <= 12'h95c;
        src20 <= 12'h7f3;
        src21 <= 12'h1e9;
        src22 <= 12'h6fd;
        src23 <= 12'he01;
        src24 <= 12'h22a;
        src25 <= 12'h675;
        src26 <= 12'heac;
        src27 <= 12'h477;
        src28 <= 12'h148;
        src29 <= 12'hfe7;
        src30 <= 12'h1e6;
        src31 <= 12'hea3;
        src32 <= 12'h947;
        src33 <= 12'h50;
        src34 <= 12'h2b9;
        src35 <= 12'hccc;
        src36 <= 12'he76;
        src37 <= 12'ha27;
        src38 <= 12'h1e1;
        src39 <= 12'hd07;
        src40 <= 12'h3c7;
        src41 <= 12'h51f;
        src42 <= 12'h414;
        src43 <= 12'h677;
        src44 <= 12'ha58;
        src45 <= 12'hcf9;
        src46 <= 12'h1d3;
        src47 <= 12'h61e;
        src48 <= 12'hb2b;
        src49 <= 12'hb32;
        src50 <= 12'he99;
        src51 <= 12'h22;
        src52 <= 12'h29c;
        src53 <= 12'hc5b;
        src54 <= 12'hd2f;
        src55 <= 12'h241;
        src56 <= 12'hd84;
        src57 <= 12'h916;
        src58 <= 12'h5a9;
        src59 <= 12'h15c;
        src60 <= 12'h844;
        src61 <= 12'h54c;
        src62 <= 12'hab4;
        src63 <= 12'h745;
        src64 <= 12'hf3c;
        src65 <= 12'h393;
        src66 <= 12'h202;
        src67 <= 12'h859;
        src68 <= 12'hf5c;
        src69 <= 12'h439;
        src70 <= 12'h142;
        src71 <= 12'h1de;
        src72 <= 12'hbd;
        src73 <= 12'hba4;
        src74 <= 12'h772;
        src75 <= 12'ha4;
        src76 <= 12'h5e2;
        src77 <= 12'hd51;
        src78 <= 12'h161;
        src79 <= 12'h114;
        src80 <= 12'h122;
        src81 <= 12'h332;
        src82 <= 12'h176;
        src83 <= 12'h27c;
        src84 <= 12'h213;
        src85 <= 12'h3cd;
        src86 <= 12'h5c;
        src87 <= 12'h44d;
        src88 <= 12'h6bb;
        src89 <= 12'h484;
        src90 <= 12'h4;
        src91 <= 12'h8d;
        src92 <= 12'h77c;
        src93 <= 12'hf15;
        src94 <= 12'h96d;
        src95 <= 12'hd21;
        src96 <= 12'hf68;
        src97 <= 12'hec5;
        src98 <= 12'h288;
        src99 <= 12'h30a;
        src100 <= 12'he67;
        src101 <= 12'h6df;
        src102 <= 12'h5a5;
        src103 <= 12'h17a;
        src104 <= 12'h81f;
        src105 <= 12'h42a;
        src106 <= 12'h320;
        src107 <= 12'h560;
        src108 <= 12'hc9;
        src109 <= 12'hedf;
        src110 <= 12'h4d6;
        src111 <= 12'h8e6;
        src112 <= 12'hd95;
        src113 <= 12'h915;
        src114 <= 12'h824;
        src115 <= 12'h9d2;
        src116 <= 12'hd77;
        src117 <= 12'ha55;
        src118 <= 12'hef5;
        src119 <= 12'h6cf;
        src120 <= 12'h121;
        src121 <= 12'h5b8;
        src122 <= 12'h827;
        src123 <= 12'hd4f;
        src124 <= 12'h5e8;
        src125 <= 12'h69b;
        src126 <= 12'h77d;
        src127 <= 12'h7f7;
        exp <= 19'h381f9;
        #1
        src0 <= 12'hb16;
        src1 <= 12'h5b5;
        src2 <= 12'h5ea;
        src3 <= 12'hfd4;
        src4 <= 12'hf9e;
        src5 <= 12'h997;
        src6 <= 12'hfe9;
        src7 <= 12'ha25;
        src8 <= 12'hfa0;
        src9 <= 12'h51e;
        src10 <= 12'hdc6;
        src11 <= 12'h1c3;
        src12 <= 12'hc40;
        src13 <= 12'h6ce;
        src14 <= 12'ha5d;
        src15 <= 12'h36a;
        src16 <= 12'h181;
        src17 <= 12'h896;
        src18 <= 12'h59e;
        src19 <= 12'h42f;
        src20 <= 12'h8dc;
        src21 <= 12'h77d;
        src22 <= 12'h664;
        src23 <= 12'hba9;
        src24 <= 12'h95f;
        src25 <= 12'h1b4;
        src26 <= 12'h6df;
        src27 <= 12'h844;
        src28 <= 12'h442;
        src29 <= 12'hc89;
        src30 <= 12'hff1;
        src31 <= 12'h502;
        src32 <= 12'hc48;
        src33 <= 12'h462;
        src34 <= 12'hfcc;
        src35 <= 12'h82f;
        src36 <= 12'h6d5;
        src37 <= 12'h92e;
        src38 <= 12'h539;
        src39 <= 12'h279;
        src40 <= 12'h16b;
        src41 <= 12'h890;
        src42 <= 12'h3f6;
        src43 <= 12'h58d;
        src44 <= 12'h22b;
        src45 <= 12'h8c1;
        src46 <= 12'h2d9;
        src47 <= 12'h221;
        src48 <= 12'h6dd;
        src49 <= 12'he2c;
        src50 <= 12'hd5a;
        src51 <= 12'hbb0;
        src52 <= 12'h4f9;
        src53 <= 12'h4a5;
        src54 <= 12'h76c;
        src55 <= 12'hf29;
        src56 <= 12'h428;
        src57 <= 12'hbb8;
        src58 <= 12'h227;
        src59 <= 12'hdbc;
        src60 <= 12'h667;
        src61 <= 12'he41;
        src62 <= 12'h905;
        src63 <= 12'h2c3;
        src64 <= 12'h891;
        src65 <= 12'h8f8;
        src66 <= 12'ha95;
        src67 <= 12'he3d;
        src68 <= 12'h748;
        src69 <= 12'h86a;
        src70 <= 12'h8c7;
        src71 <= 12'h5ef;
        src72 <= 12'h95f;
        src73 <= 12'hc33;
        src74 <= 12'h42b;
        src75 <= 12'h5c2;
        src76 <= 12'hda3;
        src77 <= 12'h22f;
        src78 <= 12'h3d0;
        src79 <= 12'hea8;
        src80 <= 12'h407;
        src81 <= 12'h84f;
        src82 <= 12'ha43;
        src83 <= 12'hd14;
        src84 <= 12'h360;
        src85 <= 12'hd7c;
        src86 <= 12'h326;
        src87 <= 12'hb35;
        src88 <= 12'h9e3;
        src89 <= 12'hf88;
        src90 <= 12'h9cb;
        src91 <= 12'h435;
        src92 <= 12'h1d2;
        src93 <= 12'h24d;
        src94 <= 12'he3b;
        src95 <= 12'he30;
        src96 <= 12'h375;
        src97 <= 12'hc1e;
        src98 <= 12'h115;
        src99 <= 12'h271;
        src100 <= 12'h748;
        src101 <= 12'ha44;
        src102 <= 12'h229;
        src103 <= 12'h4c2;
        src104 <= 12'hb7;
        src105 <= 12'hef;
        src106 <= 12'h822;
        src107 <= 12'h2bc;
        src108 <= 12'h99a;
        src109 <= 12'h5ea;
        src110 <= 12'he40;
        src111 <= 12'h80c;
        src112 <= 12'hab1;
        src113 <= 12'h758;
        src114 <= 12'hf07;
        src115 <= 12'hec4;
        src116 <= 12'h563;
        src117 <= 12'hd5a;
        src118 <= 12'h794;
        src119 <= 12'hd1;
        src120 <= 12'hd87;
        src121 <= 12'hfad;
        src122 <= 12'h258;
        src123 <= 12'he3e;
        src124 <= 12'h196;
        src125 <= 12'h8c9;
        src126 <= 12'h76;
        src127 <= 12'ha88;
        exp <= 19'h408c3;
        #1
        src0 <= 12'h4f3;
        src1 <= 12'h752;
        src2 <= 12'h299;
        src3 <= 12'hea9;
        src4 <= 12'h512;
        src5 <= 12'hccb;
        src6 <= 12'h79c;
        src7 <= 12'h881;
        src8 <= 12'ha6;
        src9 <= 12'he37;
        src10 <= 12'hec6;
        src11 <= 12'h738;
        src12 <= 12'ha0e;
        src13 <= 12'h434;
        src14 <= 12'hbfe;
        src15 <= 12'h43d;
        src16 <= 12'h9a7;
        src17 <= 12'h99d;
        src18 <= 12'h88b;
        src19 <= 12'he95;
        src20 <= 12'hf9d;
        src21 <= 12'h535;
        src22 <= 12'h5d8;
        src23 <= 12'h606;
        src24 <= 12'hc27;
        src25 <= 12'h275;
        src26 <= 12'h1c8;
        src27 <= 12'h2c8;
        src28 <= 12'hca;
        src29 <= 12'hc3a;
        src30 <= 12'h6cc;
        src31 <= 12'h756;
        src32 <= 12'h4e;
        src33 <= 12'hd4e;
        src34 <= 12'hff5;
        src35 <= 12'h5ca;
        src36 <= 12'h5f;
        src37 <= 12'h85e;
        src38 <= 12'ha8d;
        src39 <= 12'h1d4;
        src40 <= 12'h380;
        src41 <= 12'h7c6;
        src42 <= 12'h554;
        src43 <= 12'hea;
        src44 <= 12'h18f;
        src45 <= 12'h537;
        src46 <= 12'h75d;
        src47 <= 12'hff4;
        src48 <= 12'ha57;
        src49 <= 12'h777;
        src50 <= 12'h6e2;
        src51 <= 12'ha5;
        src52 <= 12'h5d3;
        src53 <= 12'h20c;
        src54 <= 12'h1e;
        src55 <= 12'hd07;
        src56 <= 12'he67;
        src57 <= 12'hf7c;
        src58 <= 12'hfd3;
        src59 <= 12'h116;
        src60 <= 12'hd98;
        src61 <= 12'hde3;
        src62 <= 12'hc1a;
        src63 <= 12'h52b;
        src64 <= 12'hf58;
        src65 <= 12'hf3f;
        src66 <= 12'hb4d;
        src67 <= 12'hf9c;
        src68 <= 12'h6d6;
        src69 <= 12'h27c;
        src70 <= 12'h81d;
        src71 <= 12'h573;
        src72 <= 12'h561;
        src73 <= 12'h77b;
        src74 <= 12'h2f6;
        src75 <= 12'h829;
        src76 <= 12'h7df;
        src77 <= 12'hbb7;
        src78 <= 12'hb8d;
        src79 <= 12'h9bc;
        src80 <= 12'hd1d;
        src81 <= 12'h78d;
        src82 <= 12'h96a;
        src83 <= 12'h8c2;
        src84 <= 12'h4d4;
        src85 <= 12'hdc3;
        src86 <= 12'h5a7;
        src87 <= 12'hdc4;
        src88 <= 12'h5a9;
        src89 <= 12'h79c;
        src90 <= 12'h5dd;
        src91 <= 12'h668;
        src92 <= 12'had8;
        src93 <= 12'h6d6;
        src94 <= 12'hfff;
        src95 <= 12'h5f0;
        src96 <= 12'heae;
        src97 <= 12'h3fa;
        src98 <= 12'h5d3;
        src99 <= 12'h7dc;
        src100 <= 12'h9f0;
        src101 <= 12'hf0d;
        src102 <= 12'h3e7;
        src103 <= 12'hd20;
        src104 <= 12'he7e;
        src105 <= 12'h5b0;
        src106 <= 12'hfa;
        src107 <= 12'haa8;
        src108 <= 12'h943;
        src109 <= 12'h93;
        src110 <= 12'h886;
        src111 <= 12'h57d;
        src112 <= 12'h360;
        src113 <= 12'hea;
        src114 <= 12'h613;
        src115 <= 12'h829;
        src116 <= 12'h147;
        src117 <= 12'h97d;
        src118 <= 12'hf03;
        src119 <= 12'hacd;
        src120 <= 12'h47b;
        src121 <= 12'had6;
        src122 <= 12'h5a7;
        src123 <= 12'hb1d;
        src124 <= 12'h85e;
        src125 <= 12'h5a5;
        src126 <= 12'h5c6;
        src127 <= 12'h6f4;
        exp <= 19'h40163;
        #1
        src0 <= 12'hc9e;
        src1 <= 12'hc35;
        src2 <= 12'h4bc;
        src3 <= 12'h623;
        src4 <= 12'hc5f;
        src5 <= 12'h4a2;
        src6 <= 12'he9c;
        src7 <= 12'h527;
        src8 <= 12'h8df;
        src9 <= 12'h5c1;
        src10 <= 12'hb64;
        src11 <= 12'hb00;
        src12 <= 12'h9b3;
        src13 <= 12'h478;
        src14 <= 12'hdd0;
        src15 <= 12'h289;
        src16 <= 12'h25;
        src17 <= 12'h991;
        src18 <= 12'hff8;
        src19 <= 12'hf09;
        src20 <= 12'h36;
        src21 <= 12'haad;
        src22 <= 12'h825;
        src23 <= 12'h91a;
        src24 <= 12'hddd;
        src25 <= 12'h474;
        src26 <= 12'ha50;
        src27 <= 12'hc37;
        src28 <= 12'he0d;
        src29 <= 12'h8d8;
        src30 <= 12'hae8;
        src31 <= 12'hcad;
        src32 <= 12'hf91;
        src33 <= 12'he0;
        src34 <= 12'h855;
        src35 <= 12'h66d;
        src36 <= 12'hb33;
        src37 <= 12'he38;
        src38 <= 12'h90;
        src39 <= 12'hc10;
        src40 <= 12'h451;
        src41 <= 12'h9ce;
        src42 <= 12'h448;
        src43 <= 12'h9ab;
        src44 <= 12'h7d6;
        src45 <= 12'ha22;
        src46 <= 12'hf51;
        src47 <= 12'hc5b;
        src48 <= 12'h4af;
        src49 <= 12'h946;
        src50 <= 12'h714;
        src51 <= 12'h7bf;
        src52 <= 12'hc25;
        src53 <= 12'hfe1;
        src54 <= 12'h434;
        src55 <= 12'hb88;
        src56 <= 12'h6f1;
        src57 <= 12'h237;
        src58 <= 12'h1b2;
        src59 <= 12'h1d3;
        src60 <= 12'h86b;
        src61 <= 12'h66b;
        src62 <= 12'h8ad;
        src63 <= 12'h864;
        src64 <= 12'hc75;
        src65 <= 12'he7f;
        src66 <= 12'hc6b;
        src67 <= 12'ha77;
        src68 <= 12'hcf7;
        src69 <= 12'ha0;
        src70 <= 12'ha90;
        src71 <= 12'hb3c;
        src72 <= 12'hda6;
        src73 <= 12'h80a;
        src74 <= 12'h5d3;
        src75 <= 12'h124;
        src76 <= 12'h9b0;
        src77 <= 12'h74b;
        src78 <= 12'h7c0;
        src79 <= 12'hff5;
        src80 <= 12'h29d;
        src81 <= 12'ha3;
        src82 <= 12'ha5a;
        src83 <= 12'ha5;
        src84 <= 12'hd93;
        src85 <= 12'h8fe;
        src86 <= 12'hee5;
        src87 <= 12'hfa8;
        src88 <= 12'hfd0;
        src89 <= 12'hbcf;
        src90 <= 12'haa3;
        src91 <= 12'h188;
        src92 <= 12'hba9;
        src93 <= 12'h5aa;
        src94 <= 12'h46d;
        src95 <= 12'h294;
        src96 <= 12'hb51;
        src97 <= 12'he17;
        src98 <= 12'hde2;
        src99 <= 12'h31d;
        src100 <= 12'hfc5;
        src101 <= 12'h729;
        src102 <= 12'h923;
        src103 <= 12'hd22;
        src104 <= 12'hf21;
        src105 <= 12'h7a2;
        src106 <= 12'h770;
        src107 <= 12'h111;
        src108 <= 12'h2c1;
        src109 <= 12'h5d9;
        src110 <= 12'h1ef;
        src111 <= 12'hed8;
        src112 <= 12'h581;
        src113 <= 12'hf18;
        src114 <= 12'h552;
        src115 <= 12'hbb6;
        src116 <= 12'h980;
        src117 <= 12'h6b8;
        src118 <= 12'h495;
        src119 <= 12'h9b5;
        src120 <= 12'hd8a;
        src121 <= 12'hd72;
        src122 <= 12'h470;
        src123 <= 12'hd78;
        src124 <= 12'hc6f;
        src125 <= 12'h73d;
        src126 <= 12'h275;
        src127 <= 12'h83f;
        exp <= 19'h469ec;
        #1
        src0 <= 12'h391;
        src1 <= 12'h3b0;
        src2 <= 12'h18d;
        src3 <= 12'hdb7;
        src4 <= 12'h226;
        src5 <= 12'h26;
        src6 <= 12'h61b;
        src7 <= 12'h61a;
        src8 <= 12'hfbb;
        src9 <= 12'hac9;
        src10 <= 12'h779;
        src11 <= 12'h43b;
        src12 <= 12'he77;
        src13 <= 12'hfab;
        src14 <= 12'h49c;
        src15 <= 12'hc20;
        src16 <= 12'hcca;
        src17 <= 12'he96;
        src18 <= 12'h130;
        src19 <= 12'h883;
        src20 <= 12'hcde;
        src21 <= 12'h3ea;
        src22 <= 12'h804;
        src23 <= 12'hc4d;
        src24 <= 12'hcec;
        src25 <= 12'h30d;
        src26 <= 12'h270;
        src27 <= 12'hf9e;
        src28 <= 12'h3e5;
        src29 <= 12'haf;
        src30 <= 12'h7a9;
        src31 <= 12'hcc9;
        src32 <= 12'h22;
        src33 <= 12'heb0;
        src34 <= 12'h17;
        src35 <= 12'hd8d;
        src36 <= 12'h366;
        src37 <= 12'hcab;
        src38 <= 12'h6bd;
        src39 <= 12'h949;
        src40 <= 12'h7a8;
        src41 <= 12'he5e;
        src42 <= 12'h404;
        src43 <= 12'h835;
        src44 <= 12'h876;
        src45 <= 12'h89a;
        src46 <= 12'h38b;
        src47 <= 12'hfb2;
        src48 <= 12'h9bd;
        src49 <= 12'h13d;
        src50 <= 12'h882;
        src51 <= 12'h2a5;
        src52 <= 12'h792;
        src53 <= 12'hdb2;
        src54 <= 12'heee;
        src55 <= 12'hb52;
        src56 <= 12'h5b3;
        src57 <= 12'hac5;
        src58 <= 12'h706;
        src59 <= 12'h3da;
        src60 <= 12'h6e;
        src61 <= 12'hfd3;
        src62 <= 12'h817;
        src63 <= 12'hfe6;
        src64 <= 12'hf32;
        src65 <= 12'hfe0;
        src66 <= 12'hed8;
        src67 <= 12'h890;
        src68 <= 12'hdfb;
        src69 <= 12'hb45;
        src70 <= 12'h5d1;
        src71 <= 12'h123;
        src72 <= 12'h923;
        src73 <= 12'h19d;
        src74 <= 12'hfe6;
        src75 <= 12'ha54;
        src76 <= 12'h3e6;
        src77 <= 12'hbab;
        src78 <= 12'he44;
        src79 <= 12'hd51;
        src80 <= 12'ha37;
        src81 <= 12'h8ef;
        src82 <= 12'hff1;
        src83 <= 12'h914;
        src84 <= 12'hde4;
        src85 <= 12'hcea;
        src86 <= 12'hbef;
        src87 <= 12'h417;
        src88 <= 12'h3c9;
        src89 <= 12'hee6;
        src90 <= 12'h626;
        src91 <= 12'h869;
        src92 <= 12'hf9b;
        src93 <= 12'h61c;
        src94 <= 12'h624;
        src95 <= 12'h4d3;
        src96 <= 12'h5be;
        src97 <= 12'hf98;
        src98 <= 12'h358;
        src99 <= 12'h467;
        src100 <= 12'hd03;
        src101 <= 12'ha28;
        src102 <= 12'h319;
        src103 <= 12'h714;
        src104 <= 12'hcc3;
        src105 <= 12'hf16;
        src106 <= 12'hc15;
        src107 <= 12'h9eb;
        src108 <= 12'hda0;
        src109 <= 12'h641;
        src110 <= 12'hdb7;
        src111 <= 12'hf08;
        src112 <= 12'h276;
        src113 <= 12'h8d3;
        src114 <= 12'hdb8;
        src115 <= 12'h2f3;
        src116 <= 12'h8f6;
        src117 <= 12'h5fb;
        src118 <= 12'h1fc;
        src119 <= 12'h1fa;
        src120 <= 12'head;
        src121 <= 12'h2f9;
        src122 <= 12'hed0;
        src123 <= 12'hd9f;
        src124 <= 12'hdea;
        src125 <= 12'hc52;
        src126 <= 12'h1d9;
        src127 <= 12'hd8f;
        exp <= 19'h472dc;
        #1
        src0 <= 12'hee2;
        src1 <= 12'h9f5;
        src2 <= 12'h1f9;
        src3 <= 12'he8f;
        src4 <= 12'haf4;
        src5 <= 12'hbfc;
        src6 <= 12'h22c;
        src7 <= 12'h47e;
        src8 <= 12'hbaf;
        src9 <= 12'h1d8;
        src10 <= 12'h3f;
        src11 <= 12'hb6a;
        src12 <= 12'h70e;
        src13 <= 12'hd72;
        src14 <= 12'h4fc;
        src15 <= 12'hfc;
        src16 <= 12'h797;
        src17 <= 12'h23b;
        src18 <= 12'h58e;
        src19 <= 12'he54;
        src20 <= 12'h558;
        src21 <= 12'heb7;
        src22 <= 12'h145;
        src23 <= 12'he61;
        src24 <= 12'h859;
        src25 <= 12'hbf0;
        src26 <= 12'hcc7;
        src27 <= 12'h1f2;
        src28 <= 12'h70;
        src29 <= 12'hc6d;
        src30 <= 12'h45;
        src31 <= 12'h54f;
        src32 <= 12'hedb;
        src33 <= 12'h169;
        src34 <= 12'hced;
        src35 <= 12'ha7e;
        src36 <= 12'hc6f;
        src37 <= 12'hb18;
        src38 <= 12'h785;
        src39 <= 12'hc8;
        src40 <= 12'h199;
        src41 <= 12'ha1;
        src42 <= 12'h356;
        src43 <= 12'h431;
        src44 <= 12'hd31;
        src45 <= 12'h197;
        src46 <= 12'h2ff;
        src47 <= 12'h506;
        src48 <= 12'h17b;
        src49 <= 12'h2b6;
        src50 <= 12'hcb7;
        src51 <= 12'hd3c;
        src52 <= 12'hdbe;
        src53 <= 12'hc2a;
        src54 <= 12'h92a;
        src55 <= 12'hdbe;
        src56 <= 12'hbaa;
        src57 <= 12'h193;
        src58 <= 12'he5f;
        src59 <= 12'hddd;
        src60 <= 12'hcba;
        src61 <= 12'h6ce;
        src62 <= 12'h790;
        src63 <= 12'h29f;
        src64 <= 12'h159;
        src65 <= 12'hd81;
        src66 <= 12'ha0b;
        src67 <= 12'hdec;
        src68 <= 12'hcad;
        src69 <= 12'h750;
        src70 <= 12'hd0b;
        src71 <= 12'h816;
        src72 <= 12'h666;
        src73 <= 12'h8e0;
        src74 <= 12'h71d;
        src75 <= 12'h793;
        src76 <= 12'hfa8;
        src77 <= 12'h411;
        src78 <= 12'h647;
        src79 <= 12'hbea;
        src80 <= 12'h219;
        src81 <= 12'h12e;
        src82 <= 12'h1b7;
        src83 <= 12'h58c;
        src84 <= 12'ha3d;
        src85 <= 12'he91;
        src86 <= 12'ha22;
        src87 <= 12'hb78;
        src88 <= 12'h32b;
        src89 <= 12'h1a2;
        src90 <= 12'hbb3;
        src91 <= 12'hd4c;
        src92 <= 12'hc7d;
        src93 <= 12'h281;
        src94 <= 12'hc30;
        src95 <= 12'h39e;
        src96 <= 12'h7a2;
        src97 <= 12'h102;
        src98 <= 12'hb02;
        src99 <= 12'hfb9;
        src100 <= 12'h1e3;
        src101 <= 12'h6ed;
        src102 <= 12'h7f2;
        src103 <= 12'ha5d;
        src104 <= 12'h24c;
        src105 <= 12'heb4;
        src106 <= 12'h3ec;
        src107 <= 12'hc3b;
        src108 <= 12'hbaf;
        src109 <= 12'h992;
        src110 <= 12'h73e;
        src111 <= 12'haea;
        src112 <= 12'h41d;
        src113 <= 12'hd3f;
        src114 <= 12'h6f9;
        src115 <= 12'h93f;
        src116 <= 12'h18;
        src117 <= 12'hd4a;
        src118 <= 12'h112;
        src119 <= 12'h87a;
        src120 <= 12'hf8d;
        src121 <= 12'h653;
        src122 <= 12'h3fe;
        src123 <= 12'he2f;
        src124 <= 12'ha3b;
        src125 <= 12'h22f;
        src126 <= 12'hb91;
        src127 <= 12'h8e6;
        exp <= 19'h40189;
        #1
        src0 <= 12'hd83;
        src1 <= 12'h871;
        src2 <= 12'hcea;
        src3 <= 12'h740;
        src4 <= 12'hf26;
        src5 <= 12'ha7b;
        src6 <= 12'h1e8;
        src7 <= 12'hb2b;
        src8 <= 12'h9d7;
        src9 <= 12'h115;
        src10 <= 12'hc88;
        src11 <= 12'h3b0;
        src12 <= 12'h2bc;
        src13 <= 12'h4bf;
        src14 <= 12'h5af;
        src15 <= 12'ha83;
        src16 <= 12'h7c9;
        src17 <= 12'hc84;
        src18 <= 12'he79;
        src19 <= 12'hbb2;
        src20 <= 12'h726;
        src21 <= 12'he1;
        src22 <= 12'h1ca;
        src23 <= 12'hebf;
        src24 <= 12'hee8;
        src25 <= 12'hb0;
        src26 <= 12'hd4c;
        src27 <= 12'hccb;
        src28 <= 12'h8ad;
        src29 <= 12'hdf;
        src30 <= 12'he59;
        src31 <= 12'h1dc;
        src32 <= 12'hf4e;
        src33 <= 12'hd82;
        src34 <= 12'h23e;
        src35 <= 12'h463;
        src36 <= 12'hd2b;
        src37 <= 12'hae6;
        src38 <= 12'hdb9;
        src39 <= 12'h4ac;
        src40 <= 12'hf75;
        src41 <= 12'h6fe;
        src42 <= 12'h873;
        src43 <= 12'hf24;
        src44 <= 12'hc8;
        src45 <= 12'h4da;
        src46 <= 12'ha74;
        src47 <= 12'he78;
        src48 <= 12'h6d9;
        src49 <= 12'hde8;
        src50 <= 12'ha06;
        src51 <= 12'h514;
        src52 <= 12'h8b0;
        src53 <= 12'hf16;
        src54 <= 12'h700;
        src55 <= 12'hd61;
        src56 <= 12'hb50;
        src57 <= 12'h1a9;
        src58 <= 12'h233;
        src59 <= 12'h17e;
        src60 <= 12'h97b;
        src61 <= 12'h602;
        src62 <= 12'h52b;
        src63 <= 12'h3ca;
        src64 <= 12'h8ee;
        src65 <= 12'hcda;
        src66 <= 12'h68b;
        src67 <= 12'heee;
        src68 <= 12'hc71;
        src69 <= 12'hf73;
        src70 <= 12'hda4;
        src71 <= 12'h68d;
        src72 <= 12'ha05;
        src73 <= 12'h23c;
        src74 <= 12'h6af;
        src75 <= 12'h43;
        src76 <= 12'h43a;
        src77 <= 12'h27f;
        src78 <= 12'h325;
        src79 <= 12'h2cc;
        src80 <= 12'hbe0;
        src81 <= 12'h1e7;
        src82 <= 12'hb42;
        src83 <= 12'h1df;
        src84 <= 12'h1f6;
        src85 <= 12'hf88;
        src86 <= 12'ha9f;
        src87 <= 12'hb6;
        src88 <= 12'h974;
        src89 <= 12'he0b;
        src90 <= 12'h8b6;
        src91 <= 12'h761;
        src92 <= 12'ha2f;
        src93 <= 12'h41e;
        src94 <= 12'h58e;
        src95 <= 12'h9a6;
        src96 <= 12'h778;
        src97 <= 12'ha03;
        src98 <= 12'hdcb;
        src99 <= 12'h176;
        src100 <= 12'hd5d;
        src101 <= 12'h5b6;
        src102 <= 12'hfbc;
        src103 <= 12'hdb4;
        src104 <= 12'hcbe;
        src105 <= 12'h88a;
        src106 <= 12'h7b3;
        src107 <= 12'h9fc;
        src108 <= 12'hf0b;
        src109 <= 12'hc01;
        src110 <= 12'hd5e;
        src111 <= 12'h6e8;
        src112 <= 12'h3b9;
        src113 <= 12'h1e7;
        src114 <= 12'h4af;
        src115 <= 12'hc41;
        src116 <= 12'he3a;
        src117 <= 12'hd46;
        src118 <= 12'hec9;
        src119 <= 12'h1bb;
        src120 <= 12'he5f;
        src121 <= 12'h426;
        src122 <= 12'haba;
        src123 <= 12'hc5;
        src124 <= 12'ha1e;
        src125 <= 12'hd89;
        src126 <= 12'hbb5;
        src127 <= 12'h166;
        exp <= 19'h4469f;
        #1
        src0 <= 12'h1d7;
        src1 <= 12'he34;
        src2 <= 12'hc52;
        src3 <= 12'h2fd;
        src4 <= 12'h749;
        src5 <= 12'he16;
        src6 <= 12'hb70;
        src7 <= 12'h54d;
        src8 <= 12'hd58;
        src9 <= 12'h717;
        src10 <= 12'hbe3;
        src11 <= 12'h28f;
        src12 <= 12'ha3d;
        src13 <= 12'hf3e;
        src14 <= 12'hbc8;
        src15 <= 12'hc06;
        src16 <= 12'h978;
        src17 <= 12'h646;
        src18 <= 12'haea;
        src19 <= 12'h9de;
        src20 <= 12'hd18;
        src21 <= 12'h2da;
        src22 <= 12'h647;
        src23 <= 12'h8bb;
        src24 <= 12'ha3a;
        src25 <= 12'h404;
        src26 <= 12'h6;
        src27 <= 12'hdbf;
        src28 <= 12'h525;
        src29 <= 12'h9f4;
        src30 <= 12'h680;
        src31 <= 12'h293;
        src32 <= 12'hf31;
        src33 <= 12'h306;
        src34 <= 12'hdd1;
        src35 <= 12'h4b6;
        src36 <= 12'h1bb;
        src37 <= 12'hb39;
        src38 <= 12'hc54;
        src39 <= 12'h651;
        src40 <= 12'hbc6;
        src41 <= 12'h67c;
        src42 <= 12'h25;
        src43 <= 12'hacf;
        src44 <= 12'h1dc;
        src45 <= 12'hdb9;
        src46 <= 12'hacf;
        src47 <= 12'h5f6;
        src48 <= 12'h51;
        src49 <= 12'hfbf;
        src50 <= 12'hd3a;
        src51 <= 12'ha4e;
        src52 <= 12'h626;
        src53 <= 12'h58c;
        src54 <= 12'hc08;
        src55 <= 12'h78d;
        src56 <= 12'h20f;
        src57 <= 12'h3de;
        src58 <= 12'h834;
        src59 <= 12'h510;
        src60 <= 12'haba;
        src61 <= 12'h4fa;
        src62 <= 12'habd;
        src63 <= 12'h64b;
        src64 <= 12'h39b;
        src65 <= 12'h447;
        src66 <= 12'ha02;
        src67 <= 12'h7fb;
        src68 <= 12'h6e2;
        src69 <= 12'hdf4;
        src70 <= 12'hd90;
        src71 <= 12'h2d0;
        src72 <= 12'hede;
        src73 <= 12'hc3d;
        src74 <= 12'h177;
        src75 <= 12'hfb3;
        src76 <= 12'h864;
        src77 <= 12'h6d4;
        src78 <= 12'h973;
        src79 <= 12'h4cb;
        src80 <= 12'hd26;
        src81 <= 12'h447;
        src82 <= 12'he6;
        src83 <= 12'h99e;
        src84 <= 12'h62e;
        src85 <= 12'hb23;
        src86 <= 12'h8bb;
        src87 <= 12'h901;
        src88 <= 12'h50d;
        src89 <= 12'h4f6;
        src90 <= 12'h516;
        src91 <= 12'hc0a;
        src92 <= 12'h84c;
        src93 <= 12'hab7;
        src94 <= 12'h26e;
        src95 <= 12'h38f;
        src96 <= 12'h6be;
        src97 <= 12'h77;
        src98 <= 12'h39c;
        src99 <= 12'h4b0;
        src100 <= 12'h20b;
        src101 <= 12'h99f;
        src102 <= 12'h765;
        src103 <= 12'h55;
        src104 <= 12'hc38;
        src105 <= 12'h61;
        src106 <= 12'h712;
        src107 <= 12'h519;
        src108 <= 12'h1ad;
        src109 <= 12'h846;
        src110 <= 12'hc5a;
        src111 <= 12'h1d0;
        src112 <= 12'hd32;
        src113 <= 12'he63;
        src114 <= 12'he55;
        src115 <= 12'h30b;
        src116 <= 12'h5b;
        src117 <= 12'heb5;
        src118 <= 12'h3d2;
        src119 <= 12'h50b;
        src120 <= 12'he33;
        src121 <= 12'h5db;
        src122 <= 12'h6d6;
        src123 <= 12'he3c;
        src124 <= 12'hc4c;
        src125 <= 12'h82b;
        src126 <= 12'h896;
        src127 <= 12'hc54;
        exp <= 19'h3f516;
        #1
        src0 <= 12'h4ca;
        src1 <= 12'h3e3;
        src2 <= 12'ha2a;
        src3 <= 12'hcf9;
        src4 <= 12'hcf9;
        src5 <= 12'h66f;
        src6 <= 12'hedf;
        src7 <= 12'hbb7;
        src8 <= 12'hc34;
        src9 <= 12'h9ae;
        src10 <= 12'h7fd;
        src11 <= 12'hbcc;
        src12 <= 12'h53d;
        src13 <= 12'h490;
        src14 <= 12'hd39;
        src15 <= 12'h2ce;
        src16 <= 12'heb1;
        src17 <= 12'h51c;
        src18 <= 12'h59f;
        src19 <= 12'h48;
        src20 <= 12'hc9c;
        src21 <= 12'hf7b;
        src22 <= 12'h314;
        src23 <= 12'h9ed;
        src24 <= 12'h746;
        src25 <= 12'h35f;
        src26 <= 12'h488;
        src27 <= 12'h46e;
        src28 <= 12'hd6b;
        src29 <= 12'h665;
        src30 <= 12'h903;
        src31 <= 12'he02;
        src32 <= 12'h45f;
        src33 <= 12'h8f6;
        src34 <= 12'h34d;
        src35 <= 12'h8e0;
        src36 <= 12'hb4b;
        src37 <= 12'hec9;
        src38 <= 12'hc0f;
        src39 <= 12'hf8d;
        src40 <= 12'hf5b;
        src41 <= 12'h6c2;
        src42 <= 12'hb2;
        src43 <= 12'hc7b;
        src44 <= 12'h236;
        src45 <= 12'h1c8;
        src46 <= 12'h269;
        src47 <= 12'h4f;
        src48 <= 12'h5c2;
        src49 <= 12'he6a;
        src50 <= 12'hc67;
        src51 <= 12'hbc0;
        src52 <= 12'h9ca;
        src53 <= 12'h53c;
        src54 <= 12'h2e5;
        src55 <= 12'h64a;
        src56 <= 12'h951;
        src57 <= 12'h833;
        src58 <= 12'hcc4;
        src59 <= 12'h2ab;
        src60 <= 12'h84c;
        src61 <= 12'hfe5;
        src62 <= 12'h5da;
        src63 <= 12'ha39;
        src64 <= 12'hf92;
        src65 <= 12'hf30;
        src66 <= 12'h971;
        src67 <= 12'hb38;
        src68 <= 12'h3e5;
        src69 <= 12'he3f;
        src70 <= 12'h7fd;
        src71 <= 12'h6e7;
        src72 <= 12'h34a;
        src73 <= 12'h464;
        src74 <= 12'h2;
        src75 <= 12'h245;
        src76 <= 12'h757;
        src77 <= 12'h2bd;
        src78 <= 12'h4b5;
        src79 <= 12'h27c;
        src80 <= 12'hd93;
        src81 <= 12'hf33;
        src82 <= 12'h4d5;
        src83 <= 12'hb52;
        src84 <= 12'h9b9;
        src85 <= 12'h15b;
        src86 <= 12'h840;
        src87 <= 12'h857;
        src88 <= 12'h310;
        src89 <= 12'hf2e;
        src90 <= 12'he9a;
        src91 <= 12'hab3;
        src92 <= 12'h3f7;
        src93 <= 12'hc9a;
        src94 <= 12'h909;
        src95 <= 12'h16e;
        src96 <= 12'hb48;
        src97 <= 12'h85f;
        src98 <= 12'h145;
        src99 <= 12'h761;
        src100 <= 12'hf0f;
        src101 <= 12'hb00;
        src102 <= 12'h7ec;
        src103 <= 12'haa3;
        src104 <= 12'hf56;
        src105 <= 12'hcdb;
        src106 <= 12'h83f;
        src107 <= 12'h9b;
        src108 <= 12'h108;
        src109 <= 12'h5b6;
        src110 <= 12'he5b;
        src111 <= 12'h389;
        src112 <= 12'h816;
        src113 <= 12'h105;
        src114 <= 12'h9cb;
        src115 <= 12'hc28;
        src116 <= 12'hf93;
        src117 <= 12'h945;
        src118 <= 12'h265;
        src119 <= 12'h7f5;
        src120 <= 12'h42c;
        src121 <= 12'h309;
        src122 <= 12'h98b;
        src123 <= 12'h1d2;
        src124 <= 12'h37d;
        src125 <= 12'hc60;
        src126 <= 12'ha18;
        src127 <= 12'h28;
        exp <= 19'h40dd9;
        #1
        src0 <= 12'hf91;
        src1 <= 12'hc14;
        src2 <= 12'h32c;
        src3 <= 12'hc3;
        src4 <= 12'h641;
        src5 <= 12'hf79;
        src6 <= 12'h409;
        src7 <= 12'h2c;
        src8 <= 12'h4e6;
        src9 <= 12'hef4;
        src10 <= 12'h1cf;
        src11 <= 12'h274;
        src12 <= 12'h9b0;
        src13 <= 12'hf1c;
        src14 <= 12'hde4;
        src15 <= 12'h5d3;
        src16 <= 12'h6b8;
        src17 <= 12'h9e2;
        src18 <= 12'h91c;
        src19 <= 12'h1cb;
        src20 <= 12'hdcc;
        src21 <= 12'h2e5;
        src22 <= 12'h49f;
        src23 <= 12'h5df;
        src24 <= 12'h77c;
        src25 <= 12'hd96;
        src26 <= 12'h128;
        src27 <= 12'h586;
        src28 <= 12'h8dc;
        src29 <= 12'he8e;
        src30 <= 12'h79e;
        src31 <= 12'h476;
        src32 <= 12'h2d0;
        src33 <= 12'h334;
        src34 <= 12'h9e;
        src35 <= 12'h9b3;
        src36 <= 12'h9db;
        src37 <= 12'h530;
        src38 <= 12'hc98;
        src39 <= 12'hd90;
        src40 <= 12'h778;
        src41 <= 12'he73;
        src42 <= 12'h3f9;
        src43 <= 12'h9f4;
        src44 <= 12'h112;
        src45 <= 12'hfe2;
        src46 <= 12'h451;
        src47 <= 12'h1cc;
        src48 <= 12'h61c;
        src49 <= 12'h37d;
        src50 <= 12'h4e3;
        src51 <= 12'h485;
        src52 <= 12'h884;
        src53 <= 12'he29;
        src54 <= 12'hdc0;
        src55 <= 12'ha81;
        src56 <= 12'h6a2;
        src57 <= 12'had0;
        src58 <= 12'hc6c;
        src59 <= 12'hd5e;
        src60 <= 12'h7a2;
        src61 <= 12'h86f;
        src62 <= 12'hacb;
        src63 <= 12'h4ba;
        src64 <= 12'hf05;
        src65 <= 12'he6f;
        src66 <= 12'ha3b;
        src67 <= 12'h8e9;
        src68 <= 12'ha49;
        src69 <= 12'h196;
        src70 <= 12'h8f7;
        src71 <= 12'ha8;
        src72 <= 12'hbcd;
        src73 <= 12'h7c9;
        src74 <= 12'h3be;
        src75 <= 12'hab2;
        src76 <= 12'h16;
        src77 <= 12'hda2;
        src78 <= 12'h5a6;
        src79 <= 12'hdf7;
        src80 <= 12'he28;
        src81 <= 12'hd0;
        src82 <= 12'h3aa;
        src83 <= 12'h6e9;
        src84 <= 12'hb8c;
        src85 <= 12'hf07;
        src86 <= 12'hccb;
        src87 <= 12'h3ab;
        src88 <= 12'h25c;
        src89 <= 12'hbfa;
        src90 <= 12'h9c3;
        src91 <= 12'head;
        src92 <= 12'h5fc;
        src93 <= 12'hdf8;
        src94 <= 12'hff3;
        src95 <= 12'h670;
        src96 <= 12'h33a;
        src97 <= 12'h5b6;
        src98 <= 12'hd74;
        src99 <= 12'h3d9;
        src100 <= 12'h36f;
        src101 <= 12'hb79;
        src102 <= 12'hda9;
        src103 <= 12'h918;
        src104 <= 12'hb76;
        src105 <= 12'hb48;
        src106 <= 12'h6ce;
        src107 <= 12'hb20;
        src108 <= 12'hda3;
        src109 <= 12'hfe6;
        src110 <= 12'he52;
        src111 <= 12'hc81;
        src112 <= 12'h94a;
        src113 <= 12'h9f8;
        src114 <= 12'h601;
        src115 <= 12'h80;
        src116 <= 12'hcb7;
        src117 <= 12'ha82;
        src118 <= 12'hc6a;
        src119 <= 12'h68c;
        src120 <= 12'hb70;
        src121 <= 12'h50;
        src122 <= 12'h76d;
        src123 <= 12'ha56;
        src124 <= 12'h23e;
        src125 <= 12'h3eb;
        src126 <= 12'h45f;
        src127 <= 12'hb95;
        exp <= 19'h42ce5;
        #1
        src0 <= 12'hbcc;
        src1 <= 12'he66;
        src2 <= 12'h1c1;
        src3 <= 12'h514;
        src4 <= 12'he55;
        src5 <= 12'h251;
        src6 <= 12'h1ba;
        src7 <= 12'h73f;
        src8 <= 12'hda0;
        src9 <= 12'hfdb;
        src10 <= 12'h27e;
        src11 <= 12'h1cc;
        src12 <= 12'h80a;
        src13 <= 12'h334;
        src14 <= 12'hd8b;
        src15 <= 12'h6a8;
        src16 <= 12'h9c2;
        src17 <= 12'h7e1;
        src18 <= 12'h807;
        src19 <= 12'hb1d;
        src20 <= 12'h23b;
        src21 <= 12'h9b4;
        src22 <= 12'hcdf;
        src23 <= 12'h644;
        src24 <= 12'h475;
        src25 <= 12'hb3f;
        src26 <= 12'h2d3;
        src27 <= 12'ha5c;
        src28 <= 12'hd3d;
        src29 <= 12'h702;
        src30 <= 12'h19d;
        src31 <= 12'h8fc;
        src32 <= 12'ha9f;
        src33 <= 12'hc58;
        src34 <= 12'hd02;
        src35 <= 12'h89f;
        src36 <= 12'h46c;
        src37 <= 12'h80d;
        src38 <= 12'h691;
        src39 <= 12'ha8a;
        src40 <= 12'hd20;
        src41 <= 12'hbf7;
        src42 <= 12'h396;
        src43 <= 12'hfb7;
        src44 <= 12'habe;
        src45 <= 12'h9c9;
        src46 <= 12'hd0f;
        src47 <= 12'hd19;
        src48 <= 12'hb18;
        src49 <= 12'h8be;
        src50 <= 12'hf9b;
        src51 <= 12'he1b;
        src52 <= 12'h37b;
        src53 <= 12'h6de;
        src54 <= 12'h76a;
        src55 <= 12'hfa;
        src56 <= 12'hfe;
        src57 <= 12'hf8;
        src58 <= 12'h52b;
        src59 <= 12'h52;
        src60 <= 12'had6;
        src61 <= 12'heb2;
        src62 <= 12'hd9b;
        src63 <= 12'hf72;
        src64 <= 12'he9d;
        src65 <= 12'he86;
        src66 <= 12'he72;
        src67 <= 12'he37;
        src68 <= 12'h7cc;
        src69 <= 12'hd32;
        src70 <= 12'hbaa;
        src71 <= 12'h934;
        src72 <= 12'hff9;
        src73 <= 12'he83;
        src74 <= 12'h67a;
        src75 <= 12'hfaa;
        src76 <= 12'hcc8;
        src77 <= 12'h273;
        src78 <= 12'h9b4;
        src79 <= 12'h744;
        src80 <= 12'h3fa;
        src81 <= 12'ha4a;
        src82 <= 12'hc5e;
        src83 <= 12'h6d5;
        src84 <= 12'hbaa;
        src85 <= 12'h771;
        src86 <= 12'he2e;
        src87 <= 12'h232;
        src88 <= 12'hf6c;
        src89 <= 12'h15e;
        src90 <= 12'hfa7;
        src91 <= 12'hb97;
        src92 <= 12'h965;
        src93 <= 12'hea8;
        src94 <= 12'h584;
        src95 <= 12'hfc0;
        src96 <= 12'h46d;
        src97 <= 12'h7f1;
        src98 <= 12'hf45;
        src99 <= 12'h41e;
        src100 <= 12'h4ab;
        src101 <= 12'h57e;
        src102 <= 12'h884;
        src103 <= 12'h330;
        src104 <= 12'hfd6;
        src105 <= 12'h2bc;
        src106 <= 12'h6b6;
        src107 <= 12'h8b6;
        src108 <= 12'hc22;
        src109 <= 12'hc7a;
        src110 <= 12'h15d;
        src111 <= 12'h87e;
        src112 <= 12'h994;
        src113 <= 12'h9c2;
        src114 <= 12'hc81;
        src115 <= 12'hded;
        src116 <= 12'hd59;
        src117 <= 12'h932;
        src118 <= 12'hcd5;
        src119 <= 12'h2a5;
        src120 <= 12'h1ef;
        src121 <= 12'h587;
        src122 <= 12'h4b;
        src123 <= 12'h202;
        src124 <= 12'h45d;
        src125 <= 12'hda;
        src126 <= 12'he34;
        src127 <= 12'ha14;
        exp <= 19'h46ee4;
        #1
        src0 <= 12'h9f0;
        src1 <= 12'h2b9;
        src2 <= 12'h989;
        src3 <= 12'hc60;
        src4 <= 12'h5c6;
        src5 <= 12'h1d7;
        src6 <= 12'he02;
        src7 <= 12'he92;
        src8 <= 12'hb3f;
        src9 <= 12'h647;
        src10 <= 12'h587;
        src11 <= 12'h9c8;
        src12 <= 12'h9f7;
        src13 <= 12'h505;
        src14 <= 12'hd42;
        src15 <= 12'h3c;
        src16 <= 12'h872;
        src17 <= 12'h3b2;
        src18 <= 12'h433;
        src19 <= 12'h821;
        src20 <= 12'h30e;
        src21 <= 12'hf5a;
        src22 <= 12'hc0e;
        src23 <= 12'ha4d;
        src24 <= 12'h9ac;
        src25 <= 12'h2ea;
        src26 <= 12'hc68;
        src27 <= 12'h88a;
        src28 <= 12'hfc5;
        src29 <= 12'h7fc;
        src30 <= 12'h6e6;
        src31 <= 12'h579;
        src32 <= 12'h3bb;
        src33 <= 12'h2a1;
        src34 <= 12'h4fe;
        src35 <= 12'h76c;
        src36 <= 12'h741;
        src37 <= 12'h7b6;
        src38 <= 12'h2a7;
        src39 <= 12'h810;
        src40 <= 12'he0f;
        src41 <= 12'h798;
        src42 <= 12'hf54;
        src43 <= 12'ha96;
        src44 <= 12'ha03;
        src45 <= 12'heb0;
        src46 <= 12'h881;
        src47 <= 12'h8ab;
        src48 <= 12'h77;
        src49 <= 12'hdb1;
        src50 <= 12'h8b5;
        src51 <= 12'h115;
        src52 <= 12'h816;
        src53 <= 12'h59b;
        src54 <= 12'he5d;
        src55 <= 12'hea6;
        src56 <= 12'h784;
        src57 <= 12'hcdf;
        src58 <= 12'h43e;
        src59 <= 12'hcd5;
        src60 <= 12'hb48;
        src61 <= 12'hdd3;
        src62 <= 12'h544;
        src63 <= 12'h488;
        src64 <= 12'hb91;
        src65 <= 12'hb26;
        src66 <= 12'h4b0;
        src67 <= 12'h9aa;
        src68 <= 12'h66b;
        src69 <= 12'h556;
        src70 <= 12'h9f5;
        src71 <= 12'hbcc;
        src72 <= 12'hee0;
        src73 <= 12'hf86;
        src74 <= 12'hd1a;
        src75 <= 12'h60c;
        src76 <= 12'h585;
        src77 <= 12'hb36;
        src78 <= 12'ha19;
        src79 <= 12'hd33;
        src80 <= 12'h261;
        src81 <= 12'hbf9;
        src82 <= 12'h8ec;
        src83 <= 12'hfea;
        src84 <= 12'h985;
        src85 <= 12'hbca;
        src86 <= 12'hf66;
        src87 <= 12'h97;
        src88 <= 12'h3a4;
        src89 <= 12'h97e;
        src90 <= 12'h6a7;
        src91 <= 12'h472;
        src92 <= 12'h510;
        src93 <= 12'hfe3;
        src94 <= 12'hc9a;
        src95 <= 12'h17c;
        src96 <= 12'h4d6;
        src97 <= 12'h8e7;
        src98 <= 12'hf17;
        src99 <= 12'h3ce;
        src100 <= 12'h240;
        src101 <= 12'h3b;
        src102 <= 12'h504;
        src103 <= 12'hec4;
        src104 <= 12'h701;
        src105 <= 12'h9d9;
        src106 <= 12'h5e3;
        src107 <= 12'h3c6;
        src108 <= 12'hdc9;
        src109 <= 12'h62c;
        src110 <= 12'h85b;
        src111 <= 12'h24;
        src112 <= 12'h24c;
        src113 <= 12'h24e;
        src114 <= 12'h9bd;
        src115 <= 12'hc5b;
        src116 <= 12'h6fe;
        src117 <= 12'h532;
        src118 <= 12'h68f;
        src119 <= 12'hd7d;
        src120 <= 12'h672;
        src121 <= 12'h8b4;
        src122 <= 12'h35f;
        src123 <= 12'h2b7;
        src124 <= 12'ha57;
        src125 <= 12'h17c;
        src126 <= 12'h1e2;
        src127 <= 12'hc0e;
        exp <= 19'h41b8b;
        #1
        src0 <= 12'h5d5;
        src1 <= 12'h6c3;
        src2 <= 12'hed7;
        src3 <= 12'heae;
        src4 <= 12'hf3d;
        src5 <= 12'h4b7;
        src6 <= 12'hff2;
        src7 <= 12'hf54;
        src8 <= 12'h62c;
        src9 <= 12'hcb;
        src10 <= 12'h1dd;
        src11 <= 12'h32a;
        src12 <= 12'h4d;
        src13 <= 12'h297;
        src14 <= 12'h772;
        src15 <= 12'h105;
        src16 <= 12'h1ea;
        src17 <= 12'h6f1;
        src18 <= 12'hafc;
        src19 <= 12'h48c;
        src20 <= 12'h7f6;
        src21 <= 12'h202;
        src22 <= 12'h237;
        src23 <= 12'h6bb;
        src24 <= 12'h43e;
        src25 <= 12'hc50;
        src26 <= 12'h56e;
        src27 <= 12'h5a;
        src28 <= 12'h301;
        src29 <= 12'h160;
        src30 <= 12'h9a5;
        src31 <= 12'h8ad;
        src32 <= 12'h7a9;
        src33 <= 12'ha63;
        src34 <= 12'hacf;
        src35 <= 12'h669;
        src36 <= 12'h228;
        src37 <= 12'hebb;
        src38 <= 12'h6e2;
        src39 <= 12'h5ea;
        src40 <= 12'hc19;
        src41 <= 12'h2f6;
        src42 <= 12'h87c;
        src43 <= 12'hd16;
        src44 <= 12'h239;
        src45 <= 12'hd10;
        src46 <= 12'h53;
        src47 <= 12'h6d3;
        src48 <= 12'hcc9;
        src49 <= 12'had5;
        src50 <= 12'h43d;
        src51 <= 12'hb89;
        src52 <= 12'hb3c;
        src53 <= 12'h685;
        src54 <= 12'hfe2;
        src55 <= 12'h288;
        src56 <= 12'h348;
        src57 <= 12'hbbf;
        src58 <= 12'hb1f;
        src59 <= 12'hb40;
        src60 <= 12'h686;
        src61 <= 12'h729;
        src62 <= 12'h5d2;
        src63 <= 12'hf11;
        src64 <= 12'haa8;
        src65 <= 12'hb77;
        src66 <= 12'h7c0;
        src67 <= 12'h867;
        src68 <= 12'h7a4;
        src69 <= 12'h19a;
        src70 <= 12'ha49;
        src71 <= 12'h4bf;
        src72 <= 12'h84c;
        src73 <= 12'h2be;
        src74 <= 12'h752;
        src75 <= 12'h3c8;
        src76 <= 12'h894;
        src77 <= 12'h956;
        src78 <= 12'hd05;
        src79 <= 12'h3da;
        src80 <= 12'h6c5;
        src81 <= 12'hdf7;
        src82 <= 12'h8c2;
        src83 <= 12'h130;
        src84 <= 12'hf3b;
        src85 <= 12'ha48;
        src86 <= 12'h183;
        src87 <= 12'h92;
        src88 <= 12'haad;
        src89 <= 12'h37;
        src90 <= 12'h547;
        src91 <= 12'h63f;
        src92 <= 12'h7da;
        src93 <= 12'h8c7;
        src94 <= 12'h378;
        src95 <= 12'hed9;
        src96 <= 12'hd65;
        src97 <= 12'hc76;
        src98 <= 12'h4f5;
        src99 <= 12'h98a;
        src100 <= 12'h3f8;
        src101 <= 12'h60e;
        src102 <= 12'hbcd;
        src103 <= 12'hb22;
        src104 <= 12'h30;
        src105 <= 12'hdf9;
        src106 <= 12'h112;
        src107 <= 12'h3c5;
        src108 <= 12'hd5;
        src109 <= 12'hcb8;
        src110 <= 12'hd11;
        src111 <= 12'h670;
        src112 <= 12'h916;
        src113 <= 12'h313;
        src114 <= 12'h803;
        src115 <= 12'hbb0;
        src116 <= 12'h26b;
        src117 <= 12'hc62;
        src118 <= 12'hcf;
        src119 <= 12'h399;
        src120 <= 12'h447;
        src121 <= 12'hf5a;
        src122 <= 12'h178;
        src123 <= 12'h93e;
        src124 <= 12'h63f;
        src125 <= 12'hfc3;
        src126 <= 12'hdcc;
        src127 <= 12'hf6b;
        exp <= 19'h3c9a9;
        #1
        $finish;
    end
endmodule

