module testbench();
    reg [22:0] src0;
    reg [22:0] src1;
    reg [22:0] src2;
    reg [22:0] src3;
    reg [22:0] src4;
    reg [22:0] src5;
    reg [22:0] src6;
    reg [22:0] src7;
    reg [22:0] src8;
    reg [22:0] src9;
    reg [22:0] src10;
    reg [22:0] src11;
    reg [22:0] src12;
    reg [22:0] src13;
    reg [22:0] src14;
    reg [22:0] src15;
    reg [22:0] src16;
    reg [22:0] src17;
    reg [22:0] src18;
    reg [22:0] src19;
    reg [22:0] src20;
    reg [22:0] src21;
    reg [22:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9267ec75ffab6a354605c8abda6eaa01401962b6aba6d8dc134e4ff3d463528a846bf8acd1bfaf7762bcb50ac1fcdd85a09078516ccbc05f6524f02cc6b7372d8216;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f5e6347d25a393882f72d80ae6aec924faf3ee978aa3e25b1938ac703133213b1e69b2489a1c7a18d2c09fe7d1ea079e47300d7f04ea5a29315ea89f800cc815918;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d03f0f666abaf510efc045cceeb67ed9439641148e8c7866a939d91c9943579f4dbd1954e78157798cb20fceb5069669d77021d8d019f731365712fe0d8c50d8e015;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd715d672aab2f62b43071434c1b3312a875d2318eaacf8219b3581dcf9f0314669c3eac4f90535e01cd90b4fd6be0c2e0e36ec6d041907119a3ef0a0c3a54c88e78c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1f8cdb5592cf43f1331dbfb20b565c0496ee4ee8e25c4236625a5cad974a11b91ece71d82d84451df7f9aeaf29987597939c690905aeb26d2e7272abe9e92ce24df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df182849528884aaf14773ef5fe8b0b5783d389b28253cc64929b756a1b91a0a89b1fff42a2d489fdfb4eda1f4ad84ed9822dc121efdc30c12506e22486e68e2b9c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16bf7c22251db05064af270e22761c1c2fa69075bac310d55470ea5442a822725a6dba0ccce7356ce3e128e7ee73d55d6da96129afda57fd70b4c3d1154cedc7a11f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfa8709f3a0b4e0554a32278d6ae9212013bff2a06bd5e3379f0052ece420c868ff83acf8396b0295a1b61ca52785c92b653676ab30371e8547c827777f854ddbedd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bd89fa52da1b5d843f2165e3062e1bf2ce473c624ef2db5a32c87dca7eafe11c8e7e63c4a2ac79d810265890534992594b23de740dafb475be47f4cc91cdeb0cbe0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4563cfca173fd5b4614833656de2b6907328f5a9317f7e98521f347845fab2a69463e185095c28ee9032b8df66d6d45c8cb931301096ee9a052a27e59025b7761dd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haaef2251cd9363c6284aaf3a5802420e245efd6b4ad8de057beaaeafbbbaf68219805f36c1f4cfeca69f12fa2b2951b0186ab0b96f2b7ee2f4e68d1c7b50367c8bff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5bfdcb1647ab3eb99dc9e2d983bc0697c3624715f03455f8344425668de25cde27c0ea0167bc866cc3250e21ebc04e34eefe5880c35ddc972ba79c9c5b69f8b487b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h201119f37927cc1ea82849b024327d18f52a0eaf7235b751fc215dc7d936ed12a042aa8987b198eb5f36f793a62ef7d043ac530c6b1a074e233126a2e81483e5b56e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa42607bfcf83d660d9b197afe5cfce8f5b30da2e9d6eec078c55d1e55272dad1ffecb96086a75e14849e95e9ab9129b9069944e6a3bcf63fb67fc9a736b13c3b712;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46ea67ca165ec46f5790539e48adfdc47366e9f5d212cd9db9e7576208bb6b651d45977379399596efa7a138f6601a98d5621695fe95ee9dab9ce952c8d0dc23c6fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35740243b52f73830db1d948c995c3aeb719c9a337eec6d5117a495b466e889f95516b597689a87e7ed1cf33d27340a515b1aecea39e0c89da8431499b9c8af22b1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac150491fa75f9a33067b4405b17f4e7715e2d8f6788755d46bd59b55415b7c341dfa87bcf4dec4a8ab0591bcd44c93c7106d02a39193397bdb9cbe5bfef95c924c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ca4114f75c7122e2c11d506dd6b2ddca62e92b2291facecd09e1b92084ca2fa57fa7ca84862b97ea64d769d277dc3247356b23be7f9e0ccb3c2d376264d8b63c256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efa11eb7bf533e8a9ab17c855ed1732e77fdc454d2b299b20ddd5ab49a3559b7d91b6028ec4550cbb76c687043d923bd9d600fd1751914abd77e3bc6473775e6ded0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf31200187bf605906254fe763a50eddb4cd0dce2608d62d15e9c08de7bf9ca777b30d2624fb2ba879b7d6865b9b09a7843b9cb6b35134ad299c90bfbb1266d8a92fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbb6d267c20b4518df851a698564a2e9a7ca51b123fb1f22993ba696e3ed8424a6600cbff4875ee15c9c3a0197db34fc65fb28953dc0e3efbaf021e15a5b1c727c3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h827722fd2b8573ea7bd68ef96db45f2d4658b13d3eb0cee8f4fc1809395f7d9accaea82d784d4b9fdbbde8e1b29d6abe7bd079a473cc03cbe8a0cabfcc3205f536b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2900581fabeeea80f1f891fb6dc2c21bc4d1523a44dd244444ac64eeeb7c6063ffeac3436541d72ac03f21d3bce707e50c4def3eac985851048ff9605f808ad7ee86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175f337d787c5be09ce28f9822130749fbc9be97bc264a1c062dac5b5c250e89a994a80c9bf7167d030234d4f2dc19968cb0a87b4a6947510483751717a8c2819b17e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a42a3dfea31db0136392dd9488725a7be168a9e4fa1a7fd6e78429af1a04c5c856c1e8b93d627617252fab70da182af69fc1c87af7e3fc40d6a31aeab2025f17b07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a866cf3d4626a226fb2ece1a9b48adb570983bc7cea2325a36eb66d752558ff0e869386307ece0dc44f08c2f97c07e3f76f8bff41527299d35c2f61b9dd3c76e99b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9a87eb0936bf02df1fc7ee968ab5c3328508948e5aaab8c645dd6ed4a2febec3127f708b03b41d6dbeeab16f01690066105015e81269c4c7a9ca7d806ff971f6bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf0dece2667819099ee8fe58540e8388c34a6f359016d69cbe2033910204b02fd19554645e1f4bd1540a35317c7683464337b1473ba421f35fadc0ad532ece2ce3c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53491b18d3c9df0009f552d8498531f134b8f648e5b37f8313e988edccdd865b0810861442b7365f3571ab6e711269091660a6fed87f233e128ddb9af998ced755da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1abca2b9a14cc88ff39f4883cc5427a1d4093150e1e1795f72d315b17e3eac9b380f6279c5960c3e17615d3581f7ed4c6b7332fe1e4b96e12d0ab9278437c574e392;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd5ae9bca22dfe22f6cf3006704cd543c40a9ae34bfe8f4095a5a3a24f404be0b4f4b708af15c92a091d31b589097cfdbd0a839623b6c22caa30599d1351aa78ba1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b421b0a2b25e8ffef2fa94ec91535d6b89007a9255e3ed419510425595186165bdcef8ace5e7d932409150dd040d4a7559f2a257b2424fa87e411149b0a9b85dfe89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1b641febdb41c86ac37e78e519db209de69b21143bb2906c00d42b0fa774454ed72a739f80f45e20dedf689dbb921dc536c778306cdbd33810548fda053b52b1599;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6c8e80a1ce288e66dd6ba0c256c29ad1bd86c927216ba3f172d5aa90ed677d438ca314c6adffb1a8db84322bcf203d2e832460fd8bb71d8773fa37fd51656224f73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f512497ea7c39051d7f4dbfe40522ed301e37ba476227d85c4419a68911c54ad55ae38c36ed97ff50f97ac92bcc11ea0ab64f55d759e19fd753e2a44aad6fbc15b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0ea04cf8c7bcd43ff4df93c12383c511126da796875abf5f0e28bbc027ff3034cbbf1ac4fd4e8bf853a6d64d91ed1179a12e19ff80545583cbc8057a67c5c7abc56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16398583a5b93cdc4c7abc88d0e0cf4ab28f5ef409794ada195632ca2aaed2009cddb1ac582f30c4edf0e6143e17ced593e65b2cb8f422638b888fc437c5fd2478842;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8d8956092db6a837e1e940f461199929ce29256d4e06d216ca6a2bc6a04b8f0c91fb498aeff627c5a4cc0b5791cf58b89153768bd6a8a5c728466c9dfba77de0e1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba74a8628c6a10d50f5d0deef3a7bdc980d8b6bcabd2a73499347ecb548ca9f88b9e913ab52d81c88645c6e6c909f4d9819ec2c7eabb194eb358d0e8de0e6c7987e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdaeba8cb1365f4e46a256dd0d1f37594dc2c7e5aedf39cd4daa77f3e54102eb2271c12efff397388f88e113c49401158c1a8baf3241ec20d8fdc85cc6d38bdec66d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c2a1edede41061a352cbc5d67fd93670f206213a4e260c84cb44f9590634de1f45c74ecf95672132d7a1a5ac59213f3f06b6df26e0cba80a63deea843677d8c8352;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fdad0bab966e5126562d009a01a804e7d7c34a7aa5aaac3620813ce6dacc5655edce199933abe445b070f6d9f81c761938fdae6975e5056151a8aa3d41a36b6c1db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5815c0a5cab81290df7864df2887040ac70c641bac313aa61c56fb90b6ff5fc8ca95618bb1e16c3ddce318332769a4ef3df86bca99c8cb4c61e96fe56d9d74051a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha71b48e0f8e8ec2e36850b4fbb34e3bf975e52a4dd80fd97e25e6703a152c070fbb6d46f2c5fc0db78a483d48abca514a7621be2b257a633c25215b52536bc868fd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4873d25df5bf3918b3563685326599270f444e2b6c2859da0fdec30f3d8df0d46826a31549d9e495d0db249611628600b79e08017e0f810d3ddb3eb51410e8bb09e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha96dc0b915533b51fd2252faec574d73ef7325af1efe058bfa51b4f3543df2cd84eb29ac6912e9b9dde0556069ea15b56686164f6deea1c7cd15ab35877f4132766;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc80d898620014bdb4ae9c36a01795679bc567d681af16cb2774e249499846d02d9a6da294df8893fab8a615697953d603cdfa874bd2fad94f6f4984e3ec541f7a7cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd7521cabc2d9d955d4ea249765465e25a3761051d4208e704433ac241aa4eb31ce30feef106390c5896fd84bedeb3b763065b3a189868b10c1b7482e4eb52525996;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6006c5b181a20b7a23e657f4f0a4f6f892731e3583791b395de9b07e4c9a727c92c55c17cc393a90388467a077fb43fb0d703261ff05c5b167e7f5a31824ae8e01c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91478af2ce67217419ab58d72c791d481037e4af6f7d67685c2ebf7cca7940e9918fb49341c0b1ffa18159dcb1c65dd7501caa395b09e22bda37b0c2471a36c38315;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3be92788b0a407e1b4cacb9267d26538a9332ba568593a27d6d08456b64084a4d863c72d6bac448f0dd929e9e8c35d70b7d42acfb74d3ed497d4c7226f7a30f794f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed4b4e291381c7248efa3e58e449691a3d27fe2e54bf1dcd3f81ef49aac573a7043a86c9c5929ba370ede7e25d556ba41dd12e24ac52bdf91a4acf5ba8b4d10cc230;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda6d7d25d9d6ee5d68c0b805ec3dfa3e078f595448159c658ba8118d02997394dceae785b2b77e894e10703c259ee6bcdabd41f296f00d54ec914f6beb3e10039d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58e93d3455f61881583f3720a25989f6533811a7f6bc2604dc74a9951626225a4e90492b395715e1f9188aa8b4859dd043007547a90796090abff7d0d1b927b61e00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2bbaf0b2ebac47357cb1c6cd28f841079afa085c38e625a199f6f24bca46d45f60fc4f6af51cb0d9d482832b2e0907a21d5c094dd440a1d227878e657cecd5d31eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h930972e881b859fedd9b405fca890d794c77428642d9ddc3e29f66bb95f30a8738c4e08fddc7e9885d86bab3730a59126966494749f2f929e04f461efb718b5a47cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcf2ffd3e8e09741d03d36f16d917b34a57eb60c0ecf8d9ab860d804f141108da873dfd7eb08b37b7d54581a579817a0f7151ea00f78155710053e486fedcf9a3f1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8814096dbf2c8b9b0866f6314d4fe0c6c318c08600fe995c1f39ba04b8042380e4c805a31d4d619aa7daedf9050279cf202b45a1575eac71bac7a081c4bb67a9b28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe8aa6365ba4cbde9ed078b9e4c14b01b69193c97211f9c575835c69d763eef66ff97cf857090a865bc86f154f20096bdf477e8932be719be72ddaf12e99277005d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1233b40faabeb9d558c7777196da11653abfe591a10b3935d11657bfa66e6fbd25f389d90cd1b34228b38ef7e38fb0c358c7ce110c20914bb5c912142808bc4dafaf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb709858febe527f8ee351d15e2e20ebf6ca379b353bbf8939b4dbe7580031b41306ec7f8044436a26f3b596f2a4ceb4073173ebba8de074e21469a1c104fc6428dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156b245592f186eaf71b4daeb7c18e19ca157ba6233488f5ae6f86e3d213ecaf46af5dc29d0ec0f41491bd702052fc26437370e3ec9b62da95279a38a0c4097e8c8e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc99abab28cc6466e7e1e78a146e76d22d411a847599478f66b0c9e9ca721e88548204e78bbc279df665542030aa1bc6b3c06fa0a7d6699fcd18a7e6b23ffc7109203;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc908d42539f8890939b777320badcdf0adbc3e0e2cbbe92a19ed6a5c736eb76fe8c1e628ef672ed38d1031a3481a93ff7a9d6cbfc20c3754a080a29bd27997a0a13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he50503dadf012ad162f56c013c69cb29cbd5e38bc3fdc7377845c3db7548e3f2d620d371d8f7937267acbbcb748fcf13554d6392ef678bd74c1154ab5b176501b373;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1277ff92e11b06dd3bee8096add12edc3d65a079d15fd9d8f8edbd1f273d0dbcff7d5afda32dcf76b82677d3c891828691b9daea254c81479e9d93ca6044016e19189;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd0950dffe3270338faab06217bd2c8aab27a7ee1b1f2a4fa5e3f5ca095e2c2eacc66b3b87b350c169958851405fb5429d4f1646fba52a7764f695a3631f22af6f02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13aa4437f5bfe7a3fd77af9a0ed687076e42be346f6ea8390b0df379a06ae75486a37f9c06ae8eb5cc1e354ef8a8a041e39da7469d2303733014462f40d9bc47a59d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd5f838e990e730c6f45ae75a82d7f456b2f741de1f041dd44c29fd2d35f02e840d5b4fa9f58f5b3145a57c58b87b466cf3fb75cc09219a6a91c488ba9ed00fb78f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d5345a34286f6cfa705aade2ba52a878d97df291c0acb48bce3b01687ff14a843b044c45fe8829070b3b78ffe34ffad9f9b1bf489db4aab254d7de15f8aa6bba9b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d72970268befed55058db4e83a4c654b83d5fd3a98f3f254d5876dad3a2226338b024583a123b7a5fcdc5fd0337234233040695053bb99c0505722535578dda00a84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d41842c293bfa99f8ad77b40614ef2411457e411b77a3eb9626f41ea5e472075466c3acc9ebf539093c36de7598572f72f7706368ea231cb82d1e442e94c0612f69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129684a5bf1e2f734d97d88e1f072cff6a756f07beed6702eb04f4c95989d239355d6fed859eec825eb1936c074d24d2149036c0a13d592c0b6185c08d571a65a6287;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73e5516f48a2f80847c6b85651eb965f0485b22439240012bb2bff901573d62819f4884d1ba87d87a97547e7ceadbf685341ecaf5c3f54cb31f8387406e56884322a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f27ff7737c19e68d9a4a1aab3d21d169169384f91c696608af668582963f231fcc858d25b7771fd860ba008d28a87161c1f44687a37348eddfb954d7237b1f93a54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133476accbfc9b5bbe4bd9b4a47aa98e381a04d61a4ac25d2b4240f8a2562314b6359e6e857d413fe49d1fcec17f6cd7bf61d8a489f9c1eff0a4c20d1cee7a7529c02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0fcb8d3e1f0c4c647c3897c67679ef17a548ef5cb14a212fc00109d0b0105bebf11826e4b57b6c9ddf7bb48425d62195cebc2daabcfe5c72f2126513b33d05d59ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fc1a2e7f80b55536662ce7576101589c573483040515409f295c89b000a99ee26a37622d932e4ebc0865e5ba9a59812aca027f5a0ebdc21217b5ef363b4b774ce58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138658cd488eff66692409c089b3ab514e3e3da673939f679b4871ce00a1ccc2414d5b1b0fb8bb951e4a3816d41a083fcfa5302338c45d416702f54f680533db8a542;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf826f5cce5eebde11053d27c87939c5b66f026a7d1a88f688cdd70abdb734aa34652b5be10197e1fda391c0fdd3a68cacc0835ef5aa9de79b495f3f8d3e253e6cc4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16810c4bdcf73c62925e41b7e2385b75fb24591b4b00ef077b9c36bf01a81a608263b8f5ab51f7f919b40b9707781e4f6c754cdfacd79fbf464e275837f1324fc42c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3b7a66dd58b35f9b19efff9b40483cc7344022f0c7fdf9b5d53e3a7b0037ff2dddc01e9df09ea5d0eb0138c853bb5c62bac3d414604218383d3e21059b63d50e4c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af03139c54f848fe5a1933dfd4e74ea9b7a645cdb4a164d5044806e9370bbf60e32db304e816fe44d8b6d538c53703630cc927a5051aad96e709d46ffa43774726b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50498a5196e5e78f52e659484f881cf1f66ef2d1325bc725b40c4ee44a547124d20e4fdd5960354ac85eb394a022b29e220280d9a85cc84df542bf37b177612dda0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5a900504e5eed506e7c9e2c1a64115d75b1db60747367fcb8c29156dd25ec214ff6823ef9ca3167782215a8d92f8abf82cd42497369745d5d4977d22b0519cb939;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffd266aa988206f73a64dbf5a97c5c3164ee61a55f832016c893268a3593cc3cac3e775cde87402ab1a8de52aeb3af86bb9c82f2f194da575fc659f01e49edd69e81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128d5e0e49a221663a2de03c29c2a9505d51b03bda4739fc06da7d478676aee4e6dd87b780b19cd977dc474db0839c9ef5b723239b348cad9c348319f43cd7b3ef654;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha388a267b2376b405dc56ed543d4c5d69e92188381a5447f2b17b7ad6193084db70394ac3a37b3a279ce98690174653023f32877752d01e33d9b5f6319dcb998fc9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d297215264f8c3280577d39927a258103c83c253790614d16d55368ff7c6348b3e6838d85ac0b0c9531cd862ee4bbc5a401bb70f95eb9fcb274ca45edcb69d945813;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4b399da6e26990cb4ffbb210bcef19fa6f2c2267c39a9efa4ccd53475f71c356d549523b88d7658b8608457c02a18fc1aa37de14d5c13fb4813524dbc961bc44ce6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f8d42e27ecbcdc912a1a05cd66dd0499afdb1d23b4ee09caac7d9aaa3d2c9abeb8df1cfdcd806b44f92f36634399f99c9e8a52b481106780b0af3f5abddaa5757c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7aa7290a2b48ea66ee9e19c6f448f068332786d409c5b91b40dd8a434ad68285a266737bdb46a0f38513cd7da71f202f7c8ef2b7464070365900dc2d66bb0a05f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae9cb99a17fee366774a7a656fb04f0394266595fecd9f952cf14de02fd54b6c02967b77ad11798dc3d01a3e444f678c041a81d892caf44f0a8b970cda7aac457925;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fe9374688910d15e791ab6bd06b645250070ba6e9e23a50c3c1d4922551b09719aa1da956de92904b4a56acc4331f9fe5679eecdba1855e9b5c153d766f9631c222;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61e501d026613ced33b4baf8b8872c8a79ffed4a4ae0b2dc099b597edb539ccc57324e388abc31e4dfc5a30e35b0c81ea44bcc535190500e562fb8450e56b4d357a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17916e5a9241561dd74923483d4451c761f5afb275e4434299c6d8fb6f87ce3ebf391fa292a078ebce7919a4ab5aa1b349254af7908314ffcbabc3ae22277fc5a68a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed0c7de48d4aa0a28dfbb3b1040d3f5ef69007c77becbb297a82a06133dbfc932511ef738f3e0dd8f97443e1e12290884dac739ac79225bf4648e56e467bb85d588d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ccf32078d3da93a8781d569945c37ab5fb68025537abf9cab30f2962f61e720b089b6fd19cdd93a5f321c6189a040bbc856e60d8846641fd3119403107b45b742c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h403ae5b20f318a6422f43abc5a9e986fc2477d5c559d9fb1d637944b21ba46df0a3c04d11b4416c6c2bd532f0ccabeeb5689fad67a6a3d1a8a59585672596011e8f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100f382e6aec06e77d4b9a3333a45e84ed52e61133a1d85b894931e7341042cf23f08efb94302b08c30c43527c958dbe7f942cdfdf7a007511464340e2890b387b584;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb7df5e68b1d0f9d596faf5c5f1f293ab4079c424954a8a088161fbb628935521e95949b2c68ba3e63046a56fd5abfcaf56058081b346e47290c4b8c037782c89d0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd454fa43ed824128d46f42311d685fc40406f713dcd6f37a71665512d6396d0332fc12d1e4f095d7bcdb891708315de92f4db4f226446f344e86dfe6251d614bb2e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he63ce8b2f764a574ca3c433eebc7d79c96e734b32d3215bfef6b8ecb1e65ae5167845265ce6eee9832a08f69e36a5be1849b515e6755f363a5652f0ea819b8929b34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104550ec5faf1a0639bbbebf0575cfe3f3ffaf0df1b8ba06e62d7fd5e9a923e23400e1ca89463299332fbbe41a4b9904f8167aacd7c39aa1679c8d1659c586462dd98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1047299b7a4aaa9a9d2da1ab23f7960e29ac6dfd1454ceb576c06b3c789769a337db7c1efd66534fca32ef750045da3377d379b5d750f650141c65d55a4916c8f3f5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf48eeccf1e5be853e5d2018c99525431fdbcdebf3aa76c63fd8b624f5e8634a1376dd01172997eeff931bc0011f4e8d0b3840ec6b071c628949a7cc59780e9c854c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93c302061be1b45bcc616e2119ab4b9ab1e470547dd4d85040d1245fed7d957bbec4fb88fc55e7d3917342bceb8ef936f4e70f3052f60a8016e35ed6c345b68e147c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c516a597e7c9d159ae7c0b2bc1dc713b31aa0806a2b39fa922a8c16bb65b16abaf04c3756c956abadaf0c579313c44c87c1f495cd2d721b840edb3b30fdd4ff853a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h600b4f11c7cb44aec551d59af4d80c76f45bc9f4531d54f99809de850d47b8913da59a19755be1639cdc6671cecb33a59f1b7ea149cb154af0980e5553371a82cc36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7a2dd483bb10968cf3c0e2c18837f6c88800879b0c548df2f57f529d99928fc2df9638c9f763381ff7d28953496a5d1dd5780308d1e1e4412ad4a03daf28bb934cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2be49933c6211ad5e8f780436bca41c1d8c3d642ff5394ecddbf68e760898add187855daf3e7c8a4eee6410e33a56dd4ab35a46b1c78a4cbae9eca2c0222ebfbcea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db897374f72d5ffb006939edf10c1a9e56f6ca57a612df7a96fb4f7ebe6d4f749b00ba5eeef0d4fd4e9863d7e8be2eb34fe581eff256f48e677cac8f07ca67985fb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a795c34d9a939d1040ec9cbff51d6088c697ea403569a620f73b68b29e6a4f53958856d831e69cb7668fbf6d213e5121ce41b52a6e933be5895bd996d687bd691137;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15dde47b8339c17c22a95d57c2c8de8fb72fad8f07ee6692590f7108b076510fd685f73d859f987ef331c6d4c39964e30191dae784e5535dbf41ff58fab04c8b5d949;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3886cc3820fc6706eb7d75b88bf3a0574d080b3b0cb4ef3977637c8696572784514d6ff281719bc197ae9205c7345e3a14dd97c1ee4361a8404e44b45521cd709ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d018367e1a86b3c34f4b33020121aacfd6250d2a8577793be3e2d468515bdea3bdb5650aa3ffb203eac0854fc724d1787672aff8d7a05d28993577dc3a532f25191;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100ae10be77622fb1dc90159cdef462645f3077c57eb1f56bcd65ba459509191a3a3214e7e2ca575c188786ac56e7acb565d95bbaa8e0d7b5a7399da1ea5314adfb2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fc084cc7d09a3c24b20150fa94d9ccff6d0716aa7c796a48135566d4f68e0ad226d1ae1cc486bba1e11356d0eb4f0cdd10337080b1bf62b7023d600bd8f471c8002;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b91c14a59b38aca69e9f1d6a33e143069246dffc9c1fc0ec13ea91675e406d2f9455c104f8bab9a2913ad06b8afff6baeac219b52783735ed2c1278bbea765d7ba1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1220f49c2d4af03d77cd9f8ec8c1b074d4b88ee7ea975ea0837cd36b4128a2ca355c83b9e64b1b8960961299b41a1c695f4bfd8aecaf502a498516a8c938db1b38f72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h967018f2d5059a3c828db6cd876d0a478deaa4811baccec3823f6efdc9beab477ecc1d1e68125813366afd6f5e6532ecaf2de2f0da4cce7c49abe1a729aaec8703ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h902c44523f6e16ef539ed06e7b438d1f93a86d3b00d3a3314f441c412fc0dfdf610dd2d3859e6f6780f82d0827140828553b7c896e5840b8cffd9b9d0e92621e5a33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8d9a65cf23f849d5beb6b82f776c516bcc40c22348f73d2290ee8da94be3c517e69bf8461a334312c7dfe1e83e6cefc5c8b472ed11ed6f6f643fefd229b23886c3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9c1643227877998eaad581a58708a1489a5764f658caa3086ed36be3b81aad7cfedd20481ebd6880ee9bd5e3291b3222197108077af7ffc0dec4055ab12cfeda3f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3fb85f5cd0e7418be1dcbce993b281423916696ae9dc38855b7c07cdfc4bb5b5d0aaecb091a6457b963f9094e012b5b8a60b53e0e666a602869a51e4dca7ffbfa2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1168cb9bedd080a0bb050cebd1390bfd66e727b54d0730446402e5dbd23e9ce1e00b516f9dfb2a8540a868e994274524e44a0fd3c9b049963e83d80f615e6fdf219d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9e9c106cf659d6f5c88a5e0252673460e7517decd37d50b4c22727d1d0b068c094722ff27d79b27b8affb94c13adadc8e3331b42f36438d92359a37fb6f4f8b1ab0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f4a0392250e3fec3bb783bf497be57e0fb5df821db4c0735c441974ce0a0274b8b66658b6fd4c651a2a90305ecd6b56f5d663d9ff6bd786ade836d1ccce5707b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2933df739abae36b65ad6ceb3ec3d70c60bcf960f354544f317c95611d2f2bcc594def126a96b56ed7d9ab2ba6242eb8cb496c3b025bebe782b27687f29c3fe0de9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffa00bb33c7320d502a82e7051a23f3206d24dd924d0ab4b1ab6d777e53710583de519f1ee0ff9522de6e7988a7d8be01262dbd3dde717206c00d24b072c114ffc6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6c8ca2f39a9aeed9ddef78947e58de1ca7bcc765af7d20de72818e52298e00f0b191bfb80b7024853ff23fea3095dc3fd29a9ecedf0f416e3f82737f37a9c2e7114;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6085d80ac82e6c1aaaa2a3547be506becfa60f6c3305e3a0ab30e1635f5b344b0dacc55105c1f4304242bdfda8011814be7034eab6fab998476ec2c00d8d52fdf45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45f13f1489ebc88c6d063de4029f578c45f3c91f45ad4ff122058d495ad1cc43fcc21eca3d1148abe8b681869c26a2972235b625a02cf3f9756fe0a580ffdbe8f27b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6132ddc896fd830f8206ed219e7b3fe16564a32d47db44760831db06b1644b0d6c9cf4d48d745f14f5bbdab8b13f934dd1c1cdf8c8a84ff4cc646ab309bcf43910c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb197e714b70beaf24534a21ce59e64f5103e89db596f65361d9059e0b8791fa04e98e7f9d6061f460540a78554f204aab58f8de459a3733cc628c1b02834ba681ef5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a3cb8bef4013322696bae305b8753ad55900dbb196eef7ea4e505f6379d95afabbee7a00c5d633e556ea76f68a8ca0746051569fa156376186ffa0b5bd3b93adce5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bccbcfd2098b9fc4e579ca4922b24ca919facde80f5e98c71750ecc8410c01cddeb2fc5d2633fd21c97e45f264fbb9bcfd3cf2c60ef87a00783173feb107af4233e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a6cd60e468dda751ad4826b1c8232e570433fb992a85b716419952efa0b26e6c858cb616fda7cde47497d73a6e04c5218da4f0d2e8fed145f44d64975f2a4808810;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87284034b4d8f728b63791fa6091853aa005afba546903a4659650b4a73646a465eb944ca56d57e807437d2fac9d4fa0d4f571fb6ebcfe8e989ed0563ed994c97be2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15eb30dd381d84b9f6a12c1b7c658e8f2b10f14c23ac96481ee3f13d06709b3b32ac50697717d259c318b6c98d7440def48c0dcf37e1f1e761ba1514438629811896c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d8d7404fc3027ca483793978a9b705a67ff5cef940ec44d0182a388a8e8c01ccab070a535fdf0554aaafd959bbfd3bbfed3b0524c58eefb9a0f9922b2874891a51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfeb172541456dd67c027c291341f45b5874ead458b3d57fdafc106895474f3cb52c61276bebc92149d5a00536d2fa6059dfa3fa1baa93f5b68d7176c452ad68c68bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff3b6438b390755a41ab241d2205f4cc8311bf0ece4cb79159136d6afba58a99c21046e98446130787a0f58adaac8c423f7d7b9242414c1c12f07a20aedf508a77c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b5b8fd474f2405cd0ba68b15d3add459d75e7a1f0aa4f53a504ed30ba27ce191b6a4f88d662ed821d4954a5f9148711a92fd64bb912c8dcc6fa9bd35c4ca5268c16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5ce4ecc64f8e2f74978096d7efbdd07f94e8de79fa5ba8806eddaacdedd045a5db745d53983b005397b5785a493de13757c70cc1291d667d5822f857f4a49077843;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h825e0f8ceaf12920450ed9df22bc9edf3a941ae11bb249034bd9461919bdd57642f21659e8a465b03db3df3881b66b375b98a77163ab460e4676d91b38ccf6a13546;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b8cac8a5ee55d073a16703ba236f31252463194b66dec758aa6a0a73383ea1893e524fe3f21d9ccaf4df3830ff8ca0cfd7ab1a90d3cbd0959f8a8684c6e3cedd8dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111857240acba7b05f1b2a76e29edb2b76a7106d1a829d19b847f6fba323807b3736125474bdb8c0022517aa26d649a56d1541f8cb0b4f4925d51132aef28eeca3e4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3acab8a1b4c070e45276ea73af42d2778d35c937cf94c86289a28be07a1d688e3237ead6f8943c7495e13663990e3e50258a655ee1c092d9b08da33c34670690f04e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec65a5eef5497209b834ad53fa4cd3d743cbb0d23a65b92f9e252ce423a009442e189c4700af02f7cc1e3b30de2c8eb2dc8e98f9d0c5b7bddb5025b37f6352b6a043;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f78aaa9534bd8f9e78c8828fad1545f0a8458c90c0f31f602d15a2f3ada317910c29b55d50df10e3e8b33532c0c5d8be98702218c80095f696c43cdb361615b9c80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109eb99f5309cb05c991751b9bf007cef7ffd27d22d6c3998b105068bbdb2cbee9b31b6efd1ff7a2216d7579f75823b8151ce321d86c7dcdd282fe43980a53b7f983;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7435abf495f3d92726b41ce876a21aeac7e60743e4ad2135f684081b8e2a58b52bfe7399173c0f477c212b4f2544fcfdced2210b68ac9ef6f5606e2f795874bf8662;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a0b4d88c85e54f5a40b0907d9ff4aea9ba09c76b7a1df2a7697cf8e2519522016e10d0aeb2adc021c0a9f7de4d5a9710833bba83bf3c88b3d867397678681b5a09c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106d454a125791141109f5423ece3ccdea45e081223f25be25a0599e4ca8ba18d714db74c54c4c57ebedad0346021454605c462706e61b922e964cb351d266afb5a98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f0ade5267041e0e09fb2ecc0c2803d00bf6eaf34f261f0c172c1578d3995922236978de6611de5bac34786a4ca40b2c8e7beb37a8349b713aae7d71e89d578139a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184fa4ef1a380ab628aee505aacac842b87c1a4acc85d05e24ad9e6683954d6fb928a71916ea9a801c7dd803a743ce299b3a2ab93ee3caca77965d70a9463a8202d0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee39d7f8c134c692f5fe638590efaa76643225b1ca6be0350e0935807b723f049e8784f64ce6f6b8da41abd7da118727cd3232e890bd3c2074a7bc8cbeffb93e4ab2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bc93ee67e2ead91906234b55bde6a896bc4a48e4457fccf612feab73c2407f31b9865e53f17c7cf3d3f232b412c6adb6c6c5e4c19b418f4bf667ae727a15a2e175a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c7f9526e49c3e369ca7e9e0047924718bcdcb520ee8c0787fcc361667ceca355c3f431107551076f6bde83eb920ccdfdfb421cdd2315739ec9a2d32ac7abed862be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1133e0273c6c4ab5a57f4032d536ca5e6835ea4b38ebc9709d570ff849cbb72900065f824e8a33c92156bfe43bc2bbf0e6550432f4b1a5c33b516b5f43f6b71315e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d271bd124a756b913e2f2f2d030f052c912b7ffa6a94a5bac7a31614224165f2065641bc9c42634566b0c09e1a8bb69fcaff31bc1f3b4511bd536d1a65bcc632f790;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127291aaeca7a473ca374464327ca6f9326de583e45e847b75aa2fed8c2f9d76c4e0c367e75effaa5424875ca38ec5e4ee39b5b65bfd3383e018aa79ab19f82b6e0a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ecb77e25b4e4ec870eebaffb5bdecead61ab4ddc97cf0df1f59c45ad1f0296c523ad01df52f599d05ef859b269c1ad83aef8a8cd0ba8e11fdbf327d1eae2be1715a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13786ff25219ff23c48e5d2c870104913d24016e57d37ba8de017c22e937b183fd64a6991c24d8cd15f07f5f5f58ae3e1ec069f189e3c76f9f8941be6de6187db8d53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138046328f00ca6d0110a77fdcc918899441468ac9a65fea630da4d963d72eb449c68ec43bf4fe14ca7215ec9d86c3fcd9feecd3a7d363c0962c583e007f489a64bcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112491d7b54210fbc0fa20281d9c40e939d38559beb62f30b0845944a2a239108ad4a20bb86e0c1585959d73192b121eb56793fb6954cc98c00e2d8f8becd65ef96a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101187b5dab590aa00cc4112b3dc907a05fa56687e8ff5ab24ab64498866367b752bc26a09902b33f5d8a47da0c964b9cb2488733b81da4b9e9811244d96b140ac297;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9e4a00e222da1a5549787284c946a0f69d633f5f5e768b9068c9547c28221726b92e843a4732c62dcb24bb8e5a6067fbd54482b63846f43bdca5a9bca1d816ea834;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187d443c1b4e8ec93a1f9a7b74c4eaf51992954d9fb6210c48eaa536564e72609004b32bebe24d019d943e6bc6db3f57d95c78cdd99b69fdf3536b0af3f28bb79c4a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d21ee6018a4f0822c6ba9689607a18fef455215583568a12af849236bb763d0ead692d336ae83ee56861b87eafbe33e1c1f593d51fe97f797a4871cfd55adb4c5c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0e350ece0ca596125d4eed678a83a4298126a4212acc69efc7ec584f987e280941d314adf4450ca248e92bbce040bf9e31f2c90c3b77f036df794c52a02be514f77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d26312c028176ad56054f6d37e3a7aff6a23899cc7ce469dadf573d7572894e479071deea7f3bf3ff346a61877ac5cb3d7f2110522a811a80a3f942b66b5d1383ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69aef726b80f4f65549bf1b200ef89f2388993e8d1a73ae0aa749e377b37a1a56e29c576a629c0f1af81441f1ffb0485978949dd8f60872ef6b5aef7c3a42861890f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6f740ac6536000079a5b1234a7d80b01ee784cf8aed61cf08cbc3795c7b6b1f19c60aa0603daa348c85bb081e532903bd2b13773da284d63c123850d9d87e2944b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e293847f53b464151cec165c42a13b3c1d88a8781b66ea4f3fb52cf6cfe9b9585e8dd60842d11d742806b3afe6283ce64256db48fad5e0b10a8c1d0e4b4920354f01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffa152ae5b8fa52df1003dbd7fde256b1b8156663ee9d1a93330a2b24725197d357b6fc39b87db395e468fe2537e08f16ef2ea83ece17a43ff93e1afc97a3d3d77e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a31e0afca8c23a93f41a9d96bf783876f924ed8f13a5afbb90ace4b1767af0576e8693ebb7a6eeead1ca22df6f08c889b8aba009b648dbb7b78e42afda834fa16abe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c41aa3150f48cf352d802da0a8b5d125e08fda9c85e4f3ff028de61de92ea9f71df348913cb163f103eb9eb7f3768f82858ab827c3fabd6b52202f36f4d0eddced;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4377c5b28d5693597323253f07da92e3481e4f9f40b8ce1e39a131dc01c451dad0559588b214af3375ec7d5b48fbb8f1c6818f0b99d57f60e39933bd67ba07514b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e723be80295a39bb46500c2ad842227c335341618a553c557c3459ddd4d41ce93838a66cee02a7d38aa0645d7578c353cc9cdf94bb5c55114f4fc7f47c74dedcc11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee381dd4ee899cfc636644293dc832f2de5c9e8349776b7dcfd72138e6d4d80383f0c15812f963864899a5e76642e307bc5f29a15374ad0f487e436673cd986bac2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137b6554ea60b9b386a315ef1e7b741f57626d1fadeb5e01839fd28112835fcd8b26f8695b6ce64ce70ee19ec33685839acf193866d4df3b853196d29604a1665eb1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac5ffb2ff2889ad854a7fe80c46c04a28e660cefd393d24f016321951565aeb751cec0a7f71348325bddf9f08562e9b223900847a3536904d8c4dd68ad7eff15945;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9786353f1bbd173e8965fd3d546178945bca1f07a7ac105535b92918d3f44997bf7c3d56b5366ab587c883de5de980c4f0ed15f719dba66e5c3ad7155a481d3c0bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e681f05b020769c659a9c99f690dcb3028752a295f6aad39ccf60a8df7c14dbb1bff14be679eb62ba1cd33ab7b4ebd6764f81299ffef1624ae400f2e9192839d402;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb734a8571f3fcc32c0630fac7b8500b7b0ce7e45b603a0a6d3148311bee0aabf122cdbd02f3afae978b44a5957b3a9d735b8cd75eb73d8c0eff57bc41f721244ff71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10435ed4878d0fcda998fffbbb6500e83265e7c304347e1e09fe95d7ecb6b6238dc10e86cc6fedb4f43d8066dfd0a65e264b2c3e6c0498952f6eff4e7f09e0a946bbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156ce5263e7df2bc6cf63a45d59327d65c20b8e0061c7db2e9ea78d58e47e00dd40b247dc4792e78fcba65062342bc6ec9506a3254dc3b1689b8cab605e878b42dfe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2cc3d6a2f73f56aeb3cb3d1291530281a87ac50695db2ef9036f026cfca3f9ea263b1c20bf54ecfdb19a19edceebdc2bd95fad6b9ffa71d101e69043c16b7f56265;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2f7fe5ca011ac973ff6bcb742b484e965e92e786804eebdff4c16b37783e05b3f1b6e542e386fae64c69476c82d05c148485769fb13bbb6434ae7281cb5e5b0966e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5b545eb9d79986dcdcd17277243893e8c7e6bdfc0a7634e71c8580e2f86df799d3e489f152ff335d414e8870a4abf3aa5c71d865976d219451470089fafe78fe97b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab522567d3d10d6725a932bca696791231863d3180e0fe497bf94dfcb37ba7cc63dcb5243c7d186e21f37b606bc61b3d882bd51bdd0451c0b548021b4d9434935990;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ebfd6b31cbd75de0161e1570797040d89ffebcd8bad744c6ae9f3bdc5401e3bdb0924333c3f0e32d06b128564058c4112f17dc96e71f1eb0d1da9ebeb71f1e79f31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24f3883e3615baef84b24d2f6e9c5d23a28a2e5aac35eab20edc0e64b9be2acf57e2673786a548bb2d43dcdb2eb9524927de5bb216998d9223fad9664f6cce33d017;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c90dc29bfc747f67528a13072551e3856aac610134b9a07cee2ba5bebd0341701e53e2034e7580cce402f6629d6616262ef941ccb476feebbe30e7681319793e01f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b733bdc0be1777664610f5688db0bfe531ed20107282478a76b1ae96babb9ece068a0b165455f84a44e72167834f698e453f452466722d0da8816f1907f48c236214;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fdbf50957049ae49cadce1dbda98bcf1e43c601a614e22b11a80366478085201bd73c52e1d290bd1fb4a2d96ee4b6c145b6461ef019899cef678d92ae840fcea77c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66a79630f44cf1d4c57a7748e630a86126f3d5a6f3c5576fced4c176d4e771d53ae1c93e35cd0c7becafd77749c46d5af3aeb4b00de7afa235e1df64c7662bd9a2ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e5f537795cf7065a78d3f61c13485233023fca2cf9aa85771f3a01ef7de4e9aa3a7e549c366dccd0735e041e21a73c2a8a3d54ee5599c5c6d65b33c1dcb63fc76f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb5e88487e106869f306290f9212619dbe6f27e95c65ddf84bb9d46101ed97ba92baf77dd62c7562189c242cb4f44d0ab64dd6b694b7070b589fb4701094ac3642fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74610ca8acfb84af31ac430b30d8b9a239cc4fb2fce0396d7d9087762565a2fd3a39cc2eb87af1f85d1235746c845cf4728075121a29599ab5654cebf90fbcc7abf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f982cc73f9093141676684061e4ebefd1285e9a4b1b23b3e41b67506534c3975f994378e2d89f80bfbbf71383b4835e68f05864d40175e2870ac886e1df698adc6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0a9c49107b33395168a80c69336dc00da7aea8d3569e3fd70d686be3dc0ee23e1aa16375c1f76374831e3efadedc4355f8c56cfc191465961c5b85bd2843b4b5960;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5ba790c68a4019a9cee3cce87b1b5aac0912936a8ae9b4d10576fcba2520570c7f0b2b76c945957077501f225b5e71e5dad7af700302c85cfaa54fb1a3045376be9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h547bdfec0cd54c5e87596a2a0b56993601672dcf4c253ae9448077746c9c46b05e371803c4715f3992e99cb5c1c927e09d39de42102cf55bd380b4f821f5e5f2fdf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c3e697a49485516ea96b5091749a11d9a6c09734ff67729271e59610fcf38ec1fce0a9c0af4a1ccbebc9d28ccf32a4a870e3005d5b8d3555ffd1659bddd5fc5bdd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h419afe0cd2e75bf8eedba925409b5d591b4f180637dee41b99089699989c58195c087fa16887f260113bf26b8d129ed40a9da37bf2018726767f9fb6bf05434329fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h869f92d1ccab6ac5117587ced1d118514dca6c1af58773d0eac8dfb4c3767889699e0a369efb9e123e7eda859c86ac23b5cb8261aa9e63c9122543b0d1d6a68ea679;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1613ce92513724b77bea12b057461a6c0ea3126f4a97faca8fb54cc82cfb3a5e01500c4f628a6bee5e02d2b025115d065dd88e85e0959e592bda196d74f0422b71efb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h800dd98d236d6dacf6ef6242d25fe1e7ca4a4a0be769d1f59c97eecd4590d7ae98ca40c56218f5fad59cc17cb0655cb65e3da420d768fbdb7048cf645b09281dbce3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132997887ae86121696cd184a392597c115be903d02289f541da214560e9af406b0b9b4031d8c3fe3f560dfcd146c3105d0c9dad32fb51448cd3d49345827a0d01844;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h754e88ecc5de7b043edce5cff8f5eb889b6dbb5b977c726b514848ce166b7fa1cd2255ee0146fca9f8a5923bf8c755e34c5582a581f4f525c3273ffea9fbc693b87b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18001feb51cc80a66d3daec9f31f03516367bafef995e78f6a48e3bd6a714a0d36111867199ed4483020b14b8a51d59b1530bd792ae4f75c3e133fb3ad4e742abb948;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h753c61b92427cb09c098a5fa274c4684368cf3955c707e7f05d6bb59e14869ee3b107a9b632a5ecc9d756d8b000d2df95cddb19ca509e26eb732bb65d3a5487e87c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7e5e2bc9d2f267d65e9426886d208f92574ca106ab7038f766b8e2f04ac5c99608443527c2a3635af0dd477cd4052b01b6946520f8d0b276101094c97707ef9914b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca6029ab5d9750d238ebe0c95a5fc14b5ea70ce7e16d115be656f3e3b3a6bfedc30b55becf06883f42bd4b609c1ea27ab42780cdac52800d0f29c66aa152d9d48e0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h624e3a5534335e232da72e7867cc8aaeefde37a8130964c6fe31d0e7c35a020dbeb3b7eeb4a51c4b05d10835c4ef7b591a9349a63e71a80478c55a2117a2a5aefea8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1107cb8500108ee7064716ddba06de3c6d29294da455711192e386b1a82a1edde187dc37a6a0aa8f1f831a4e58b269cbd418de0876025c0a916da017fbec588691a14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9645c79dad3f65b9f87dbd05039c56756bbb15927bc57c153e445f7786c3c37e8f8a820ae343a9f7e04de1c67afe526bf422de198bbf0437874b5cc534bd0214144;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cab61774883880c0a21f7ddf688ad4cb0f972875fbb84953e8963b5be5b188b40267b07c3ef3d044f0eb5a791704914da7e726a68a7aa04aa1a1ba7619a95bad8bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdb0a731449b1987165ecf1e97ba74748e91cba8b1db76237c8bc0d318ce0adad99cafbe7b0e05426b852dc6454b132f2b5f99b3694ed70879253837e022a1f4309;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14055fb22a27adcf861746ecde953c9ed337a1589f44a30572ddb446610cb2f6456aceb192990ab179646de17e9ee668de438f3d536b9f50eb129f81fb1b94f9b2256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb88dfa4e0d193cfad7381ee621401afd23c96103ba8dc1105ed782da7be69b3edb329a55760cf75104e9f8f0e5926ea808192c26945e7188772da953661e3e36b767;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ee2393626a217afbb8f693213baff2454dcb87312a8f46ebea6c28ce12d9d624b46c3a544c131a837a211058df25fbcb9fc3b3c00859dcc924680a39a2987e8e6b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1767cc449ac7bb928a617ea08bf6a0ced0c2e654836703009b2dc36071c798905ec9facf5c8906368d984f5119f863d4b3938d5e9291410516bc5c54f2c7e42f3176a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he604fc3d57fdf8e741b40fdf4647bc5387a7495c7f3fbf72a6bdf8693fb6cd2a074144820f54db8fa56a9cd2cb82f2562775f6a44deb921de2b08d845420d9b94325;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a313dc0e4b0fe752ac1a47c33807514a2495eb702424cbd0b7a8676a9df9f79c1e8c030c63bae02cfddcbcfabfaac21d95eba7cc45d6f848dfb11263f33d8f676cc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3159cb5fc898adbc11cd1e3d45b89a39ec18ceb9a79b608b81d19ee4e37c14781bb5a5120b80b35d88932b41e3b85a07a45fd93869ee5ec1f13b11825b6a180461;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1403ac6bd90d32917e366dbfcebd0b1d0dbccd657e82a6ec130ef9d41e8362f5efbe3cb92a6ee7358b5fe2a0cdb63baf3091fec1156cccaf9e3a73ee30fe0a3f8052d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19dd0bb3275cb79c6600f591f06b67ce98aef4292b82cd328bda3b18a6dd44a40e32b87c879dba7da229e77e9a8403eaf03c0d038897ef4a5f04d8cb34ec76ceeed32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dfd70441233a8b7914ef6f8d17ca2236f58aada5d9450dd9c62cfc68e04823fd3ad4b6f56445f7c6957191ac89be27ce55b1eeda494bb55bfd5c7669403d03f04c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e6b6289995e332dc5477b43c11a2efdc57b3ff4fdb4b53663b84c114c7d9d278ed5118deae1a99506793febe2a546b3d22b53027b8e356d2556d939d17b6fcc690a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h323586889e3577d7ac4906789260eed3e505c45caf0c4782783e43116cf37e66ad907ce033f9b7372847d043776053683dce751a7e39cc8ac57332ec7390568ee074;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3b798a2ac285e238a1206dd0896ee4529d325524d35635507ed2530f2ab8138e42407c492b10f58126c27920578496a71685e42a52579d670bbab24370743de6803;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc968b22d3dcb7acffd45397a8f59860cf5820eac977c31dfe4f0747fe234cf6ab0f56a982f989e7184c3ce53d2ee38cbda53bc68c4f77933602a47c139e0bf56191b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2f608fa8f444995c968dc41a94659fdc7335580843d35729a3b44bb0c86386a930bc2aa2396f9d985457dc87e963f308b32dfcaa3e4b5963d6ea730b59cb487254c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2a86658841c49e21eb77f99444db25c949ce5b65f50fc0e0c31c2ff997b0125c651e95956a70f3d874ce7e78d86bda69e0bef3d8bc19554f9f6586856b19016d0ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e8d43060663ed1b2fb6c9b7ed8e23dc533947dd3aff23b7fc98e3fa78e292ed44c1b9697b2e002e354cde6c07a164e77577374c98fcf72947cdfb5dc7c1b26773aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1439e76f529570ed6a6e2ffae57a7f5b722d703dfbce78b11bc3f2135dc94af1b28df34a2856c07dd3f51355ceb813ec7745a31e228b66d1dc94da5b6ff285eeb69fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h713855ec6b628e03071b070d8c1361d7522f035ed906d6f19c598897d09e0705784ed7df29b7d9fc939bbce9ca7a42e96feb2d94499a9722a1552e84c55dce18260a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f146ee60354fa0c7dc91f7599c2c8387ca77e59ed61bdde802ece996829414edd1c484fdce962693fc1eb1735df20a670599120969ec68237cb694f1db8874f9a1ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2e1928395dcf4dcda0ca2df981e242cdf7b7188d6c09b519d81258a8d28f52e4668edb96de13c64f90b83e5670e475e05c3f171730a70eb7fcf4a0ba8bab3c686fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1246bfde7a728aafb2553335432b77909e9fd0ee9f244dcc1626aa3263ea733ab771fefc0c878781ef1a9f1cb26fb144a2fa8a5e07e1f87fe2cded740d7c8e98304de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16843e8f3165017cd73cfdd9c85ff91b1cffe98a285ac5e1ae25222519e129f06f86cf9bf9a7fa2330a443b0f6919935ca6a3676829a6df2867b3a1be0362daf1240f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183850265ae4f069ff7647d80635fc0946e5bb92f3f014eb957f747e96cc05909f578f542908802c4ba314029f03e94f5ac8159daaee6035afb0961d84054eeac35a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150ad538cc24873ed4c2af5bf85fbd94247f03d71e45e712a8998f27326bd9031bfe9e9c7e0459c96afe69fcabb9f6958bf1fce509aaec7ef2f6af3807f65ee33e7f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14419bfb741958a4379ea31456c4fe13f8621ecdc920797d7655ac4d5a31c023302bd220c4c4891f3bd4bd7b17b0d1ef1a3a50d1060ac74912c9706eaf2fbb8cdcfec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddb44cbf16bb8d487dfee6d3e1b566332d26a7f705273467cb77303a512c789081611eb25cdb56acad73a318dbece8d3fa1462b8d5ca9baaeca4098432d0acccb58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4340f35df32edfff326357a0dc41d381da7bbb49ca705263a6a455fb45b19b5a12c7cc310b8b776aa5befd1e15952acc1d7ab062c769b9bea8f2dd8c0473330aec0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103c3cc767b052842d13e7b7aaa61abe6313703f7e260868d973e977ecd03518ac860cff239b27640902a0979b1d8e03d4fdac85e574a58fc0096a9507f3ea5b42383;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h842c1246642305b1b346e87304a7d24e897f313da6bc119ead5df0c38f3710069656c0cfa91dd06384881d83afeea42db5ae16781589a89ca99944440bf1062a74d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d3a34a6652e8fe16bc7fdfb8dacaf4a9d5128e72ae89c1cc1ff5d1d6d8cf23afe8bde2b1b834f3e3ba7739a2bea6a80738a63b1c913acebb142a7afba8c8c521f86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1069610ec139d066100d6c601eca7cfbd46cde6ae5197cddbd325f04fae7660e25c496c13be0bd7931d18e5735c1e7b5e8f63904f9373ace78c0cfa5a6ac8a3b95846;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28d759f41395694920ad77f5cff484c86350755c02fdbd680dbe5e88693db2a51bc9d42be0537f81528355a9c6d060e205060933806872701c0bb81d1c6dc591b3dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faae84a33f5d2e561136773ca0bbe2bb66287f5b8af4564b6756efca5c2845a8826927b16abb340f6d6484d6997a40a4d2b0b7f1e058d1d3f939a16e35ddfc616a62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d86ec9d2521c6b4ab45775d84126cd912ce2c6bbd5bc38d9495b8bbb353c2cdeb6751fd49f29fee649edb9a11e0fc2acd60f62b6427dfd04b80d85533ac712ec8ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee9d6384ebb1f41d5f9a67f4ae81dc269cdd6779b9beb56e592c2b3e340c224968dfd08035d01638202139aaa9c916c444a118f21ad3e938636259d8fbaf8e5b75ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff5bdba94c38702ba3e64d751b32d33d6b4877b45fc941cf609b590cd9a78df58705073554a91677d247d7e27edd534fe8af3a73a3c9e27c72db9c6260910af2fd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haef5de82e75db4fe4de32e7682d09ec0354daa47a29b9fbcfdb985f32bd763235a8e7a8d62832f5179a768f72d6ff5ed9b83f2b1dc1e63a4cd9e42e9adffa335749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a35c3059634f3bbea5558efaa8fddc657e12a1b6c9005cf282eb430b6d5494b1983bc6ed0d3e5e7862f4cbd39c5df82577366202b74815e16f1ee323f3f1017027e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd339feef9a7513ceacdac7a4e3517b83a9636cf068b8265333cccb21d387d2a5d092a70a93fb743c341405fd09e3eb614f6dcb8a2de6dfb8b5a6683a3a6416b898bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6518a035c711a5b109465e907ec8d90abdd4b45c54c530080107ea32d767ceda7531b2a57c928930db42ac0faecb2ae390f96c43f2b3daee8e898e73a3d013e8a5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bbdcdc5f3ce5866015ac1daf2ed86200a13998da10159527d52555e9ba7f0fa6ddc8b5fd18a4944811b4339c32696d4727935b33053584fcc9eb03556c33376a7bb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5384025e210fc6fc204ab481f21ac8456645383d06d8b0842b64fcd6434759a9178d410ed8911ded9dacc7bdf47e34068b86134a5916722631f6b914bae9eae903f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he11a43ad97b907dae489664b0399f1f195180d334d3442504299ba84913523f38b67dffbdc29a24fded1da73c0464cd0f3332a877b3a53835cb17529f81679683452;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150d30afb735dbc1ae94bcaa200b87ad1473f324c01b33653a9b98b779c02568ab5521826d7bbfbfdcc49af17cd552b7ba13f47cd54624a2383ff927dcd9b138493c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54743066ed1a8b231ffae3271094bca1ccedcb51ff7ca019105b3bb3228f5321e34b5a262ff42e1f735bfa59acc31839fa4d872fdffd2138840fe7d40efa1ab8bb91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12707de05db9df63a162c290023fe73e98e603f3833a284406a28757bc78f3bcd13e70235f1b4eb6db272501e32596439212dcc406eb4ee53662700aef2b45be1b305;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48c95fcb21bcad741b6402f164762b0471645b79aa54c82e5c3042d1351d20a596df80a990213fb181df62ce69a0cd122d2df95bc2a551c88c2e2f7db200c90a0ca9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186ae6fe793d3279d84e70e943606291a2095ceca956e2c4a8009e48763aa8ec6ffe5f52a36d217ff83e7d444810cb44525e59e960f80ca32b702e729d55035d8d14b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133f22c98c9ef9783958d0ae7ed996970c5fc77f0b35e5e368567ccd871da48141ea225ac67c2153d3862bc2857ce44cda29ef0eac60dfc7eb01706b54990c3da414b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11cbed7f178f4d94049f3208c7ba2cb81f9aebef9499eeb2b28b893e1c5fa3885201131cbc5ac2f6673e434e415fce92d0546ef8492f4608f8bb60793f6862ab03810;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19313a77733a7222020a57a7fb21e514d3e4ecadb921e4c4553cbf1c605805ab32bbb5e3295c662a1985691ea7bcca257d93ceb3de02c2fd1faf5ce9b628c25ed2fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d5df306d5561d157ed418c836ccb4d3488653a2d8cc4ab5995cb654fcad0a8c7d18d65c6055c5091c618210738fcb4a81ce6929b7852c562e6be15e3d081896c71c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1827198d99dd7ecb071528f2f2448d69aab822fa5560866fae40e0568a840b710b9a561dc2158a0557aa8b1bf54a20773c9bc37a34b42b7837d14030c21255b3e331d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fd9f39634feacce5b18dee3c333e820f686da157eaabe7dd060bb1b2b57f7e6d94ff922c1dc4e6ed99b5e2e22c427ca63a9e1058bba88c2eccdadba6de5ec804c26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101235ebc3ff2b91e2793b8684b776e59ea77992041d06a1842dd87bc20f4c98169b341457079de1f6c6c218c8e3df26b9288d95424ed04ea264139eed6bae046a7a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17025fc500d492cf7e8d3421e5bf38e5d9e760356829eb1edfe678c0ed808a0fc3e729af9678473b9ef8b9fca69d7afdaac9cd722912003abc82024d45d790c02d25c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4700c8e828ce3fc7b94b7602d40d61e142018cefd9d5d1f0c6f3c6562c4864a21e41b9baeba9fd237954ab1b02149a4b9b6b5d6f09c40e7ebc78990f47ea631fb38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150066d0d8703b816ab85eac8471504bbac103483fad0cb0079ac6663dfb6ec8e0bcaa0e3a1ffb6923c86f21890656a94f1d478620e5b662f927f481dda64989e71ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121fc7d968cdec015c5158e981d1b370d96ff02269fa3199e7cf5576794260bf4e5d0ebf832f12d070fad8f96353f57296b93a5b287dfaa954c5807c472221b126b84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1e03f559b504d0a49d2a829a15523799ba67af4731e620926945de75a2f4844013629fe505b236036bb888f51bf884f31d55c1968f094ee234b1b93e7e6c0bb93d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152b238126845c3f2ef0f5ee6aee3d8d71107ddbb1b7dc75a20eb4bc0d23c820b455487247182d9be79f6f1280f8b940acc49c0fb6a848370f0bb1d3c5357a8537bf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a7e6b510241b8fff51df93afdf2e3878a2b6e36abc34325f6f65d5b9548da0c442bbb87a1deb096533d1a5c7cad3e91899662d6fc570ab99354a273297026164001;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17072bf796ac83e8a4f31505dc43279c9aa72e56cce48e7bc127a82aa538e005d169300dd88cf4286b1662887a4b7bc4224b924876d3b1a5a99526077ed84b768b73c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0f44a23908d54cdd89a8ca9dbbe556b94b1a6199b23c8292f40028dad9d1b4158945104629268a9e11a9631ccef043cede48975397c70c417c17b93e8ceaecc86da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa701f4ce56f83c7a9ab3a88e17fa6ff23cdcd320ccdbc68e25966a18850eeda0db87e5441490dff01d2aae0ee1543451e45a0d0506ad102e2a9ab4cd13d2a7309eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e44f19dd2087a56022bd390d7c4738914c788362e33ff2abec78c5ba01a5f90f06a1e903e5d396841d7f38d60fd400058d454fcb169587602f3c2cf3ad6a608828b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69b795a3d133c0d47baf139fb53eb66240224809717f9c4e042b62c4803e543527a3e28e186ff4657c233485b9c1222fda19027e0a2e657d7bb589e3f1c0dcf10086;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10dee53767aca3f8fa0684818b47410a410aa2c707aca9550106aa91b51d52ecc235a8d09bfa3d116f621b7529a2e293053c6eb4e936e7637b2ff9e286cdffc68b007;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4da9f70031b717dfa9f27bfe30f67e5ec21f1eb8acd5b19634e8bf1fa953a6c35278df2c3ed714fd3f53c059d4e3b74f15344297c86c5490a668d1e94342b597daf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h283467166de58beece9acdf0454eb5e4547608967731d7aa58dc36b1fd4c4ca8e702ed22342d6502acbf6c6123562ebe206ff271ec39221e4e93cad9a528a56dc002;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24e58f156699a8149936e6a21d4a5cda361ea2f196124606dd8ff8350e1ae6d064611acfd685eceae95849dcdf98611275d6dac88039b0565bcaa412d138974874f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25387110bf1fedd6bded6003e4b8a0aa9b42c3496fe2eeb38159c8d9636749579751cd871f2278fbb63c00ddb1d1f52d7dc86eee546958bea62937e91d42e8b760ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h948d528cbfdfb91b93be21433f37460cba9436a2c954d52a12365823d69a35857d851c6f9d11f2b42a0bcfd84b930b7bceda3abff8005eb211886636a8426c2d00a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e5920f22f15399ffec96b781b163cbb4176ce7b994e466238be74f01e9afccb04ad556fe2af0a176c2c5086e834c302047b5650b4c8852d89d77be92ca725a47bda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190d3f16365596c15208d9944f12922f293a1a54ea21ca3ff6b8078a945958ebeb284a000f81b37e469235cadf8e70cc68d13ce8793388c0b6610dd761704e9d02eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h251c886edeeda6aecfbbaeece3b9215032f40a9dc950f1468da820e8baa3d9a62994cf209113d10f0a0547f6359191ee399c7a440669d3f33d31af451e65aa1394a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4a2cfd1a74e4e997f54136e411f4407f26759f65f1e902ca5c25f4c8e6c4396ecdd8b10ca8276158f02d492e8792f39dc9a966683db18fb5d2a504fc3434004e68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb3ae50f9071423457f266e3ff8a4dca0b71acc2e3e4ca9f4e7ff24773712d3accc67b49f1b7bba26977031999fb8eb8908c33c9cd56633a59b3a4dc37bc8d30150e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1079bdd6d1737ed5c10cd1c1fbb5487a94a8c907d5e6bb33d1ae0c197f944a4c0001a3e08f4f130c5957e4e46709771c4f0e829f27fcff170a0b7b2c6bbcb7d3cb2c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca989583bf973b1d289310bb14fab3c4240d93e0e3e52335befca89beaafef4d408836bb7e8bd938aa426551a05443108badc770e7657d6b060e13251fd4f49cb7ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae2d93838ee358d7aed86e4b5fd17a04e81053cc7c77ea25224fbc83f37f210e9269b5f63f06146ad40f964460b6d594978fc25bb0aa6a67b113895c413a5ef1bc4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153de337a9c26eeab51afe235ee7e06035d94b99e526fe71e73572245103171dc844f042fe775b48be3654f720cb7cfcaaaaa7cb16a39ae6609d2bb11d88c76781979;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e37017ae01d4489b0904ecb6f1893ddb3b8846e356a66614ccdb8d78f2c8592a91915c86038f8f1bb56ed74bdf0a6f7db9b5d996a93d91963351bbb20d7c1f155e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162a72c21b46d6039794349c3367a24fb3212edc68e3f49cd86a98a8295e1a37aeb454a7486c82a0aa473676fbf05d876dbf1e8c825a0f86d0397d9f077ef0407be0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127f0d41906e8d8ed7408d7435cea85bedf2e9c2af08de6b616126fe75f5fa9f6b39dec89f971e7aa1e72172060a2ef101eaf977a230c282ed67e6255831a2889ecbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa51bad6d8f9db179e70f2b79f0cf96e21db36edf7dce9dbada5b7959eef60ca546bce54435ec349b5660365411ce1fb209553d4b29fef436b7d5b882a942baa5b93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1a5709b9342c9ba760311139b10c5b2cd2c0ee519f41f6393fc30b1544caceab61d54ad9edf9363fe6d6e3baa15e81ee209ebbb8664a7a3eac66e497def8e7b8121;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1888255a2414d196e1552140b1001930b3aa7144cc15cb73ac5e1fd94afa1469ef591c9ecac980983eac7164d053f080d866a7f0d42a725a89b99117a39587a16afd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d8d10b750c8affcaa59654da15dc298ae0bbbeec6171213a88e04ad66a64658f04b44e11278a9e0c253081895640f424c00cc32054d02bcc9a0f8038a4b78545bd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3215e4b9533989a57dd2ce6b864a611d6f1d99dc6726e6da6254807a9a69878b36ddbdd346f41ecb68abb2a2fffeb8083caceb477c943471d7db611247298aac2691;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h439df94554c5c989ae0050356f4200912484bf718c1479c4d189a7398f488dd1d3a9381ac36e9ddfccbb0741f35b0c377c6176b59134822277166917c14348e0a5b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146146c064f2acea3b1fa25fd3db2fbd083024f7885b897d247bc0d532fee365126a1502becbfd8825ba4b85cf7e9dc579eb1f3cc8bdec9f87e2a7b4dfb93af984f8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116261209e0a5d8f029fcc93fa99f396a8d9e1f5e1af4e21208506ae5ebc5edcf07167d637b6f41f37b3cb031c64562b665758a8c66415d7d2676b442c20df4d708d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d0d66079136b4185f2915500bdf724e6e5c7b7ea49e194e676239c0141354aab0026902ef4680d8eb358105032cef8a798f336c3320cb58cf604fe3031b0ba5fd3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199c89473d6f09d355f88448e4dad41652e1267fd5b808862dc5ac80eb9e2c6e5a55da35e40d613c0b1d5b1729be67f4267090e4215ef4f9fbbbf0df136212bee14f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c360f291286ba5c7c232146555ef6ff0caf9d9f12368d0ced9fd2ce661e928c63337390609e3f5760f978f0caf82f11b603fde13512cd331af8112850b0932bde66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf300ebf9cef9b8c2613f190baa20a9d2bcdc8d9118e8f1c239e6c5cc521d1c53c113fd4dcc401d5eca689f64a70a68a8abf993685762d3ac875579786d56727b13be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c69f1e34ef5c4fb83f12bd7989b5b9a991f9c8cacb051a4cf07eb47bfe95db1e8200e6b54bdd7615e70bf6f83751f0e05273a5ee3c0206bd4cf25b7acea1617a6372;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he491c008c79cc70edf362a0aa51cd400786c34b6071fed5045df09045c3136cfc26301b0e2762ce6f02560f008c7e290beed37fed7bb734c4c8dcd181ba465649cfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1975ed9f9fbee8a99bdc36c51e7d054c8ca21e950ccaddd19098391492908c5558dc3770ab7dd06a9de21b5545c6f1c013218e6c2b478625a9962cdf966e3da4fea0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2cb208b0aeda86085b36ae1ce5b8a6002bf88cfcfa488302ff93357c6efa6b0112cf60ebf813bb38e313c9ce8719af7e404130fd0c49b79af0c6a078c347e7497f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h919a81b843d3381aef7890949736b1ec5f76eae7add7c1950c85e63759be34104ca33bfce0bc7ef51b5ac89bd8e11268db6df9f34d13c9041b3e2aca4dbfad85214;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefcd586e97c94fbf66fe015e3f89074bef1704fbd36007dcfd8f537ea4477d77a6039b682159ad1916e279d1266f0b4e2ed57fead3f30ef8264e12468db65a721b9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h584ce3c199f55dc5a27d3ef4aac113485f8ca7fd3a37ef71c821a8755e0c6c9fe69971f392ef184d88af23643833cfa11f05ab42e8ddc4468cd6e29f264abe23e043;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd92b3bf2b7c1cb15bcfc32496771b2b40dde741d4c39348e51686f330533e53265b856a5fe53660767b920418cb1bda7da79cd8e3ea1ff54a263d6d9953bd67b650;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cbbe730306789e222a33bdb020835a64c648c4fa765896f33647367beb57f466b30c8686bbdfecf191f12c2ae079ca0a8d9cd838163b858a57e9689067d2d0b994e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1897031c740ea3ca6c9808433a649fadd81c6875060e8984942b413c806ee2356e8c3fe45962c7c6a21006198c0cb1a8796e6d5dd063914eb8665fa74b63f5cddc914;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188c3a83240d5c10f958a319be2742632fd8b50f499f957e8fb5c39b071d0e4ada6c86d31067efe2ec4de598de43ec9188f462cfb37fc0714e78622d3fedaf19ed749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d7461798e8ced8278819b5df5bf52aba3333844d6199fe185c81147ba6aac74d23712147f06c0d43f84549283646647dc3bcc5e37dafe2ab7e22a1ba13e2ef1d4d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a09a1b4f65a9049eacd395c6444dcba9339814a776eabf32791f2ebe48e0acb93638640bfb8a820ab0cfbc509d1dfadb0041fed492e92f48c49c5a4a7ba4a4b894d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129744429fb646a85e0d05247acbcc8670e508d47ac357598e9e8fbd18e78d0e74b42c19127eeb30cc98fc2957572159eda43ad7a2146e0d2186326befa5bcf8406fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c6f870fdf43440d08c8a37f372f36e3c875d0ef5ce74860947cd16ed35a012975079123c9dea4efa1411f31541cfc1ebbfa8e6fa37568368bda288d30492c0a327a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd931e1c6fc4fb632abda865b9c0127005f61bfaf4ca3ba23fd47c783e562332d29f5b64bc2b3d9c21c3ddf08a044d77d5e18527741c998a7dbb5d63a815906f6794;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1406ab587358b084b939c593dea41d086197c90ce8c1e961889f27407556ef7cef8ba9b2c7b21a303cdd6b4e8b51b8594c9fa35c5227faac586bcb0e72d221d67f190;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eed15071560873123b5f6dbe78e9803b67c98cef4af8a37e7820bfcd9e5f4fc9b0e40f78b69a73f48dd4382830e5f1c959a5c7ba6a89e3ed4e5fe757635efcda1fb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1371c2789496ad3486af5ef88d8bcafd2e790dc39487050a6a1945029b2b68edfe4a53b3541d30700b4b3075e125d896ebb59f19e55aed7640e6f307166d83cb08eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h624064a22954d7144b5b55f2e5643ca01bb026146e8e8bcdcff428c081081c8723e02fff019dc63ea5ceab319cbfe7a4ee217d34041494cdf280c7b11b36fa288cbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4fc8acb246638bf0f8de58702c8ac27b3a59ded5f31f146f1b83203bf6eb936c92df3b593a48984ef88e965e1eb0b7f2fcee8d193cdfd5be8e55f8d69f6213a0efc0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d769e98ff5d4490b109ea700d910ad6f52459db1a3447403cf21451ea44f3fde8681fa26718231ed6175415d7c5463ff770b0f823abf63b9f007f3b4e0f582461790;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190dafcb65a65d244bb8b97bb8a52628ef7f6b862ac9b35f86710dbd927c43059a26a957ba9c957953dfed19544c5a36c94d0b36a9e493200efbc09f13023e8fd9ad1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c89163e5b779ef250a3ed7d6e693dea91c68c16dfc7e3af8edcc2d1c991ba03f102e5a33025773a80ce785429d6fb0a2c34a100a19b71cbdddf8e8a9cd783ea50244;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf8e857aa677ab58078cd4195369f0249a644af54b3f6006ade5db0b807f216fe8e827806261d96c35bd1c6faf4c202a483acdc2eb2700a307e200057a73e001303c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11299d59e18f57953733db6506ae2e21668babc8fd9cd2158dfb130fc72c1a60ce16fbb19c85f3c543705fab56a7882d29707ebcee1cbd97d2271601dd2eac5cd9562;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60be581ec448b35487bf0cd183c5d9b9516bc4cd188c293dd454eebc0cc54fbd8bea4bd4a5f12ed700d994645988805eea2587fb3c762e52b9b02f07b42ebd69edbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdefbb3b049cb574e1c2970e332e56d7054b2120feb14a6251b7ac097dfbfc25c323f890c2d4423ef4c928bd8a8b5bcffd9a32d8600047cb18578945eb64efa2ee1ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd611a8e8f0c19949f386790e047cb99a31836a368373e966945990355f8c1b02ca7d478c9a7f89a239d750da0ba17308d645208a41566c580b147eee71cb0a94fe1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb51bc107b3b74347c286e38b4393e722dc9b4b16fee6c417049aa9525e227a144eda0d2fef42e4e53f51f24eabb6ada030543a6425a8df3c55f4d42bedcc61d0e5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6846acf73334f62ec3c5d31ba9601c33aedd4487efa36eb4c1b84b32ce2d4e8db221cea33bb9cee45804ca58a17a9263f4632ab58964c4cb01b07df533f32bc4ac99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b3f7ea33abad7cfc8793b31da8ee706f7e7ffade3a095d77720d15bd8f13aaf54594e24b5a01e2700806d3414264eaeb47a02e717daac96cc568746a25b452196f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c5ecb8c9bbb7d3dd263955a6f8ed16982ead6cdaf3bd6de1d5fd7417da8ab194ed1e638cff5d240e6c734b655c518147d17cc8f39553fca9f2640b2ba0c000ae1ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc13942bde20a1581e122a79090a38c3e30fa48fe7c829255ac22e331331a7ccf0aad664f97e45ff8a27058d2228bf6242404680d7c2100c8914dd25c59c2aa4a84b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a04b827c3cde006f03bfebb810026fa28e32c05ee4599c61580f04854ce0cfeab883af3976cb4d106a9c647f47a95d3965c5e0632e485b3bb1b59d413b5e255de26b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cd0bf91cdcc6f194c2c694a6fd8f765bbb11e99500e79fc60f22bbe086b44c3f5980e59dd22ada5c7efb2cb0bdc6c6e4e9bde5ef183b60429111ac48a1fe7a778aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe94340c8bd6f89d23dce395bcce67ee6a41458f1d912f8471b3e2fc67c46fba58a0460b9f8d1850988aba1bd9d0ac7519915a59c00b233daecdb354d5b564c6364a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8ccbc52ce7586d94da5880e0eda70216328fa9af14d3e598887edac4c613d9b0800ce7a07db974633060d6c8d31f1a3b0c83c90d81d8d9015685ee7bb83d74e3160;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c98771de91893cfecb8a5456ea034f3c1b6ab2e1aa215a9ff3aed1ec866a0894792dc07b90b35d6031652d50f9ff35dcc073fe26fbaedeb78eb4f1b333a42f22b41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17cf7fe8ac75e43fe628474c7ee676f85584ee8251798739387a0313d9f8b637c259e876ebb2178213990f5813bafdbe90c57f56e9e16d18f8d290b78705b20d6c4ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ba3a1c507ecf39e688d95c91609f114f348bf67e017a4c00192065ba5e0b1c7b3ed53e285df7c048be8fd3e1b1dba0634d9b3b22728b3c7ed2b03981823d8cb9d95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c81ec931acbf64d8de8b029342229497e97ff98b4c80e8e443b366f9ceb8de95c8db9d540ccb1f714d2af217ffcda292759e3400401ce7e8e4e5848c3dc13c5fa47b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79402d56a21141c36be4879218c223d523ce0698899f95e0ba32b6e9772d635023edaa1c8fcc3f0c0cfb1037f4bfe153010f23ec40957c0cb862303a5320f9473e85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164be81e39fd5fc0541b5b22bcd2702c549bca9c2e11dc730d6a5fc4f18998537f5a86f827485ec2cfe0eed74673d7c247bd1cd5ccc092d100ec912fc1ddc67ed4c64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89d2cbbd87c3ec82eca7de4fb03a5987fabb6bb3f500b3c8d4ace48858ec40acfb67a0bf3c23d3465b24b81e4d500ac6be6b15401812e9305a52fd6db0aa008d6c19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a695a7b005c8fd06ccf78f6a3ce017ae8ac40cd5a069e1f806e378e978afe83b1ab0391f89ee439c28dac72f04bbb52d071d69c84675071e037b028f1acf93bec6c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6ba9d479561ca2e9e6e2df32947f53f785908dc9a85e395285446bc6074ae031e5139b4b3baed72d3ef7b449b20aa27c01418b359acbb93bc7c755995d45a5cd573;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf421d48896fc0d646fb48ada69a15f77a271eea39164c8f735858cc451f823b472d959cea9e59fc3d9b633bc0b35d9f786cb516ac558164e93cd4b42f137b2687995;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa30881c4c72424b926ee5678102fce40939b3a45de65cf3ecf28de714690957e026158e745a5a32475938542563a6a39a5f46e8ba438478839c66a978baaa7bd3dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9962a26aaea0c26a3595522b897e85932adfeb0a56778690f0e4b5fcf9410b84f2fb44b99a863788664489c796e0c45c667f6e372c5bda099b4b07d0e21c7f2e566e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfac92715641dde990278519d408d66121ac514086d791a2a4cb21694af9c725f7a296d60b5489ee3a2230d4996f4cd7a5a3ddcd5c4a43edfe595dabf48b5de61a85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a0198ee7a14e5b310d028555da4bbe17dd3ef521484b98dead317a5f8c9af82ab171b72d2f60365bef62619c34aada12db936172d22de4c0a5fbb95a34fd24cb7ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf511313cb9363facc0c0d44e8001bef038f00821618dd3e90322eef1fcc4896ff7a331b39d35377aa664c119a53f0b69a6b512c4c366046cd828142c4a90436c1d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h348477611cd45834c820132a4a6bccd00d5131661f4f74b5b0abc9ce4d6e36696b50bf5150426ed56beb6ea2f642fb5363155efe62b8abddac87ecf61d2c45a5033f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c172a8081e95c6f82e8c1c3d5a6a47cc984ff30d116184695af91b8c0384b4374f2f020e9bc9b8844a532fac474f1e435628654ef0aa071537a9ad6d07bb74f8a16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192914a7cf892c0251fd8cfdbb59eafe18ce7cccce50f473ebe9c7cafb9ec21234b6dc1c51f1ef3659a4cc8bffaa4ce2e5c639da3f76f303dfcc0c5036ad301d15446;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc2d15ec8a2d49f9cb4a4b70b064e7a24c8dc17ea51d8c761c2ba3390fad3c22e88ceac636fcea7e604d55d01d861c1c755bd1cd36c7f4dd66d608b814c267206c4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b298b514e4d2aef6323014e00e8d758c96b34af2a607b5ddb6dce8db9c1e7b35301675d9962097cf35306b5a2bcf117aed0a0e42cf1696bd2269d12f7830544cfd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75129eb71dc358773492497883f0811d917cdf1b588709ffddc8493c2c1b613911a317fdbe8fe203f55e7d4187f428695eb60ca96602834d97eabeb495f03fd68536;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86b4f90f0f0b0a34779227aced0049cad46ae1cfb2012c5b57f921e6a9b264238cae96faa6e8c5d44bc0f38afa281901d465b52497c6288306471dffa705cc8be614;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbe1eacf3c0f201f73ce1d5b65ae11b9f0f61cbfa3cbf0baf06794dcf485fc63df7a0a0fbf1359ba3a4d8f18b1823b9b6ea8d60bd8a7d337b8a46e9f5a4011f4c195;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0f496619c2a511bcfd35f0c45fdaa091141b43ba71c6d6d262dfb704151460d09c86d1a090be3d4c1aa3f29579722117c8dba988dcd972fe046dbe1886679bbd729;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c50ea11d18f3a6f48b7cce315c2cdc7ae6461578793b906e76cf990ed36b251739cb39da19228aedc45d79c202c30e3365bacab5aa1f4654b0d27b58ee1e0b5487b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c563baa26d9ef2129089307651839f8a452775c490e4914d3937d9e9086814a5ec93fdf805be6fc766d7982388d5f945f020324b34fe811cf0c3c2695d84cd522a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127dcca2372c4e4b26ec5ded364ed635b4ac6dba1ffed63999c4ea66e2b12932ae6b0babb9040087850eac7eaafa5890d4092f330b3cd8228badb3d74ce95193abaa0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80cab0b37ae499cb8d82c56f7f89fec3c606ca356f2dc66e5a5cb3a4d062649e88205ccb948e4f247a95cc9a79b557c14c48c5bae45568ccafb2c5ef4ede1665b237;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad162f1f92cd818847f777e48964caf5f7c710367fc1abe26aa285f02c133d8908f8cc6ba7b8defb96ec2c0eca682138e38397712b06011909731bbb66d2a2f2f065;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfe27cd43909789da0aca1b2b13757168b12200fc8a6a9c9d312f46acace427a5d0b85b1098330b6145d1e35422eb3186e85debb2712fa81d2da7f3991b8712585bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2ff77dc1e8739943a3f3254495cf25a42164a573f5bcec4b435cc9d8744e28e7ac4a62f96fa42bcac838abf66f431099a401655fe78d3fa79ee6fe44ef47c8bf27b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8ce27e5b915f289bfaf913c534d2fc085ed324c4ae215e9ae5d6ae4611143f65ab9e6aa992905f88a3ddc36d1a42a2d2fc010748e197c512a2f4cf4552a66993b7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7be62c8fc7f82fbad65bc487b65e9152f66260a24d01480c7ec2595e3a4e58ae8816e97323b01675c02400056e9c7b0c355456d3451b931211bfbafbab397c918261;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cdc998bd0779daab7a2055fb427afc7cc1783bb2dd70312b5f18eef986b1fb4b0eb94c6e1208a997ca7f3ca2452b5222294768ac639e44d59321d7ea1fcb99d5eb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d659c10d6a35dcef9d1efd52ef05bfcc4f5bad21d9003c95de33b6270f16f04be76d5de3ffed103ebd826848a626526cedb8be5303bf7aff007c81315e2ffffb85f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ad8ad249a5a1b9afecf331632d35e1c4d129f0ce0c6abd22643237621ae999492ab726d7b47843b0d02efd7c2945d892a4ff1e2e12a2ab6ce4d21c821794659f2ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9c962d4e7cc820fe6c8e5d42b82c04bf1962019e3bfa038c3b18385b166f5c2951fe8cf50a66117b4d89f63e076083ca2f08ab75471781704b27fa51768510bc9a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h325f0a8ea85cce72693223b13d99e92633281b44da4cbe5e6d7287db5ba9cb9ad247acf31c9219da471a87e6ce40abacce9dab460b10d3397dd497ee958fbfbccdcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186b6ce26d31e8d257b380241f3017242f16718618b92b08770be200621488e654f959a4beb71510c3db4cefe96af402df5424f2653b9bd503a85428947bad61d85a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9df5caa38b9439d6b20910ad76fab8b4fa8fe1abe6bccbd7be95def78205a6497b35db8fdebb9abf9edaf890479970bcfada11f9222d25945c706f62bc010783052;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83f74aad40a23c721621271da8bdbfe2c7ff99372d3df604008ec092c51fae153517dd082a5744915b338324148af320653ad0f1abc3202178f85b94702ac1882401;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47af79e83b8190744a683f0d37d745871bdb0343fe411d32ed9c13c34bf3da5709af83238e11e3ca1ae66c3418f6bb06fa68dd03c2befed83712115740069ce42cee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6e7b13a8d870f0f2228647146554e5bc2753f61e64d50192016e5cda754e8b1216abded88cc0848cb0a21ba947e2feaf53280ad72554ae6593a77b9c204db641908;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191883e82725a19638e9de81221b847e6e688319e0163732a8b8ce2d26952f315356bd994b664cac8bf36b9f220f095a7df5971e439c5b796cac36fd9c6ef7baa514f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f70f8669feedd738f2af62d956707f604e505da09f2683ccbe87b94d374bc00e1530b0d168ec7f6ba1ef6b57defe836ddd11bee1ba89147d7826b6c9256aa8675427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e9deee6faa16fda097a168511c1d8aefa3a7ecb3a024a82ebb09c7afa3f803476e412c5582c20cf83705064659dd4cda0d1257a87bd71d854bea6a8c63cc755f932;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5606a90910fde2878a7148a940fa9ae078daef9993e35834b5751f1b8ced6214ba65437cb196f757b7e4b4daf7fea1f896abe4e9c90763a8ef09f072d177831441c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc557d294aecd6808a50318ec95c9dbba5b06f510528b81c9deb5c5d8e3e157d4410cb9ed56052b7b49e047d20f20e3e82c418cc66ac2f87507f2bab58ae2b093122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afb584095ef61a8d3530ee1cb8ef4bc074dc8ff800b6bf9911587a9ce31017f4d3fedf917119acff8011c7fee2dc33418fdb10ae127836609f6bfdfa4d652f83602a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118cdb7cc01e9db4b24111c49f841d0946c7ccff3d3473f16eb796b144451696cedff9b943b0dbaa8ddeae83273ce00669174ec12ee6e3fb31a2bac683b3a18920e79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11986e152224e339fdac8a831b37d07647662cb1fb2e7c80544bc6d3a3dc001b112e5270015b1b3ff31c22750251242bc9f0615a821353ab6f651f696cf4b6c3ae536;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1888dc031466abfe774dccdaf8576038e8088211a8dd0f086d9db93705539b3f944eed1402e2d0ae958997f601f38b868285fcbf9cd0f212941a675399f82e6bdac37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19dd1de206bd1940f157e4d152888d2951764a12b8a598569d631a45fc82df928b7a800bfb4a743e096213b6428a8cb760a1ec2a8e11871e7248551acdf06c8392495;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1414fcec46ccba332bc83213ccbc2cf5bbe2664951b48abb703890dd9400b08f9c4b8087caa629559d58047f78700d51368aab33316f8421c0eaf0ad166b0b4a8d556;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h945259e8689c59eddf292263841814a3e7e887ea4f1740d39f0eedc48e88b0780a22507e81e3d3c619afd431602e9181f3a5363ccb3e901c447d5481c53fc7e164fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181c08ba2a2578dcc74f20f4938960b0ac28d003e3bdee24d036132ecaf6a18012470eacd73f8c89454c4212aefde978fb46a403ea3bed533683a4393aac732ecf69b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1470b5c8279df447a6a78efd2534a8296219a8c359fbd8a9af4eedcbd8f87f8b60e30b992a500d338a835e5afea90ee26265058d96c7f699a5e483ed044baebb6f1b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86dbb567174a7d7e9bc7df712cd6e8a32d7e327e07949dc58585d1d7cb262507cfe61229b953fc2da9827125bc766d274574497a109e918a5ff350a8501a59504ae7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28c7b76df76b1b1f83d1f54ef684a55e2dd847a03e959d317f4e04fc7d59075af50c797f735e0fe5cb7631714a1b8cd44f92b2d761e092a181667508d3be4a4140b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d25bd53ad0cef70be31b231012a4365ae0c01c851142a3c382123bdf4a3adddefbe8026990783c5dd8982ecc7d8a58ede2f411c4f6b3eb42e626fb4dc5cde8cb1c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ada9564217c310b2181fca1739b98b3f00e34935a918800bac9deb7cd1bf9423626179c4066c92eb7e5b62e2889a668b8081b375a4eb69152162ef74e1e43b751dc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf810516a128efb1660db0d376e23f55a8a26d6b18c95d929f71f921276bb2ebfbed671125626fc603c3c770c92249b87d7320d19691a30a924da553176f44699bec8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h336c058620fdb1ced65c39eb4536a35250506b6bfd8208752a1322d57104da034606b88a697144a8669731c21c99c11509c7c65dc68a8acaa1f0b425ae0eaa736f0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94e7039c55ed4fa470759f5db0180c747924c63c64dc739959f963c84cff0befd34a5c70136439d4146fb43b542573f08fe82bb02dbdbf8de2ebf1d1a63b6d44ee5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149c8047571920cc21b663f970a87caf02b6a64879550cae3a1f2dd29f15fe77b9191722cc6392483395b74fc6d216cc4da433d38a89b44b8dbc9447fd7bd408732c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ff2bf5a930d6e45d91c1cf08f3f476beccc9e17b7d65df2dc3d370c0f55a65679aa936d1db8780e29a8d38877d51939eb3d3a4b68dccee1e31f480629c68378215;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b390d3551c3afe7f69a1f0edd2c055b6bb8daf0abe523a30f0cec39553a00fd655a5039ced5ee0191df0416acf62f3d4951bf58ae0df1594c14d505e349e2f6e04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc69144154e913845a0a8c2d970a2a23494994f6b43cd573ac7a012055dd92110afdbc94a3f854c3d4284ae25fbee211f817929ff0c2bbb7086d7633ac0a7b48c324;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18719418549f305e9b5cbd52c5b75d0503c9acccb8c1f1a0a18ca7cb208168bc066c336fa3f64103764ee79df2396e05b4ce9545740e88f688879dfd8256b84ae1e64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd01611fa80bb96fcfea646b0692fb26010dbd060dfc0bda3662300fb3dc19a0302216fd0ec586b38a1030fcf5e78cd9ea69744ff58eccecc74c15afa9254353c620;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138ea132ce48571c0f6b8ed4bb01d427301f34efd61eb3e13ad7f59d53b1b9982c02901a92078ce01d42a334edbf28f8b738b7b1aca793b5baefa0c7bb75e95a8b92c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7144aef1fb2c101856a36be5ec031c82a88af3001f0ae3e76777cb2653e2a2626c650891424b055b28cffe26f14568542dabe5e9c98278821875f2e46b83420ab61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1364f3db32198af7ba87b33e2b610c69567611d040527bd2938df9504b5a85334752fa35529495d73972835b144a628a1c56b6f9241e699dec172e062d67082fbfd69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f71a56fddae18212d7ee82e3982ebed8206db8083f49de0b86b9ff92ba746aa4ae33367ef0075d76fc86619024ea41ca05a1c11fbfe1d2378509a8e09b915f166857;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f04d49acfb2b31691fe6f855257c5005344487e5cb5a11ecd7b530392765587666c7c7eae5c414654564bb3805fe5523b4389453d5f4dc3c66dea7dde11c6bda53f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cad63e842e6ee60d0edac47a653b1bf4fda1c03e68a37c39c3210f5b75da3ebcbe181e8698e62200397a6987ae29c70f5abb3a795bd4b08183a0b306f632c5af434e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cbdcf04460d921edaacc96ad8f66dcb73565e4e55e852c4928f05d6b8aec4eaa0be7613fe55e9d7a5593debb4ab2120317183e445327eb2c1fb117b23880c42021c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa133e463c00b6ebf5c54d2ea33e1350298bfe85cc2a0afd6a3a2758f584f8e446119b40bfe68952668707bd4b199db11824ef7eee5699b22e63072c21b3d6b8dc38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19dd573357802eca44a9b3e541df15e1bdf31205c0756fbfbbdf8a539c0460a1952719c0707ba4e23933ca33f01ebcba6218cd9b310873038e041900ce00c8cf4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182ec8c479f28e219f1302fa6be3df1b8e19c72c9ba2602788c28fb692cbb6b3d7cbc56854815329064e61208884bec4c8d4ba393e272918529de961e29a353dd5bbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he65fade981e05dcd71469cee9f71937543ce3138b7fedb78b86c55a77e3010e366e5fcd154dd5a319a01199bdc6e55ae9b3029cdad3b2d6f6e8452713bb9d060cea9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3193907dd5de6da610046a595a3ffd8477c73e0862285222c68095a9e23018e392516fd454bb5cb3dd893be4d5e5ca0968a2eff51328b53c0ec2025250463d22b97e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea6dc073d0711e5b25afc61fb43972940aa9419e474bcd962a0fd4c3c21a2ae776bcef77dd12da0207f18ccc793b6fd6ab8500f4e61ad4ab1ee2aa5e27c2a9505476;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcce779a86ade5e3b65490256a7c73a7fb4b9473da60554f134330322fc6dde0ea63cf2d05c529c201901757b85e0103097a93bab200ee979a5fdc0eae0e7240527af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3507c6c4e79b9a44084c6c891efb826bc7c942f10895a07ca9f906398eb69f0a21cc03af7fc374e11cbfe79911c8f89253c15730a7f2453cda245799c9fde327e59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16de1ce27795cda2b727c10a07e25b95931069422bf2e096417198c8cace8791873ca85d9fdf55453d84400f35273125b99ff446b797cb807b802fd86e7c1482f4fe8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6693928a7427c601c120625bb9545877fab24ed8dea2c315831d4272d4359c57ef11f9d0de6985e90cd15090384d4b3aca980e7601970559962c9022167fea90c9ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c30952539194f1b1a2d7b1c36306001307722caa3cc8478871042596808026b99b80f99c507e50c87a6b4a40b858f3735af1e1cea88bbea543179d42f4caac66566d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9def11a9dbe2f426be8a8fbdcc7156c69aadf072e6ee7bff90254807ae306f4a4bb2456da9a48c01430192f757dec041cbbeef876c8a40cb9a6532c3ca45d7df147;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdcf6f644d9a3b55456f7ee84a32d5bd1f19981ece8edd197fc7e3f7a3d3b7523c891d086f60830a3b26dc8b6519789c7c7f696d3bfbd1333911a22b0e518aa1a0472;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e350455b8a6447b04bfa4ab023bfa7d8f11de667e4699f70d692747c643f722434bdf278284829be85bf7318f6fe84f910cc8a52f5b73446220eafc6228d8296024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5ad8c6cf2d324347724747d4920139a0cd8a848552ff681a3179fe5804cbea32a331b2b20b32f8cd7de7b3e105c8e56472dd075574707dad441798e301518d4e56b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192b9d19a29cddd9f2860fcc2cf4208a57212f2f58793f1c5e67c71b264f45198600e38ef7d7a6607d8c14195aba6d797056b6dc40af091d1f286a3fee2773950c81c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h197aa45a5ae1929567b5da2d802c933a5ea4b6a874c92a6d6219c99b765897d8392ca955533a650a8b13d94f85068475c5848e9a7adb589e9361ecc97793f88338c28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b344413fd89b276c632d8a16e75291f6b83cfe54828daed52367efe6e3d58f223035f10ba094c09e0346129429c0f86fa69c180ce2e89bb3497ce0f6bc42b52f07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9dc7ea4c7c7af008090642aa254317f169daf31178901112e10da0c5d4d440fcb9738154e5e84f82ff7016e6af9cafe733a55a17ef87b2ac212757ef5befb4909ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106db0065f022ea03d893ab616afaca89c3c31a435fa69417ecbaef2376efcea7a8a8f761ecff03a7dea5a772c6eac843527aff0f51b9b4e7d62e3a95a283ab107e9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ae2c8dfd3ef882e93bc7fa52c6a085f437dc9fce06ee8aefe7557c40b425a92bfe527055aeaa47dc79220e322d23ef4df0ab7db8f7ab162f53d60ccdf9a0d3373c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b09cbd990f24ba77992f57b1ccc4dd1e04f0aec1fa05f73660fc27c95c3d660da54480c7b84b0fef794c0576483f2a3ffb8c05490dcfba8cdabdb75c0f27a19f1be8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105f7e4ca55bf4f5aad539e89b44e2a2d3bd512acf8b9e1a3cf77bf4b5b250c1e3c30a3c3ed7a401e9273a892801d87c6a04726a9ba1bc30a5e8dc7e31d6aa6ae7594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2d43a93b0819e79ad4d4ed96d806e0b22256df02642ffc95b7ec4779b86e5cff17f5791cc8b168a82d273ca0ed347e642e6515592a725ca483303d359f387504bc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aac1cb18b9d8ab9c5c322fdc3393b4f367a27d8c3b726f6162f472bf20f66b23d0c4804832c81785ecb2dfd66c34d973c42e09f8802f39b7d37fb751dc842a038718;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147d46c88162402bfb2cb9e33cfd0a6b57cfbe15aff5bd0dfd764e55ca8a93de06bcc77eeecc2d43e5bca2104521a249d54d1c5c9c13572ef224874cd15b7fe29c9af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ac354f4178fb9237b5cce9943b18c06df52e9b082926d9e880298a6ce95792fc4fab3d4f76a25c8f23a5735de1b2b686e2f7adaee6d07898d9e6c78e56f0ca8936a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a989b7b6118e86985118588603c96c3823270333a6c70a87742470c7e9195e260ac24c22038d7d1706f2ddb08003252f688e1ef535d755147b31fb83843ac0ea7360;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f79a31994ebb5ccc3851ba024d032d9d8117f9f8a20ab61cadfde245c67b10d063ed56084f8dd2fb590e4077eac41dfa500d439f1a62a0094ee0751fd459268a556;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95e11f8d2865cdd86556b1133311096d4708909ec2118c18291bc90392c63df1dd3af9c413f686f8745b012db3a26cf99941db407e6b4109b27cf3e36fe86f143921;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1c7b0c6beca441932a77e4094fc82e0c4ded3c490a4108f0cbc871d1345439b7a5393a1a38aac883ebe70056b90d0907f6632765c07ee1871e336073eb12ad505d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150ff36e7c3edae1ec9e4fc49d22068787e2f1695f06b4dcd1e5536b94322480061a123440ab11a785bd5529b9335c1be4e87bdf270d45ddcd7ed2a77af27f212efd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf322aaf9d7ced2bdcdd2a1420e9028d4f4fd4a0beeb47a4b2ba4bbffc65cf9f717da4ebe9cf4cfb4191e7039e18869763745f0b50ee1f8dea14c4b9bb5ecb8eabf91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c8a36a221802644cb6e276f07a9f504aebcea5414b4e467b74fcd72fdd77485a596f8204bef1e5f98ed687780161869e8d7aac71871afbb66aa48dee7fe01aea4152;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc917af44ad98066dbae624b2d42202ad790780364161637079226af3380be469feaa2ff6a20618a0fd440ab8145c09e246da5199f9ca0a9f37d258a0e5155b1714e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57377ff6676aaf64bd9b45a2a4989d3cc65ca472bf44e5d3afcc8c957719333faf3d51fd9f49034241cc7a3277c015db3b665ffcc2acaea636c40a17d8971cb416aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4191011a0f7a9ac9eeb3a61c008bd4c80f14f8e02d5d11c021edc2f7c0d14354b839d91763ee3de0aa53851100331a7a9871fe4058a6ce8572f2df98d6a8cef9180;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdf96d879d8d9a635059b412c735da69941ee7ca14fbd7c3ee15fcc43e52de753b2cab03c4b15e3a1dcf7a9fa67c8eefb277c9b14c1047a493cc03e96a5144a86c8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8847a290ccdbca99df2fd4ce9e819ab84e7a9279e7786f92a272134d38fb62040aaa5a7215ca8aceeb264b59b24695760c3ab35c9b2b52482b1bdc196bf2eea5760;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135471d3d29e0ccc596175990a5e9177d1ca25d3b27bc8aeaeebcb595acbb465f376aa571f2d616e80f76461a3baeb0a265c3a8c4378be1af3c192183636457d5939a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d22f00bca75103ce1c432387111bbda75e69161cab2975e58e5f6be8c5d4b8cd86cd3587ac0a14488a6d784b830bcf6c255d38f9dd8075643ad2b8055a3626f9403a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6b7cf691b232b8a4c00a8f07c07412a5c95a9915eca2faa29d95dfb5d5fa9e464e31f06b9ae91e741a29fc9baf7b872f183d11ca0cb37fb80944d7ee7e226824761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3b52710fd907ae0b1873bf299b873c588755512a339fae1f7d7ee491882f4c5d605fb091e3af146fbbf6cfc6d0a724177ade12647df6b3ae7713f831c6c928f5856;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e434f2d20c0e6f10afc6949628bc5fe96e0d43e54ae81ed33a073dc9e7032cc99362cfa919cb179201fef128106dcc91b63cf0dc909514fccf0fa8c44817f94333a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2909dbb130fb4eb18d8091a18ed4a7dd9debbe2babffcc82a5e977c611a5c2dabf9a3e714dd1ac0f6539bd7b96c8b4af8f7fda9990aabf49a794a0e1f8afea085fd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa5d3cf75900a79eab96010c21c95b17000f4910f8f6b7c39c1cef31dc5bccec3ed74bd43651bba36a715c78714532fa56e22b06ffa9ac81ade85782d063359edb0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b81f45e6090b3ba8c0cd98ef613ecd9eb1c9cda1a90970c9986b0cb05c4cbf99f95312cee35bbb86b13a4f531a7190e0695913fc29d5b75b2b8ea1ba9647dac885d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1202d046f8d1b09505ca029067c00e620bc99ac897ba2e81f0326ec6099ccea74ccdfba47be8cd364864cd3522e294754a7bff48c180a4d0ee14b1f77099848d2d491;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec16787e31f9c42aa8747e279b9c82d0e9cfbf34020c1c63e2bd6f3891acd5a9612ad8efba3c7d525e82cab1fb6f3ed3cfb1fe16d79404e3addc981789895d1eeaad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ae5034f62405ac89ab9fa28ff205d1d646983a5c968a26df3e64f6273d8e3d3be26184ea9ff02bf91c9ec2e69d316a0efaf4e61df5314bd329618ee322d8b40016a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6558b85007d5f00248e261440a1ad8a43050c6b6cf0b4b6139e03588987cdc5d6dbbc3ae571f41607f9a9f958fec7e25d2afeae74860287642fc05aa31c7bcd1eaf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa1ea2051d1f80cd82ea9f772d83ec3a621ffad6b4242b5ea033f89fe07a3867a59bcace98a1236e3d09abe4f0a0c8cf0cf8333a8f100db51d5743531b388234ee6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee9526a711eccd22f641981ff52d162ae41232f8279416cf0b793b60bc5c2411360a5dd377ff9cbfe49b6ae45addfe7a1d2a5ff5fe009dd3a5fb8e91bf0fbe078450;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5741e9d79f3332bbf382c8b893cc1d076753fb9d9b097c987698c1ebf3d8993415c7a2881a91896f8d5c8c1ea2c2f6801792eb6bad72b0484d7ca4af500c9a5b1f5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9efe48ce0c52f83fa45823a32799f310b3fe5193ccd71ffd8e1962d27f967e48149ec471906872be868669a79703acb3c5c0a195f34766b36d05355781499a58fcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc87750a1172614daff117f2dd082579d6cabd578dbfe2ca13ec10a5290b82722c41c45ca47a7844901d66a9e77cf19bddc235c9c6cc8f9493b65de5420848ae08670;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf867847860f059ccb20e1ac02879f29c52ac4fb0d000afbfff2cd34cfc4b73c364db8921be2329f4baf870324a0cec9e6b0af7f8571bf08b86249b8012d8960f98c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1427a8e135b2c328e4d4ca68f74ddc95765b871ce17be743076949c7a4ae41bea84bddf3ee49c5551500d6b3aefb9c49d7bcd6908a85df9fbd628f2ba99a4ed2bb8be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec9b763998f7910fc6150f27b0b312e50072d8240e1425fdd5b4bcba8bee8354bc5afd87860f64ffe1f252e719a2b1c94e30f5d4440f1f4a074db2c055f20ad41762;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he89c91d3d5e401bf4f6491019d6c19ed19c61b62fd3f322818940ee8844288d07ad949fd5277907ef2b9d944dafb994da4910aefe034d3fc289ecd008fd51e577cca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e4b6b4c02a4b551617925df9d33a8616a217de77fdfc623c5f7ca0bc49ade37326e37fb587196f285f3305222228042c584625ce6e7811bf0a70de4c0be30146a69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118b278a9361084074b8a77aa6af3d8b6e2906f894bf9c1f555832f06e77a566f07ac5be187cc9fe3f410fe88ca2e288634ed1b4bcc0725a61606d6e817a33441a3cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113d6351842498865607292694f4230037f6f8ba17a0e4508844f38f656194dd4389fd2bf9a08afad22c333e4ee5fd398c27ac94101f9835a7c316174abf1b060299c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb67f8e12681ca84538c5da1a5e7162f956788a804a711a7f03e58ca0ef503b5769804e2c9c8e3f4c1fae2f947d4a7d12a7e108f2326ae1e5c55d8fa3c221f2b1dac1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f44ea89caa1f83e54250bf56c0f49da2079fe334fcad4a414cdfd693285875efe7dce5d881ad7a5d148204a641f1bb2c0e52051e5e3c75d831bfcfee08c8b22cbe5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46eb11436673e72707cf3ede04e79206549c8f894b4fa8687f119ac6ae5c48810d03ca971778300f97329192a63738be84c575da3e523d6a69b6dccfb0a64bf164a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f761c644b29a76f6dedbf14aebe980e6ccd92090191c43345b1b50ff1e63bb1f43ea6a6bdb6a2f0bf0e99c83da20e0a8f95c15aaccc7916c41ebd2b765e508fe6030;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bd5b8540b45d9db04d460b1ba378118331dc44d122bb828efe4ba7e6461318e89cfe3d0ff464a2697ae97d5c26f49d792dda21716e347a2c31de147d78c931e7f1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h488fe7d450f88a512f7cf78b2bf53f9f8aa70862ff231a6dc1c5828b5715c808fae0681f990ba84f454a783617549bb6a27720bc911d590202a3701dc77a6f2215a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4a3e88c0ca32590247d66fbbd19de5b0a11cc9ea7451f524badf8d7b373fcf69c64617354090e26d0b5530b0b1051a283ff1492533f2fdb70a45d7fc0e8d9f1a435;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134bbc01dc5e8a45ac4730e41ff176095b1cffeb05e67a549072fcbcea100d9e767b535285dc10145310da5942896872e266856d56319a6d0efd6c03a59e5ec3205d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e734a669e2bc63d9ea96008861f1a35591f0ae1255cc689c32998bc34434f42e6d1dc3edcc092fbd260a635ff6646bb26627c6ce8880086dbc2202c8ecf9864da0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aacf45323fcc758428bc52414c52590fb90ddd309c4bacc82f1dfe2ad2afc317380ce5233304f815a98691bafdc9f4a119c621cdb27e20762d9d4bb11ee8aef534e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb2c92248c8fdc17e0266eea1d8746418b5b07fcdc8009daf6bac4c7d61dbc34cb803c374c28d09380edaa911d628d3dbd46721adfa24de61a80fbc8309155e8d91a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h232edc27afa8a825339f8c4c1880ca987a0143761fd70956ce13150a097ea7c355fe009f313318cf3c25de9ad9b866d4cf4f5fba42e460dbd6cd7e309351235e0222;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b883288486dd003e744d176c41e081906544313c34099e36f61aaf7ba67efbf3121dbf560916ef26e7667a2d865298fab709581b054ff44ecf1db2f3a9178fd0d11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171d4b2044f60153b84ac65efb5dc99bed8193b7aa39b9c37e0068ca2122ce1fb5c23bc57f90b99a7fc6be823f7a70bb109a612005ecccca8802a852ad8de995caaba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h92b715f0c9fc269664a1f548f11fa0211fbf268073bd6bfe1f14f641e9b90d8aa0165e03570da93dadae9d7b35aa08eb70d0e1218ff561ecfd807a1a41008fd30ba1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h531d7ac3bb3cc2866d4185d08162b9316e64b490e324af898eca43b3d1e8756b4a1fbc444296db5e4f23e53cbb8f520955ffff4872db760875c54a75bdd5371bde48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4b80486fbcef20f57726f36e1b1bd295da3dba1c5793a048913d1a812af536bf61f518d58b8c724ec0ebbfec5679037a730ea55aa4ff853953f824c0a4c951f4070;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfcc182d5e456dc45ecb2ed4718dfee4213453737eee875bd2786a57c0ec9efda6810ce11338c04dc410b0ba97286cf590fe0cf35f91c86b2a35f899cb36707b0cb0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb091aa24f1a8ce830de38ed97c2afcffea0ed3926e59f2f7b1877ee5925050276d76bdd3503dab9d31faa551c850a1b297f2f71790785cfa90237e103c3896ac6fbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9610d2f216e677f991dabf9f6884eeaf34f13832d735774df00f701d3796ea6558da5070de579c8a2b867d516b8c5c0afce1f2c2cb62199162b47ece9edb092b5b26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8130deb5c478c33712ad61bf6cf07174c5cdca6439bd68e29e481d04dfa18e229064e5e1bfa7d63b41be12dcc2cf88b075f2ccef857936a692e12fda1382350f93bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe8458cef9e5efbb02389159aa3b6e487974a29f2956710ed1a7a2dcff7d4c7f09209b675116124f9801c19b4ff29e9e2ba0acf84d92f9af23c981cae2018a907cbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fe67f986b13321918e8738abb19c41e0b3595569965eae8b9f8c273c37d68e0721620d201611db20648dc545c3f9e9f3c60d96993f06257738119b6e196e62f7a94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd67746a32402786d4940a6aed93c3ffff747c51a34b7f320847545b346a8d3fa6f222e21acaca4689d306cbbabf40c1958a6d688d77c4f054190f152fdaf93c65570;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea938e325d857a62c9fb1e726d4f2c60af402fcc146b2124f99e1945077d31e28d98390b49af30ae148f09e34432a30d142343b7a5aee9706b2f30d593867fca3048;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8857c83a2821dc6619e5e56604d0003c8aee5d7374fb9950d1aaafef30b4b6ea3419b93b9e8d80d10f3b97f5e5aee271c87f5ca7e7ecfa3f38e555b867d78241e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107cd5d0063ff5f7c9ab4e2f041972eae6d02290b59fe966d54593f7463c2bebf807aeea6071291b26fe64e9a4ffe71a8b2788860266a1cc374e67ee167e1d9a7f115;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e2d1b8604c2c7d78377574ed3be287bf5bbc2ce574420a9ddf4f82ec5ec22a055bc0d5f788451499aaf96d41a0becbff700fe3a78e32ba7e0be88a42bffdfaafcf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e20819891bca8c3a0861952375b3090151157c9a209e0da514205d61742ee1ab8c2cdce68a0726742c143a17d8451cf45b7a20724369e232b4e888f786d184d23d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da9e051a5fb0a599a382cf16b30fa18e0334a19621179f9d0c79a9f3fc8fe027df852d678d216adc928a284b4cce4603652deb577d6790b1107f3740b6cc52faa435;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had81a743d51506ba107e4ba4e8a4bf6487ee781c2bd9d790e753b8076ca9bfb62044ea0ef649618c55fc34e3c783bbd01c762a44f7d95a7cf5e486bcdfdc5861baf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd1f9685462b5839e7b876d27432c3249b7e9400b6c47c2ddc0ed239d01db14cb8c6e029d98f3ab0788381c489519f06c376131923764ed338bacd50ecc600257ee6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1209649aea68d9444fce9509624db052ae9349352b60ffcfbf4f25ec22cff02543142a4dd2cab388dc1e9d4bbfb9e93ac5d3d4d0424ad5495cd36b0491f5ecae34293;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115f397e2415019863a39c2e109e081aaec444e4912c43d36d50de905ad3a8d8cf27eb4f9d748b7da3c91f3a319dc69f2796cb1ba959d5747fc00ad45407a47dc1f86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c73aae706e2a426a437749c445d3074022a8373e196bcf695f85fe25a456d4d0fdd216f35bde17469667016f15a23e4e6d2ca1c1e6e34ccaefa08f713970a94c5aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c06698b308a76d82f385591cc31e93846121e8d25c17435b69ae4a6750fb742a86b87894babe4921241bc9e117c06ad5945e8f15faeef7643464ba83b01b47782f60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5569b02cb3974a833ea7f950eea52b74dbffc818706342c476bb1156489a901914733f6b4d61a29c0c439de98fd11ef01345c8d313502e372f415838a2c3639da05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1f2e0b7b00ee7af058dc35ac11c801c51d4ceb188ca958fd66d4d9a66151391c88ebee67fce82474b300dbf974517da6f4064f42e82474878e366daf7979d921ac8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191dfed06391c14a9ab08d5dcc9832b2ad5c201b6d2317285e1e6c19ae34da771494147aa77faf0f3cdf21565141f7261c2e917730bc5263d6975c1e8fc966e6d3af3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cda2ba30e080cbea420d0972761c1fc89c99adb003589cdf60451b034fe03452de020067d069ae73e508d4852dcd4705a025e7248a1b760168387ee4a40d9a911c64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf291c5761847dec3728adbd096e9c48a99ada7c4635322204561d2f2866c64aaa60735e8837267b7f8afb2ea833d615c3dcf5ac2fef6eada7c5a049d9fe110b2f94f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0495cd1234dead7209db23189df08a30896815241ad5985e3638304305879977dca26a69212d65f16b662603430cb5eecd4186a62716b5edd74e34f6b47b53ce782;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c2b956b9bc6b1b8e35c2506953bc03303eac4920944fb60b137544668752bd3dc421893b138db20b78fe7519a343ca2031b960a2f4b62b9a0067ee6bb992e96fbd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1774cd0a6a5fe9bcbe9848dc886eb9ba4f8f71128add0b9b140afee6e3d9bef7843f22d4d17bb5968e7f916c4c0fa7b69e4296cf53888b5c9a5409fc4124897f8ee2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bb9a47d46cae7a17a28a3ecdaf59d2b04efb34871a3815f75363b0b4c391aacb213b466fe271b1a1d37a0506f8f58ff1ebaea48d0344989bc30178cc037c59e0356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d58aa23b0c80b5dd5f5398ea0baa341c4f179d49fe66793f5e1a77318fe71fca37761918ff98f28eb79df015e01f68ead40f75eb1a9ad8a92298e753ce78b368857;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87aa2ce822a0935c60397f7964d5974b38b1ac0d875d798e44d163cd8df99f6c28e620bc4a3edf6da03aa7a225b9d8e425b85850fc5a90f2199cc51a9a1b13a22b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af6fc3724fb15ed3092bd4cf64e6b3b38d9ed71b845891cd802024b02fca50684054ab874ad6ac5924c62f35b451b9a05def06398413a923adddc538dbacfa3643e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95b61dcfa49acd498cb4d99d16a92329f018d1fa13f0482fd27a01856443d4d4bbc61477431ba0636277be74ae2b3aca7e6ce558850a04488614317c15cc8e44aa21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d1b7370fbf36d32f293ddb3b4bcfd402c7b13ee5f5bb06a21239712ccb4c9de16f47e211f111d06065206b3496159e2c2bd7aab687a3df28b76eaad6698db092d9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a73d0c5aed46ff4d9fb9e8cfa192c55f0e8ab30845f33e40502b91ffee61c6b311fff408be0b76f17247f18c400af90f5c47e17d2ca8bf827470d8a14b75d3ddc70a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1749587f0893f25bd61fc7286f0e6836e297ec2b8460d36b9a7fd401f9aa6ddf57f8831868fa5207499696b1fe594ede6df68d303c7fc29c355f8e27144327c7c1401;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb9f24870c64d7614bfa137d37a209e25f817b7f849869a1bee953643db9bf9ef6df359fdc21f8ed32ac5a7e33a42087c87dd179b5d93165758b5066588f8ca7fb80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1533d8028e8f01f3234978cf8e5ad343401226cf70bcf54fe089ba16198d3f24113595c05833784e07b8ea8ae0baca4a59b181beb30e99ea382074ed349369c8b51ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h446cc7fec479c589e32997094969b98791aa1c888aad259b7b951d2af9588c85dd1c90ae579e6bfe2f913527c4db49cf4395cb40a786b0777739bdb2fc1f2c7b0053;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167dcbc6db680c4ca73b8cb11ab6b1b18f776b76dfcde34010b807068644b13f30e11a0b006a5c171abb379babc8b91151cbc12158a8ab86c8e605b3b199cdbfa712a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c3d3dee1d8eae24590f58a4244d298f8fdaf6771a225919bd4444386bac660c0dc370f501e5a68b948bebefaa0f54efe730441c32af050f0522ea0800e36c26f002;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c0b69ac3bbe835f56997c7bce0f984786b659fc5ff4e22b8583c3732ce78e185bd9e1a42fc64eedb70edf124468d07c2a15c73f313b3283e0a37482219eea1f9843;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b36dbe519a8dc2e98365e7a9f6c7a8d980b27d731332c2e91b39dd0e993c1da8000ba7113d6d328f402c1be6d0df3dc6cfc300ad15f6e6f597f8174acc78ab2e4f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h930fcc1e8d69603be0b3ae1c03e9df371191e26b9698be4b4b5631937030ac5b56bd7be9d952db9bf23b6689a5c2efaeb1cdbedb8588e1676b63b6a3475974c70e11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d7641bccf6319c537dc29186dd0e3d5b2896f9bf719c451dd6ce08658ccc6cdd069fd49ba735b86e267a0fb2f94b0c997ceddabce389f058be29c67f88e9ddd467d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fbb02cdb84428e4c6716d2043e138f061904c1d1abfa96bd2743404d54464edec2e0b9b72e0befc5cbdc416d748867cdc9d053c26818b75639619c1d53ecea6828d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f5879f209e0802f82af3f6b0e50a55c150dd8b2a5c6e993d6e416dd3cc491a3c9a5cba621b77fde772b12ce1a5af053d03571c471c1cda1b7d24232a3a7f528a30f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38bdbd2afab35ddaa2dc268c0ce3bca560eb9f7cb42429c22b9344cf36fb49a73fb67df64a4b43f140ab81d6ebb78f990c834b212799c258106a3e4e1f5978d043c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h602eb957b003a19ac3af4c4e023caf5c38229bf30a53b8cd8bc6520b2b754b08548f666c38cff88e20ea9d3772cd0683f285d12effb893a656ed1e1e56769348e9a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b84201c8a15f119033496d9d1e4dcec38fc716c32245dad8825f5af7b4ea3d2e2a29057dfdcb94da3d0f87fc5854b187d4724dc8b917dfaea09d3b4006f61d8a8274;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heafa219196228f9fc7b715ca92151746a7814d6b60f81a8aa72a6089edd225ce5bf72bbe4df6d4e86badc23c478a03d4717439652c5001e78418040bc25f33ab393a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f6642026d5c005a17f528c96d939078912fb19b606204fb298abb0e4119c49835d6bf5ad5233029d3090554364b5a7886752e2843327c21dba381726d54416de16f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1197f71c3950112efab84b1c976e46381bbd2b5a242768a74c244a7155e226770690028e8d9b0bed8d0a68a247ed996f122dea8441ba8fcb0a04dd0ccdf935bd5ae4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45f1e6ada55ef56eb178b746930c1527bd8978446379db80c3b2eeca8c848773c7e3b4d185369ae890bdbcbe69c29e3d08f91bf617bd8f9973d9f883d2b5c7d43132;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141072bd4c27d54326a3c201e0f11b7526f97fff34f57afd908e8fc4d98affeedc65a4ee8843dfce735f8e49b73afb235b92a3c172d19ffc1c9b10833c603968438c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fa10de58ef396b5e7481ccf30cff9c37c29ece234883a90dd93670b123ba59288ae9c7ae3b82ddfe80772ae20f840b9959c4d1a352f02a40852d85a39536c0e6ac0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2a03831d408f1a980feaa7ccc8dfcda08c3b1170906873e2fa0bb9fb711345bd92284a38b2f39175f5deec47676f70f817bc6bc99d875a646e58cbd92c14d34719e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8757c1c013f33ca699921320a044c29347320d2cac6ad903a9a0b0ec8cb24cb111b67094ae07790a7fe29b5986d3eeefe71d47adcafd9961ee8b601c85711b663f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc858058aaf40c7d1edb59d609beb0cc6d95141d55960a3bb773e32bd39bcd351a81648e4328c29cb756a478b14db76129dbb8ff4c627438520b30e4fed78889a6e76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45e7e369163606f13f1c9829be5c7e98d5d0cdca61466e19f845ba8d09424a39786f22f7499850152adfe4392051885875ca2fcdce600e11aa7f65feeee291e09963;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea28de60a19c404e8ca393905bfee82140b96ad238e0abb34d5d6993348ec4244a57ba9c580a3b15af8042416bf04bb5f5a26b5d3819be609f7f6f779a18a9e3cca2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4532d1a74aafad6751859be140c9e3a9979620f6e26c7d883af9330213e5773ddd0bffbae10f2da0e2a591d6394e379e83b7b7db0165ace634df37e4349083321f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcab50c4f36eb2be21c1c758809a170d1922afc5c12d61389ceafe260e53e5cf81b1a5a2c9acc04cba8cf56872d2b26600388867f6e68a1c108a0979bbe12eee2afe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcac7456ff305f7ec7a82c16f1dec94c70376946591feda4d2e68d5e4ca25722eb70b58695d4775b5145ac2cecdda3da637284a6d04125317b69253618e23acea5909;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc5ad74c9811577e3a3b29bb14cd153a2e24d2f5c00fd94f5ab8010a4e4bb497979ab8005af0cd4a0447f4db3fcf178275bd38174f454ba113ca5f6996328d3de835;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee1a7300f931155fe7cc3d3d09db816b13281358a9b7e32bd696ce611abc68134ccb9f6b946c4b7364675c9fe248e84eafdcfc9d69d71cf80bc496f965002d357ecb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5cb813dcbb1a57fcdd81cadaa2646cb52a5c0ca73af1c10d7c031f5eef763d7de572153e77cafa051b308a3d7843657d4cb8d101298c8f39eab4676d5aefaa7bafd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fe342e732f18673e8e47a1b7c997a18303ff91903916df908d963280a528f17b910dc4047db55f492da304039b5da6960adb52b55f2522e66e197258504eb90c00a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bdc68986febc6b6c61f818f0a251a72004f6c0038367d004ec2ea310923be2b450805b905fa3a90afd94b84988e148c46638eb2d3f38543d49e9d738e7ace9dd15aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6025945aa03731f1e097723b5ebc4f6c92a9577d7dc041a81205ab6d2dc41e5697081b671d62dd73860dbd384f53269f1ca844ac23a91276daac4ce965c946c45d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17059ca480249036cb9a85bf71b1203f0f4d1937b425a4fbb3eb63e31b332870b624a921de155e8ffaf8d82a751c54872fcd52c3fcc2012b586bd83f3ecb8b0619ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf615c375a3519da20dd8ff0219f0a7ddc7e63e2c23507116d39fddbf4ff9b94417b05019baa5bf8aeecc92025e045b7087a03532e9d7f1057116d0b1868050c040b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebfe0d3eb25dfd0691ffbf21775836a1e482883b08e995d2d57fd5d19c633da610c9420d825ed7e3b320fa0a5a237e929485ad3dc1a10c5f81b0942614a74439270c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cefabbd2f32f506d8afff95782c846c2f344e9b7a979292d7ef9a396184b41755901af2a08fc6e1872f57ad10a543885682debb6ea60db4b929b17d0436e3c9eb41f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3905c30ec8d726c5268ea76718fc10a8945ccbde687b0d8ebbea1093a5db57beb811ac6d277aad223e3571552cf667c52b4311e17e378761904509a091bc296771;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5136d449c32936e23cf0f4550c8faf1a0cced1247ee94660cd7848df0259bb6dd0aaa9d28bf88d5136649b5341d0e2cda86d2462b6e24ad30d4a784a46072a4ab57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haefa56ff2dc604e185ab1bacb07018c4c99874fafbaab253973cd89f7c7ee8e6ba76797187a96f16d77ab843b27741bc51b5d6b7838414d876a731922c7a551a8293;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27f7b2b9b62b6fea7c88bd1b57c947b5a0926b97f40f19cd9a93305802985c637d4b3a9b1cc3a109d1a17f95a3680a8d4f5f84b1cba9388f23ed65e4b76abfbe1bdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f513a5fcc9145d7c5616d285b9b3c65ed6d6affbf9651045e1dd94de19be2a35a6e53cc243c7255a470f511a17b8979fb4d08414b6b819aa2e0aafb6c7bd29f0d14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7f4c421f1aaefda7be88e4b1bd8c396d125b0043a5652238b2ff4f58b54a6acc0b0d7d2dac7b2f8a4b7cff6074a0c08b9a5da9a3d9c64802944008dd6a525ee6931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h253041f6448b66cd7e1f04f89e3f187c168c48bb7d734564c36eb9a119319583b1915429607aba9c4b735951356e304d60164e0e9c72a2898acc8cf94491008edb6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b86b9a62de91ccc41c8c64b2fa7d84fb6eb8dd9060b3c9c54ef1cdd24922ad81544ee702fde685639510cc9549c306b13bdaf01823a44324c4a121a3e9d100b502f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee5a34c069d09611a545edf202c333ccba55f28d8a4a9ee3b428dce8245dad7bda42cfa5b97cc7c6106e0322f7dbbd05d1c9fd3cb77eb9687bcc5f895bba9ee84793;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h762d6169c7f39d51f8e6be651774358c1c1aa255f6b0db2092bcbd92ef0900cc2d038f96de18d579161eff4d1299b6f19db8cf5de951f0bdd59119992c4dadc8350c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67986d9074ebce122f924e03c9173fe938f7329654122e10b5fdc707dfef39ecec719936123a62223891800efb5089b56eebb58d457043d21324d38b11a73f9c9b60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h197f530766b6566321082a0b0659a999d7372ca7ade4d9142d856244483e9d5a8953ec672f836aadc0b155f559a8efccba828674138f87ad75d2ebdd7d971fd173ee3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1339c88eb99f7f69d55ef7b845117b885f24fc8522ce9e144a2bb5b7f992657a0785fd007e7a00b6a84c6cb63b4f53d1b7fe0cc7335040a7140ba795826a695af6496;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a820f4636fb9ecd40ae74f835373f7c93c3461e07919eb84d3fa59ae601b03c99d9de37715f3b6469c9b7ad72987e6d07cab02c9a6d4185c594ccc2b62da7014898;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h945ca3fb37aefc6e6d6f08f06e400b1495a36352013a7e98a900819a21aaad208343067a4858c5045601a780299981ee0c2e6f66341094aeec5e4cc2a2c5288e49d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4acaebb11f2876ba2355c860fa89d3233b45c77529830238bf877990dc9ad54a7452df2dd8639cb9c8ed9eb65c3e4186ffdd82304ef616ffc7a72e3c429e1afecdb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d71b2ed2a817e8ea862360f99fc8b95113a98efe5f8458121fad88e85b7910ea8b30308c99d94080c9e92567eae6d13de6a79aec5e7296aa4cc66db2992ce54fe3cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23b11b2dad8e574ea9c23b963725a2aa8cc43668b4d30ad3e4a65b6844d9544d3ea35b58686b7236552ce5e565df192573b6c9b96648ce88d60df36c10642e2698e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edd941c9a76cb1f4bd9c75d5eea8f2741c66b865a2ded5788d55b70d653d2aa6d8e9e0ed0ce00044f23c08aca8be8fe6b043fdeae672079ef4989fbdcb622c4e6699;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102486942986f51642bd1c9a9f5bdd63d605afef34aa7a85459f754b32da1e1331bddbfb7b905e524823561c5f23347541e26ec44ffbf664bf9ae968fabcf205d0154;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175673bf9c07f05cb20188bdc328d208464d738002333e199f31c06595b972766503f270c420430f7db72d4557361293e8fbc0e910adf448c3d1106a3435408e14ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126408418d03e81b7d7b36f034eeb4193d50b173a0bdcbafd45fb682c7b89b914fd598553cbda5a77bc334c1fc62032fdb5a6af7665b190806308cd5db090d110fe41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc89082252f8a82bc062bf7d3f6c3836d0e114adb4b40e78b6580a855c11b6064134ff4c1429f70f748c1ad94653ba4634e174968a5f90d8e0174e236a320dc3ec1a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe594ddec139fba69fa16a43040bbdcc350221c57fe8f5282d3dda3dbaa5e5fd8abe11de0e20dde578e8523cc7f52275aabc7e0160d30b1604675b265ec4b496ea9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64edfc3fc74bf5d8573839ee1497b1a7f3fd1b39fe1bb6d9e730685875501243fa7be63bddf074301e9928b7fc7c8925078749e49b259bb64304ed0aaa81522c14ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d1335e4f64b7e5d8eae443cc529e171696bd39c0bc3782bbdb641071ccd4cd1ccba8d07540441d329b92b301f8f65f45931f4f33e45f3ff8f3f39fff262dd13a5a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e69afb92243ede582cbc0b46d1c7668c88bb6f7c985b98a64ba466348810598578aece84527e88b62f495e384f0137b61c43f32cb45bee2a24621bfe1e8ed1ee722;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14af6a77c5cb3ede20616f387e700b70b5df26ca4ec7bea085d3b600cd6ddb5431d4cca91edd7f6e246289098077e50750ef44a861c2db234a39973ec17d0fdd9985b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f818230a1d00e5a5c2afc75ee93c1c13fc53c2712e52ca6167b69d68c8a7a7adc304dc855c6048659baf5b8a00174a1e8d6e555c7818f4c650bd24b9e4768123055;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0340b614456bb8817666e6e8aca7220d82a69690bd2cc8688207fadbc5ba1f402f448648034cba6e022c6919482f566969d582092b558f6fc1e96ebe89925af8ebe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h838124e265f255df2c146ff83d1e29548c5a0b04bbe6420554ae173c6269ca873876833c95ec49a461b7cf4d52bff986e8e18447291781a37675e3ffcfe8e77cad04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1567e505eb28f08a612edce4dd2ba1361d3efd7b2b8c68ae97cd729d995bb01ca8eee9cdb71bea52acd1eed82744724be77fc00eb9f5c83a6074da5057afeed12ba97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16589a8e446f462ec8324bf9c25a0c134521a67131c19a9c3dd23239603e72b53f0b17cc5b59ab36dacee009b68251cd47f33c597eecad2dc8b6f117f08a43cdae45f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94676eb5ad2b2868c8fb541dfde66213633636c6dc9c67e38ab367c49d4aece089906df35e3eada4add41707f4de971b49b900530d4e1fca6809b2b4f0d5cec18b43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ecd1ab0670113ae99d682d0e04b94073b028bacd3049fe35fbe9405aadea134eae0e85a9c7066bda9b3f7bd54aa3b50562c37e1fc0a41d6a4cb7c346109f1be57fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd638fee0bac90ad32e4645ae4f41ae73bf8927fc426098607fea4f5fc193b0960a5338b2cf71532b052745fe7b5f03b9239280e171ede5e1e637429483121658fc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3de092a685eb428252bd34df91d36c61ab8b3a7480e391d00aeb14f347e0df2046786bc00799376b503a287d3a0a719793a2a281ba3d34b6817c55b2815a576114d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161dfa3ac8f667db819c3493d389d35df8e9c99279f6af497af08a75a3d32afffe7ad3223a86f0bb21e0ec99b37ee85f8ae3c443b57129b13537f7ab72d2734f62526;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e671edf40e2fb47f5aac2c9700ee97fa8d176d57895b6101754bd6fa53ec30f0aa7c899663c680c635e9b30c26c36936d71d8477bb333fd1f13939cdfda65c46f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185b9b6c8622c1b65583232aeb3c3fcac718e98bc541d2e6248da31ec1d5e46622114e9343ba3cc13683414af54c98690c207926eca2e8ef894bdb0e86603aeafc6b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1d9bd249814f2e1ddae5be4bc0ca9cdc83d51cda39f66ca40e71bed4525a6da695cd1eb31ef507319c3e8e7395d581cd8b8c4e78508c3ccc0f9b1b8f9fa6775c00d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ef6cda032cd9d9e0b21a2077aab452c40bb7a12b512309ad04dfc6502a3f67b9f8b6386843d5f1e0097f6871dcd189c45d6b916d5e96686fe13183e41c173f76cb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126e4bc813939619c2727405ba8f8a3fcae453ce4b97e385236fb5f1183f40e70ceee107b3494bc13995f28b30ebbdcc9741d9c51a4b1e5823f3c912aa62fc158a0eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1428638a2143af16f988abc300279b300a1cad64e1e510fcda5cbf21a182f247b6654649ed740ba0cccecc027b8dbf3a6b73ab09648dc19fe285fd37ac29ede1c18d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25e03713b18f18d22dfe23fa3650a64948eefd23c6d2d8700724b2a46c7ffa08a4c704f95b40b52b2fbddce87a1155200035f379c95501df1d68a14272c6bba3b4f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138fcade4f4e52c2911eb9e7345dc109441164a4ca269a7218a75ea28df8b3114825d0b84fe56394f1510e14a24938dd82534d73f96b57c8c603f8a4e94fc23b81475;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bac2384eb418095c4a68c50630f6ef2183a03edb6ba35e45cb1cd414560b4c0c8618e8610850065ba247c1967a5f8407c8ae1718abcdce2d2151ae1dc0cbc32e3b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfadf0c76024e8c764499d00554af8f8bcf482c9e40022a743efa7bab2d4ea9bc302466955d60fbbc3f52187780d93552e85dff89324a7e96abf6267d3a4d0122486e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc7b7b4c0d389ffb3023f705e118c865be8663b4803a8e3fd1387fda5240c14ebdc45af91b14f0e41a88a071d4daffd938cccd023ef7c019cc4ac4ca35e2676527b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a5f1db9713f1c81c4d3d72895cfbe61ff1813728eeaa0bfa704cc3cb334b472eaa4159bfc9e922f34de88baef73bdb277854a55988323d0c8ecff8ff52e651ab112;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1499666ab08de538fd3f635c2cf7888d20faf848cef9e462fea4f77eff4370d12f9b82c89dfe9ad9694be502625178ae3cf0ab1cdaeb80c81f802511408ba2bacffe1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165af6d7fb07e6486bb26c54ac686e8f7027c5dbb4edde806e0a838e8bfc6177170d6faa6292f2b005a273523967ad30cc05796163296b68646a116c03a243481c076;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b60cbb43d681c56b407074c015c46fbfd7bd2e1dac815165b46ed2d958af00eb5030e0920e413ecafccd99877d360b9e1f57873261b793ec48321e830ffaa304884;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9c7d95e57a49182bc256b6b45ba47d5f96113651a8d433f230bb10332a17f002fe1f68788ca96e6aec8340104a41f8df5652e6a9637eaf391a0c11f7c2ee035a533;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d3909fba5314fe75010f5ad58e2289cc55bdb7dff10afefbaf376275f9d676899bc8be75ad69842beaf0c71443d64eb38d470a308339305693ed61a671ec92ef895;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f42aed023834c2c59cbbd3ffa50b450a0e5a91aa9ef94a552c5bcce04ada8414c4e4a09dfe564201a35a093081bb551e959c8b6cb5ccb90fb1174c52917fabeabf3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heac273c4e854d68a41a310f866cb44b535a950b01bab327994ac29c715f5d149b610ec0118b12829501ca8284a394157e821608746a4edc580099ae65fa07338fa21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1606a7011eda48fd4c452501a36bafa17217134341ac7a343ae0b44a5ae762c30c5890791c173035ad47a911e18a2f9ac480b09b6ba6d809369686e8e77c9f2e22ded;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13555a1aea7bc989d228541ebfab0be5db3121f11b8a5a3c445b69bd13c2de2ee16b07de50d7c96c7e9c5db73c1fbee569f48299bfeab97ff043ceb0eb2e650a74ff6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd98f5c8277aac40b099df5b064cace6b8ce7b5264afa7929a8baee2f4401a6e2efaf6aa0375b36a63fff738aa13b27ad3611ec2aec4de057db386c8a8c798577c053;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haac9f3cd455845c739a003e2015091b3d9b06a1511e09d169c0a59d2c597d24f6ae8e30c496762dd4c6c4005889729c52f9fb5e5dac44164364d969be8b1ccdc2ef0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6be1f820193951eeb653145fb9f7f7b8cc72fb2effe96a331a2a5db8556c536554fcf9893659b99223b154609f6675bdb3f90d2a6755ef04f62c29328ac8b8d14d23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15362beb13da88eb111a8fc270ff57c487e10fb38c56ce91963ec56176c77eb0b15bae9cb5b87254ca460d919d155e0501e8ee74fba98819a398de2bf476cdb0563b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13facb0bc80eff97c098b72fd54bd60e0ab29355382e49d20e4c0ed3f4fef092fd6c29aa08a360693a0106afd85c75596b2fe1da6758c6b412bf6fae360eaea7e46e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a1f932a605fecdb61df558252b8478ac85075ad5b48095bd3a375da1e1d0e44a3a9fac40f030f7374e2e229fead50c92b05a41843bbde97e4741992bf80d6289cce9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147416a314df59b53bf66a5dcb844fc59e1ca879d96f22ff74178badb4ea840aba76ec58ae6e907b3468eb5522491a0d50e364d6b10bea91c980a68b20efde8c18b90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fea5c8bc694534e6a41e13456a4cb3eee83ab1a461f44f0ced32e5d371cd1bcb9656f0290acf61f14931e757a7f84e7318ecd86c2c764586ee511767422a708f01b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbacc148a67ef9970cc916ea66f617048fd8aaf40b6e641bc528e51819fdfdd2be37554dbd3490175d48a4cba889ef790b1a655c0114ea86568284971af4f2b7064;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144607e315574ea42674ffab8c639a6e49730f6817f69d2c7f3331ac87baa866d34db866f150a677fa887d311a6bb721fe09331a8f37c908bebc1bb613777ebcc7568;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17016ce70bae140da0d1c89c1f4833de81a85542b227c450489e3f5b8064acc7ee78ad3f7fd271b547b51fc956538b35e27149294c4bb02c27dbb950f383e72b5f37b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143d5e0285bacc2f28196636343424b9589be01269567b83140155ea8e0887a0055a9fe4b0ccf54029ea1bd8a69a4095ec107a0e8e28bdbc44d3d99e0d0671ea5e4db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1876bc1c3a5ad3e621b9af2e32163485892cda34023cb52a48dac70f7eaa4b58617a036e07c8f89039db6c7da02953473eb837c24b31f384f3de4cfd969e8f4f90ccd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac84b8fb0130ec9a888e4027a7da8ac1a3249cf414fdc0a0d3818ec9639abe214403b2a62c187cfb4d7b869c68e53cf38a0ca0fddb4da574c2aefecb0eeadd295b71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc82a23010006eb4371a0849c7d254720200e472fc392ff1a130e8472483114fc1686aee7132825a5051ae1eec3ea9adf1f0adb8e273e1d2e93927452da85e0f7ef2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fad5757b01235d89c37a42dbd32044c9d111068143baf3d478635c697c8b651f44453c5a447757c30dbdb0fbfa00660a12c6ff65c158fe3558133a27c51f3e0b6719;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60faf65d3deb1b107b0eb373442bfea093f25f11b4bff9a0e23b413287c315a66f006b490d97b3ba1a5c759280e4c31239fb52f87a6a0f19aebe9145cbfa935e7779;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125958eef4da31ccbbd1b8e713337f636cdef0b2f290d6d5099eac991b5c0d3afc07b9b7f7aa2d76939027d56c79062705da5f04973a4da821ffe85a957d07f9fb03c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb59524d8ab5d9322d422a48919c7c5d1a9015980038af4f8da4dcaf4ffa44361347f9927c1b91098ce0ae8310457b0c15ca85c93371c8b5d2b4b4747b05ac56058;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97456c0f9610f820a945c28024f3ca222893958d29a5306f77d1d2bbdd213a63d23546fea2b6f745fed84e08feae84da407485d73a30cef7db6c4a086c521302d2b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c8d36fca42be293ed1d5e266b911eebdc5ca6046ecfeb4bf44c65910cfa4d4068253c2a3e2179dd2f618872f7e907367cb8d10399c04e114b79524e060ef77ebec80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fde67bb7caa3469a5f54d4feee94d2d91f2c7bf7824dd0e8d24d464afd8eb5c1787f30cbbbc3b08d682bab003ccff3d3ba0a1336a20f26c1c60b5f161f0c061a585;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d131e72564603789cb47b2fa13fecc812d1766d07b707b2450b0dadad3919442801373835963d1d9532a5059961fef2a472c639444ae9dc0c6d5803a248906e82422;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h271223b68dd00e0423c962d59f1af30a35e4888fe92de074e11bd1ee16a43d4b2d7282929b6d4c7a652efb436d2d137575b39a8f9d02c53a2d5ac45294ee1e7b1563;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c31bf3d9ff34ea9aec1a72b4396beffebd5506e845a18e923f58b6f9e31170653696d45d8ed771372416aafe51b85b1854e35970aab28790463f599bfcf44017324e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h786a6116a9cc888d86535228159619d6db9e3e12434dc6ce804f315c15a75a1f8b466d9241edcdb6ea32caeee55a322e7c9b20c1aa96fcf2a62c4b1d499f8167e044;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116f100128402e24e9aa049c3e2e97384b6b15da1f93ab6f65b2d4ad18b25900114c51c9988cdb458651e68f0183e1ce25b3fce2dd8b312ad261730deabcd966bbee2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16fcb6a5d96568339e213d79f6c543ac22c225832cb3c85abf9fb1c9d55d06cb3f40275cd707280ad0c7899dbc786e815e353f1349d344c339ac9af88aa1756c23e7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194b716577b71d4c26da229f22eb770c64bce879dbdf7fb38d51676e1dabfb2f744d2809b8a5022c451898ded88b6c4526d7717a8ff9950295f6675a5bd9394311244;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74abdfe976b4ccc2ed22dbdf4d0d7d0d7ee75bc747430370173329c7474ad3e7156c0c2f49fdba2e0c044f18a4c34804e2cfc38f55ef02bc8855e9277a8bb6b3207;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd76fc435aa4f8eca23476da5ed98a0855a1d76f2ac2ca597c8a8677553ccbb04f615ac2c2c1e21a5d515d849d94fc91c57292718f7d7f411a5ae309b270341cd17e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7922649e48e2892846fb87ebe967c180b46ecfc6e08401cb73dc12a872bfe4c0d9f003e4fa006dc7e178e8abb32c862b2be46c7cb41386381595313bcab1151b477;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccf94fc6c73b6e7605fa0ed0dbf62b8d7fc4297f37437b1e56f3c636f0edbb22ebafc9691f56d36f0ed6bb4099f8719836fc22b729903f4748a219d3b13fd273553e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcea93e819308acf50cd0f15e0fdc14cf5483b21575d56d45d11709bcec70a44dfdb9647d14ffff2865185fdac688ae38d11d4c682db66c0ad3ec5d6a288104a7988;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fe8cc8bee77eb2a5ff36b05271e8806aac1b3051d3f501006d4846affaa3c6b800cdd1b9f872e6ca3ea19510c0b0580523f6d3c8ba541c59c304efa93bc22900fff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16837ede18a5ff84c3537731105fd14dd6d3fde7a2772206cfe69a8b1c2ab17a3766c0b1de23fe01748a71cfc0a4a6ecac808400155cd380a67466468ba1a31f14c44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1465f6cbed6946fd96844f52719cebd88f222d6ccd9ff87b0f1183de47ee9047f59e94ffec3e3b2f5e847c19b77e0a02e0a89c4b8f0a2e02e2c7f0858b1da18eaaf8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1010a7c03e27bf6d85ffb82944f38a70ccf297176c04548288ae320bddd65635ecd3545106e508bdd8e9cea3ba415a577e0765c0a3105967457333a22ffa31397a74b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162319cc9e585c538e3f58faf4b16098e848f52f02c75d328c1ba54781a15087b88cd1d64f8183753e0947a32749e40d3cf46e4d2a88aeda75b653ac9c2f6298d032c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1634061e7bcc517c777cdb2f6ce2783362fd2ea1d1593e175bb106c87804d60d8d3a7e28a5e8553fa30ec818c529863b2a8d54e4650d60b70983606e19fa9135e90a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38da57bb1e155f3d92bfa45293bbff6e404a5bd0a9d333c114df1b374bb0a5c29ddae862f6bb3693e864096fb49d33ddbaa22cd89d359cee4130f23c63865c59b70d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d1d6ba32f7485dfe04d2fa18c3d411cb12c06b07875070710f01ed2a5b07461b024abaaf41bd5f8dedfc6d634bb67cf9c6e4e5e858169b43fee245a022e926a34fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11363f90060a8666d5aa8fb5a7a036ea0fa49437dee6389519b4dbfd66adee775ef4cc00eae539f07f92b78bb1ae2ab44c294a1defe749a3549e3f36c19d68df8d65d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9096165ba603aff2c5dcabfcc696281ad3beb7b167064bae88a958fbc37f9e9538d4b2503df82fd97ec756aa553156d758eb930e7a1efbfa2410e8c32fd22b1593ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf817cb1a17509ea443431f2aeeed055d1d6de3b0915be8b374dd6a50e4754ada42ce909b1142967920baf8fe070bf23f35da5ec350318da8e20daaeeb151cb0d67c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6519178f6023f3089dbbc3375a630b7061de12512c5ad4f020351405d21fd31aeec500f9294e7f835701423da49cd8ab6736d98e47510316057ece9c82a5e1b4dd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b0c496b969bcd80bf640dcc3df448b598e49350814dfe6542f221d12c962328b38d2a8f4a68e0b11f9c47d436710747bde88711fb8140f5362ae6c28629f570195;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he86f7640b0339b1f1f712bbad9c726720cd32f18f0e61cd50b040b3cd452d1e592830ac088760e68a37d7a06a2c015f9c472099699ba56d4ecf1750ebc533d534044;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174600b6ca9e8aa38c327d19f35a29389c0e99444db852549b9cc5cc751acc9ad59c712bca5b00ca0d4622142e8cb5a72205e8048e1c3527cd5129f3d48d84d5b86cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a7ae2970fde4d6e813d53af1bfe558620044c0a34bde50e68a477b871f3870c2d59c8bcb2a13c3a8c1b289da8a0e12dfab358c425515ae316060103d2e3acf2e3a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8545feb3e949b38a9e37a836d75d5501d839dc7767587fa8993f0ba630982cb9408e8a81d019e9b25acebb1c0e2e6687fd813da1afeb343b89f15ef348e60270615e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151263e637ab36dae0bb271eeef42623cd4bcf2fe3dfcf46ea44ff6c5f3bac9a6434e8aa7a55e0ce3473f05d77542c0fcf31d0dacf78261c4fe97e788a578dc39a407;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166444fa9ebfcbae739b5d938d75900641fa778bccbd41fc1cda0d041e75d83af930dcd9700e3b9296465c0bc2559bdc3b3c779bee88bfe3c01450cd12c54e56ff64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df432644c824d073ac424a6c6600dfb18590c91b697d97c8193277276e7491d6796b27f5a685c499ff4003168491f6c9116c77399e5de1ddf92f83728a508513e1d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97eed83dd18743472b1e65c118d3e479d05531509bb506955a887ebf29583feb849fa3f0d4defd8bcb300c651506abebf1dbb5551d33523ad2cb59848b16bc3334df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115eed5394642b915999d5fb4a7cc6d8ee9787721cccf7206837ae0a2f416210a69ab42b497c38ab6887e3a861c28c7ef2a2e4b47ba87d4ed157640923bb59fea1aae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b26426c02ad9ca11e22b173b51cfd2cced879e36c8da967167f664962c1d2d9ce8175bb8c26b35668470f55bf9d499fb41c879e48ccb307a34476e2be509d2920a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c3dbdf4cd190c2202ff212f07c566f2ae3a41ad5208b92d1c72ab80456d520dfa8b9a4d1f32570655e3e61c6976a30e0868564b639f667675dabd354ea3c3c2776b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had740db8ed75649d397ed14092d62303621328fa7a3e8a09b868c331d4d66b9138518b42c645df1ef386f1ca14e66f1daf045216f7f92b70e870fa7219a221cdad08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5f13db92ab7cb8eed6c203836af23be27d8a07cbb865814cc12d249a500145ddd4be564bf17790fb0092b065ee6154e34100bd6dbb60b3060cf91e417dd0fe27a82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18037672ff20680d60683ed2bd9af12a389ad5433e7535cff5a348c43ba1135487895c777297fde79701c02ff934a3b19bf0350ed08889c701a73e7ba73cf099c4278;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16cd7d24e38af6b58ba816903c4c5e490aa9f778da3f3d134e8e557dc8a4d174a767bca329b9f9d35f1285685489486d9123de6d4b05de688f0f553307766158dc178;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7499c093370054dd9ffdaa3e1d9b0dbe0512be9e0db2d214639f08a3cebc284a61abb10a2050fc459258fbafe653302dd35746146ac4b0beebb6e63bc850371ac0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102a817ca6ba033956cf3959cb9122d7972b8d43406c277fd8370ba0a52c5ca3c54e7be6c09c44bc26e7867453df79e7271c17a7b6e7acc605bcbc749a14781a52228;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152a89185a47bdeb10ef029aaadb52a122b2cadb31f2044fc60f8ac100d5b8a01caa0ea6f6836bc7e3aecc0bbd225f426d2a9e9dc275559ad9ec4ddb1154020d04828;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1599afa8031f877979688d09a1e3cbfbb91e6987bd87962c2df21adf2f80b3fdc5d3c6ce5ae71cbbefe0ea11d289bfbc9c4141953f0cdea72c49d7d9c01bd41e47558;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18176c43517a58351cda4671ee87fe50ead20b383c29d49f37103a8df43b638d385c52c9f35a4e8dfeb4494aac1644f1aaf27e2f99a8e7035b987a6bd8eeb3f980ae8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb2dda9f44917a2498db341d178a9107501dea42328445d226ef978ff41b04a7e439f7b3c925b1acdba28b95130476f4c09033d7635b02ec98425c3d83e012589614;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135f77ade09e735981305dad32c7493fcdb8d246ed2fe9956737f25d4759c060e08b6b24e9b97747bf387638ee375a59c14451b2c7076dbb769a06790b061dba4867b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c384dc3be927afbb92a2d207524ac170ee1821a687e82e76a556325f648133075893d88baa2df3aed2d4ccef79bda684569335e2369174ef6a2a9e2f053e0d26635;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187536b7c54802a164a9f69a1a7f536ec81ec1139b2bde8a8ee7a142d5eb60ef3d6c7c36346ae32f5827ffbd92cf84539907c39b28fb9d6e367158c449f71a4de998e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4cf4242c99fa06ba8e8bc7c18882ea2af3fe5f5e2dea5df5ce4e7d11740a45dc36f9c4258787bd02f04664fb981c4e1e0beccb72b1cbb3cb3f73c287e414ea510897;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa0ccc944b5f423d5898398a07709b6d8dd3330e84f087be994ef9b6cb258505153afc0ae818de1283bea792eb679f74b0a09d254fb8b3cacd559fb5f87393393068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3b2e87e9fceb404fac38aa8f607fc0b52ec1a8e1678252067945ca4e630f439bfb792e3d32a6d1b105a6a1d4c89b558a25e00a3afa709df5afe19f51d00e1a068f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1010447059b1d0681f818dc8accd3ab16279bc0c1c719d2fb7d33d2d54b1f3cc4898896850eeb00f822ab8e17c0261b8abb4755ac930aaa0bb1e4b2253a19d39c0b00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ed61f4786b071dbad9c3e907c46b319e87492fd193e5428427772dde7a63cfd4a8eec76e34083ad09f5ba13eb3c983d2c7b55d9d26315d2726696e7b351af561bd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dc0e55b251f9481f1897245605d7c0cd834409bce6459c0c69dd829969b1fc3feb73e40a145f233bbe219272345fd1cd2b072ac5350e52a7c1704acd90ac656e205;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h63d5a10d2f7f035c4ecbfab331fe012bc3e062e779b1ecb5edb63840c3ad7ee0a9158e5a6c2441776f83029a17bb2d6ded2084775b645accddb3c2bd91cfa3ad4c88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121cddb78093758b30ee9f2b3b3e02071377005006dbeb6bed92afa71eb16cd368fd13cd136edca991c43943453a38a31d26845d63d9f4b6a89e509261fad27051b6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc4afb47273cb5097fc7a85d1c60e096d52a938703c1b125aee64b1cb8d968cd7f28005bc6c2356383f758b2e4c7c29d52a5f2e82499847eca3515fb4050b9d51b42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9345f586565d4e5f21128826043a5f20d329407303fe576a805fe213e31af51a788e34e6c6290566e487cf77232c240883013de4fa947ebe6cad54bce3e9fbe25e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f162d7174424eecc20b574c62f5c3d812577bda774e319f2ae87e0d6e85a15265b9bb81c41fae996ad9d6d6b547e865a8747ed7d7d6eadaf73e6ecfae99cba9cc2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cdc6c8f1e25328d688d2b9679703f6d0fe8448004b34c0beed3d24e199edc865cc01208fb73634c5c58f426b1d8501f1aca8ad81f829d1986d039ce7e0d20ae0e1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h63abc8b88d6fd967890f7942a85b53e20b8034cdd8783fda84c7b8974277e7bdc9394255bbce9916e5ef7ba3a754dff91403b3b26b663e73c37ab15021e245e1816c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he44dc3d5f00b4b065ce37e50bea5d172a15107af2a18bba010c8fdcbbbafeaaeb67f87665c1c7551790c29bc4f929867d3e43f4855b5c7b2d2527be682be3135c63c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h959fd0695e0e2778d257bfe7bb41c76daac9e88cdf7bddf7309ad225225fc86fb2148dcc4f5dfabb7273e9b3529cb8c610a49043ae55bd5f5a6a0a65bae171a4287;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2379d28709496390b7f45b28bcb6c1544f92cf8479bcfa3b7ad19e0aeb752dccef0b752f65a8d996f126ff6ec9b02b284c58f648172a8cdda1a9864451c7c9d1e749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8b64d073a07ed6e685e56030db2c1377e2956a34ec3415cadad427abc26f20880016041047121cb926b78ecc3a643c4ce8d457a4e67357a2193abecc40de0676b5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4e35f93512a06fcf5f8a99cbdc44889969ead8e846d675a7b8ba290784679efe6ff5288cf9a026e96731bb6a4a36dabb5db36d179050dcd5cde7a873c65f52ce967;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc026ba93375c0bca4d5891d2c74c4192b3f51f5e32c72b6125b5278f9377138ab020d99178e57e0b672d1e0948120b3d240eded91c8e3fada4f84b3842524705d119;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb30f4d1049e8578e98445df6507c738355055ad9d99062bf7690f8a82d98589df41325de84f835dc71905b90ee7dda8466b746c144f027090810fdb910d3136dea02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79ea2257b1e5ad01bfe9f2f837f57ef9f3f733cdb120b2be9d77b0c0fecb63b9ccb026812e887b4bd6644393ac5c6b7a24c69704b033030bc57d5a1b26f39428a6dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h346a118dcbab40efb48c63e1a5cbbf2825f5badfd87dbcaebdb47569fa93aa4fa62bae5b51584530599a698a87623b01b09f0a4fe1020cf592900457f2f51d82497b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198c8bd999696f0f46b4d17107b2eb0ce6f85453fbb51a05e4bd2e9e35b1ea923a826ed8f6b3694f157339d83d794ad31597b24111f17d8064c4df61224667fdeb12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8b31423402aeeba671718a6a24b07a93d07f33595c35d8b4ffc56084ef53ab8bdbebc0c1ed5be7d71078859f3f69560c987e6ed6ac62d2b567895172255e8ac50bca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b25a665201073fb4dbbc63cb580c1693559bdcbd786922af87dd9fcf978a63920a251b36962db2793bba6c46aad903133587d644edd275be3c64886b50e5e327c73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h622c7a77fe3cc87f23353c3732755afa47ca2a6e597e0cdce614cb31eedea4a917d894b76f0d29aebfe7a65913dc543335bb2fe0a4b9ccca45afcd10865266788b33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4bae13f3e2f9a2244c7b6dec5fc882611755ba85110548030c5927fdcf3740ea0be8eddaffae9b91500d4bc6d6ee5bd765244cbf4a423cd36321ec9f9108beb02b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19cfc7442e42d28ca2e795db8eba55cc3a1faa1fa1c58fc43d30098e0442a81b27770099a694021ee342a374f332ceb2049e97389f31dd48f74d6f1b210cac3db5794;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffc9b30cb2de47c82041e22c28838da2cc228f106309bba38e1e337f741b203bff611c1c639c707d055dbab86848fde8a66e841d90513d72869a9caa2f06551f3b36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf26a868537df0f3ede2eb04af40ade1d85b636149bd6f79c87d5aa1a080637836e39ad78735021a6c865cea48ec2348418b153d98ed263ebaecefc600702d4962aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad96dbfaf7213e8a6698c8f9e4a417ac925524d0487df967fc39cf7a763c4e12e78ddfe1180390306e812eadb5236646ea9c62ec2d348bf73cee5a0503aae677595;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55b16bb2cc1ca49fb607afde5c43586f0d7bae8e70fcac51d307aceab9bde2446916f4f0e69996d0e292b0e83427bd30428e478df8f4bc0491d2e81e022dea109dab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haafa1ca31331bd11b8c45a47b2c7b4cfa96569dd569b72282e6570f9e8ad85a8d0a36da70e5e882ea68fa4cfdbbe30a9f932c7f1175948388ea3edaa4a4de9171ead;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbb7a86bbd4b156c4dfc53b38b06c550073a12c8f2105535159b994a4640063f102c47fd658ea8f8016ce01474e0e94f9978fd3a6adeb92c0c390dccf41a6e9233da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f847caa9578cca2180012c38fdbd09f84fb75c1685b167a0b639c3a246c83b4d8edcfed502e993a6826244e099aa4308b0b763aa256127a82935c08378ec1d2a5b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5c64b247e8a3e793bd3784f93a3778b54985be84b13a42dae588f5edc42c7b138db63e2618e874c2dca22bd6153da58c7c28b16ef9f280769829f8b77a723647326;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd19904660beeb641b503b1a5dfeb65b810a8e78391b9a52b6785ca2e1d0ff65fdfc3b2c05f69cd13352208cfae5826addc94f7df22c835bd4163b2e4cd42e5d4cc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab23e13cc7c8f371d95cad854b5d0b39fb4174556ea3316835f4fbd94d35570555694c5f0c95345f8fb1cfdac70cacf5af3cf8be701a3d2c29ccedd02b79f7e8c7a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ce3cd63392dc0ba04a11d8531c8dfec006f519f4dc0d1111a5378e38ca30b2b4ad40d46d934fe84217ca236c108985213ec6587da021bed101d4fcc79cb8f57c498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he72188593ce49d0acc8f2ae3fe126fe0a3b23b77cdc8a9d4b1292893eaaa8f8f4767c8da3e22465c2ad860e8b29b4ad2d15802516cf7ed4c35a7e53acf5f4833fcb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff9f8b133f6d29c0fbecaccf74dc5214efacfff4f844ada32066690fca41ce2c654d3bdd3c44efc136a79394c1f014d5be81e5ef08fa74b99dcb88dfceb70d97eba1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123edd14f8967bb3cb5051014fb1558b919c0c171f992c5dae03c9315f2ff3264f9652419f97c93009c421af5afde817998ef4873fc57c892688fd0835a378a55f780;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc089e49c7deb915efbeca33e7018fa6a180459603c22789b83beacc9f7c731825c875fa250d4cee9ce8a178b9a32a264cbea7047dea83f7f226e7da4a5daaa1d8cb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175a30825129e6357897b1b2659f4fb6f2bdf35eb5985ca8cd7c72205e3e13a8b49308377a13e5f57fba1125714eaa9c3d986d12f46a00ddd03b45f967f32a7625f07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c6384d6f6f4d43ecb7cbb0eb7d26d9490f19b322024dbe3092a9abb9ac761d5b3db5bf30c228502d099f14a78983e3f8f299d67fad652e7a2c1e1072bd95f9ce301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f65a5adbcfc3fc59a43c936627171d37022b9f2f97af4e260f3fbba2bb1c2f80a7544f2db9b8b4086d19aa0bfee7db124ebad3851c3d5797cffe6ee9798c81652eb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h288b31b7b198411a39bc3dfdd0a481c80f671ecd3fec219e696d3406d2acdc5b3a1cba316e0027f0654019e169e7f8719b9e4d404976cb89c97eeac4b3140afc0237;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152ea1bf651deb467e85a68329a97e32f75a7e16cc09714048b14d4d58657674673a0a68a94ad82d537b3777147f8bbca08b2aa8999443380af74ad9aa5a13b0b11f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31bd57338f586e23da242f79d202cfb30f0077656d17de1a26b872b2f4120458ac6718511a53d8d15530cc4f093096c0605e553d8e63896602e94e3cc7970f4a6648;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127a934ffb45499d7a62a9cbc69c6eb38bbd8cfbb0801674bdfb626573e25e6dfc4a09c84406245a288cc9ca237ee454d581f797d5c2e1bf2e26135010f4c0ee6d699;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138a8aa5a78a39825fa1a9ca5ab73ff99d0661b4eca5aeba902c1607d11f15bda68bcdbc74cc4de7f43a267b037fe480ee0e9d1b5c6cae88958dbbc13dd7b7f283291;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d2549b28dd994279f3bdb342983a8ca05a9f83ba05b51441039f3e65e9ecc22a8e3340ca9eed2e217a00a44a49f475d61e21db177026fd984da9d9db41b10d911e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180dbdb5c06a9e20bbfda15a1cd5dfbaa9afedff42d77ed9970ba3fcfd1af6d54b1fd2c73f2d4401d61dfcc4f614720d158f60b0cfa4b42725662bb7d8ec4ea77a242;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fbe8188072cdcb1dd4207cab07f4e23331f7f2c106b514cdb6d406cceddfdc54c3067c8f86b8eb91b01ee364b4b1f41c49b5a8cd4b8b2198601b16318dd35bf5776;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187c56a0ea6f41ae7c878e48a94647835fc31ccc74fdf0700b315b4c5fa13460c4ab85311e843ff93509d95f5556e53aee3d68764d8f23f0fd2455f6d60bffa9a2eb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27a3884ea900dd6a096107c60a7980f207ff2fc410e2b8a255c9f6caa84e6058e48956b6a151fbef8809ec248181a2de8859ace100491337f1afb2dd605585c4a241;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a56f20504e67e566c532781c2f4564bee8caf08bc72c29c06c06c24c7fe1f6390bb91c20f37c83d4a5ec9f69773bc7e9ae8b0f8b9a7c6deebcc549b893c3c957a31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150b6079e469ebf0a17327a0a150b90de8f6be47522b003facbc4868be10af8c61cbdc446167a9ce1fdf8aa87ab3cc6a2c14ef709656d669ce9f524a2ddc46207d4ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he84d9a7c964bb7a44dde1393c20e8fb47065d3f1a1ff03c42f296503f8822da46ec9888c78f7702b454066bdc1d5c6523fbf661688e66084bf008ba182c4295092bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f898bda467e4b599de850eaa56bdd38a99a5698388e5367311a7cc1810894f3922d37cc7f3d0fedd7814631131d0120b4ea79578132a9851210be3f8c9064245b56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a9b5161bcb0f7ad64413448fe7d18ac16bd3d16a8aad139d09fe3714f41514c37bdd3afdb6b06fdd86a1884ca3187a167a784292272f5aec219b75d5944786f901a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f1382bd1b5c22bc6ce491112ed62bd8626a5bac4d8adf4d5be34e5edfc2310f2ed21324a72bf2ea2a1a5a245eea8b92d6ab24a036d0aad5dbd0c3e8abce57effbcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98e9c376adfdcec107459fa73c6e61a8b392646ece3505d16593b21244c390511db6650064b934675fee6583907e3c8169ba21f3b59c34ee450c785a8a10510dcb9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c821e39e96276bd596653986ee57872d9d4304cc7a5843fd694fc01a2f2b6105fd2d78e2e69999a617ac837acff63176fcdc1d375543514232ab665899e2cc27ea61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4092780591e31f0c94c52577e6fa27c172289cdc8c254bdfa0337947695b82fb7892baabe38bc407acea91de7e06bb56322944e8a73d5d5d10c583e54fdf933f56f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7320d3b4b1f4d71d177aa86b9ec3c74588d80a4356b5dfeb02ea2cc825687a0248ef9ccb3bac412c6d38fd04947dcf41dd0da0cea87e76a9831a109553de9b4f9c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h619b3c559e6127167956c1b432996035701dbe380dc5ee543ffe6c125b2dc67d5c8c5080243e8afc86411cc0f30dc7e7373baaccf1f5d9505b34e28e99305a2424eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2edba76d181dace19a04dcc992cf9b97a6817e00c10b3ca9e75f265b7cdc171f559d65c62a2089dd6745be059df2995c5b9ddd8a80ef8e26ffa5c0d52c46898a9327;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b356e3ac20131df44c7a3bd90cb12e853e58455b9893a0801eddab9aff579ab5e6c7b15dec52b5ef447bde88b778ca53add0a1ba12dfed8de2cdcc7cb21cb531a78c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f850ff0a8f4320955f88e55500a2eef391f2688fc8313abeb792fe5aaaa23b3483619350aab19565f8c7e9fb1341344fcd28940db4c492a47830572abcd55ce9fe23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190a7eeb9b1d9be8c6b78fd25417e7f45baaaa56b391932bc9e618c9f75738d36cf7f5dfb90ee98e168901b78bfaf15ab7a7fc9fa108afe2b8d3a5167ff92ad6cf395;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1793ccc1d7df89c88d3619a9286f1143f0747e36a33782a637c318cc6fc02b3bb3ed95a2f45f66bdfd764a8ba10837530fe28b7832719e791ec0d78682c0b322c6594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193ed16db2b47463a706888da03f7ec4b9b09820e64950aa689a3c25e19663b07b7677439a1f69dd4cf818e0a2506fa43a77881187fed0aaf3476c2c7a1ef65a0f955;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79eb895ad80a3299508d8717a73a5f03d4709c3b86ecdbe2a0797fb0584be6bf1ffd438b6b13d9522a148c2150a98e2e6b4445fbbaa7736a1f74d415c28e05ef47f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha872bc6dbaf174e4456877e3753bce083b48dc8593dcddac7b4065a040b0909ec93a70091cb76a2fd4b151719e9c6fd8c6a866931f6f17f446543c714dc6357fe4e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18747b65039fc9ef09735793da3c3a1cad8f67cdeae0a97e23e14b86818cec59630bb1110cbc3b97c6dd588a276c39aa7b3934bcbf109152ee1f851249f7d8d93f0d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14079d2ef7647dee8160964d15753da924af5682a3c24d61dca0eb9dac1872a1a1f5fad15f71a644798522c4a5ed164c4c39ff1b90f04f49bd9a44c0da9f733f1a46f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb934a65847c9521f709dc08f7aab63919bd01a1032091664aef81b554b3a9d6c9b995c06aab7502b8e5de39687fcfed9662174ce2a6cac5f348a1bb80c41567f3dc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ecb0ea9e571abee0d1a1d4e46b6b486fab4e5dc54a7f8ce20df276c2dce630e96fef17637d96428d655a88b17d34be5be74f3028462b440558b72b1e3d1cfb67c365;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d54f1003012369434fbba1ac8f088b09a048cfa0daa7e5da42214a54ad3c8eebf7b88feb75b8f6bbbf2063c8557394db6214b57d31983827bb40a245c5520f88af81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1384fde29163310a18a8f55739ff91a129eb1d1179bb42af167389e1489a2c39583fecbf0fd4b81a36c8f342b1d3e635c9c71be53765c58dab1d13122780d276ac9ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb9481d4bbe8d9dc9f2e82ca35c12ae2c141ed940e736ab5c82490d7522e9848f7449e91875a7ac3ae6eae425726f5acbbb386f06bb754b714d7627764f0401f0570;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9f6d63e3b03758ef0b79a33b2d719e49f4e7036d4a61716ce1a62cf733419d56906726add7c4e827fabe627579951734bc5c66c1467f8609db0429859e43a4e876;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e11115ee117c15680dc08f973d768e4cf0816d476ced0f63f33bce29b0aa4aa530e0b3dbe962a25278bef2136cd1651bc33c235d34e9a35df030dd189943aac1cc9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ca7b156d25ba471a9fdd7b4e6eb1ca889740bccbc5b7fac879debd59dc2c98fe42b1ed5e0b5b96149c67445b491f1da633598191b39e16a906cf146866038a6db09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab935313f585cd0e0ab62b7bf4bc62417cca08f6517616659cfe53fca51011b6a722de8ab69f0a1c2c42a17a5c0414959365fa3dce91bbd52f9ec4e5d195bbdc8ec0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2041994f135814d9acab23cf751b81080b15eec0d72f515f2cd0efbc7f987b0d4b7a691de3803fc7e880fa0ba33f5e9a300ab20b5f996b8005f04d883fa01744752c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bd9c2b671299e57c85ac93a1645827401b6aae62577996eb1a9377d71abb9a8ec184156dc35265ee66389de62a71752ed1758cba7f944282702d96dc3868c3ab7af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff18d793c7eaf9645f9c9c1b2327e3d4221ee749cf1662b45392e3e026b37807b137ae84c388d5285034dd0d818d6c58162424fc55ceb86a50693d553bb582ba711c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b280218da4b2be00d2ac038f800ce7a22c139f20d3d01dd8a053e1fd2a7424c4ea5df2ba81f8e78de8336f8ac8c2a1d05323f55abd0f148d8b3157160a1d75223e87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d35784c3d35169ab9a042907156b52bf89ce3f6764b09e32477604536b528b42aba60fc0e70087a54fcf080a0b93a4438a2440606726230a22f2083641189514d5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc2d5ee021f710dce708a65dd41dc52bf79953495f9d3bd436827c3ce6ecdda8351c3a1a3d3d1ac8cbb9fadfe89d962b60513bf289f146ecccea4d3292589923e21c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34a49a0eee0f4242a9cdd493ee9506e9dd7afab2faf0ca6a5f8008970fe4511077a30b418e48807448323788afcae34e491eb5f46c88b985b1da0b8583517697ef08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e5311e11b1417d1f1b74ee901aff4db6f98d63c92ff78004f60b5b13d2da889584e8d8e2f5721a3b9a36c9e7108cfc8f7b912e944982ac7a171204e397d0d3de8c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9aaaf6230c75b0d3caae6f3379f92ea006b828fe7bc3a69acc94a82b3f52728226efdede56ab546466a97aa4680bf5fbd6e26150a5972d4bb52aabcdc0a32ebf61c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5cdc850bfa6b422fe3e098b13a654514dac20a198041392d3b20a5b40fd333ec085eeee7fb646aa8578915cf2b557de86c4c1faebdf4b340c5a8e69a7d6dbc6472f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73d80003c26ad7a31825285e8d490de539dbe099f58b637f67a812123350fee96f40d9cfcc03705b5ac6c27f9cfd0815db6f9ee35cf3d09c342f4cc61df0806f3eae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfd41693e9878f98722306a1fc9a79fc2da8df9e9df6a202d12b62fc422651242e2de7d3764581fafbae4c8bb8e7146ecb3f09b42c61706462adde735a2253f6e82b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb65b20accefa19757590fe3c697c6c0cf56903508b53723b22f7b158941db142b88c3ab84c01cd860237669017422921280e0155727945ad504159f2e708493018d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h939603a72bb3fa60e2afe669930ce8a5b5d6fe8a659bd33b825e14930e946a443c7fb29c2b198b0a31481a2526f1edf5d6bd3cda1b175c3f34f979b9e167d346751d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107fc906d9500f9e5c8e8086601435a501ea36aa3ed2b1e4a5c174bf4d89350e08fdb3790fb4b5663761778b6cc32b69469b572250949671d8bbd2256802b0aaf2b62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45a29a90198697268996bcbcde489818d24b83877d72e188b763f80d17452e581851f503cb51a4b9e79a7ec3ecd6b88725b35d9e16d2d905192a0bba1bd00870ebad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb1591f1f4ec4d27c8281126fb823771c70058b64b8e60cf0c1d7fb7e9f6c117f61cc15668f93a211e6fbfc4f21830b1bc3b2d39459b0f1791f531e270a3a8cc57b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb96bdbf72cb71175545160e67666061d19c74e29b32f8123c2457d06ee99aa3a7740b3710f899295e248a5ed3288a7169fc0b400a9974d4428d9aca51dad330bd9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b667ef133e3abbfdd6316deb263c403561dd13df70617efed3f6fdd76179fb935d93353d7000eadf4feb162752230ab0a1ed2374e52185817c0897f10e0cec6c9705;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb71643e206dc25cbf4d3ecf5d797db17112d8c1541ed62ded3c760d0382cde45574dd61c3694f4c5c47aa65ac80bd078cd5a28d8160b6215548d923870ed376a9566;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96a9a94392f0d561bf03fd3811f2e436373351044374681d6ef5a95b8f37693c97ac7069c7b9d41843798782e6097c92b007e3ea1149bb3b00751e59cd1bd767f228;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f92ae0bf517bd1f82e26a31b03fceb9c0d8e245a4b719f4c7173ef61269b3a345353c9c2ca1192ba3c4f32663809b7dce59b6b0f86b9c1072b332406387e8319b099;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128c30ebc49c467b55a2719e6e681733884b413c9b4a5ecbb15843db408c97d2071fcb403519e59c3ca29fb6b8e7356027350827d07cd6d8fcd6ceacf61cdbd13f082;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f77ca4bdc0a2fd7bcf758123654aa99b84f46f52f4a6919eb706887861dab6c227b857dd950d07a10f46f53ac208ab39e1a4b325245336a0de4a40fb4d5c3bf0bb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3ae39386a37e29380a101fc403d9097ad41c5fbcd53480d5d785d17286b9fe679ebc20c2e5216679755ad833d7dedec22bdfba858b4f358dc32c95e4047fc8d5696;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f308fa077caa11fdb0d4f3fd3e7a9ef6c1ca1474cee7ebefd2c6e949496cd3d004768d00217e5e43c3394d48b99b365c2b9331a744b83b4bfb257327010e58d26e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1371fd4372f6c4d878a9125711b6df3e053b60ece70164c9d13fb70a1eb7158306daf5c214ccb55a1c92fefb4b78fe4c5d78a01c242e429d456524287d93b5fa0e1eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefaad1e4b99dbee3348d02dbc650f699722aaa73e7310edcae097e88020ea59bbc7344e6585432ac243a5cb8b0ebc5cbd5e9b859f2e393a57c01c223000a7377c9e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d830cb76ca13dee62b2798b6bf55741a5134a85847bc6618b56c05fb8c985f79fbb433e95d66861b72f03fa9141e49019ca0b66490f5e8b48d56d114bbd4d5d079dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b0642da5dd19fa30510bf337e03f26ae83bb6ba024e46fb682bdcb7ef4ceace671d9d7678dfd908ba395fb01c6f882877cd23ad988efa3d229e144e84937dbcdc59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d51dd888a391f1957de1c490be60d2913ab9038851465f3df567226bf2b7985b904da244fa0f07250298fa574e3fff6b5d9ea0f6c4684bdf08921a6aeffea9af14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1578b905267a3b446a934ada7833f596a4da0ac9c37999c6727629a89a48734d205056eb0de8ae02b3f8e7b9ca6076d2ac3f9c615dc5d2bde7e7e40076e77b1248bdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64f8a9db8715f40f5757db8bd697086654c86b9459eb689b7f711e88816bd990390b782255a445d05b26294a01b5128ef26578e2a81d00887a5ba5cf39fc76149161;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cee554ba787e344cd81c2e4756636273535ecb5ac2e00dad3509bfccc2643731b2dea1f8dd930db9428262ca22171bf47d09289375b83983b72dd9c100eb3f85fc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h662ff3a1ee3fca7575e5bb22fd7b475465b4e3b88a298a3be1b3a4ff574e2e468cf443c569321940f606b7a0a145a7fd8fbb6d399f8412fd9fb794dd3277a2f87878;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79fa10cdd78a84952249d521145c7308c4e17d9ddb2e2f5531b368f12508e0d8eca286b47a063662df1fbcd8bc2a824136810b9c78be25171f14a8d93f1af5313244;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eacb72944ea502e5c8cd6e96214a248cccb186bf9eb4796178095299c8684887a5ab39e3688a7be3c3b326426de7638e8d47db3294f7fb41d1e53fd84d4d2c76c7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104ebcd08bcc894bdb2747e79de995f6587e7e4938d348a82bdb8c2542db1f6726d7643cca4f6058994fb350223c94d33c13885d0ec2a5d1699266a953c1841feb3e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116830e539aca8880b47d7ad3e8679e222c9f4e1e6ab420161b5ac801ae13b2aa4e7d26f9d612cdbda62a43e85771de10f71e493e386cde3c86eb36b7993041f13625;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a1a95bbab6d085524e638050582249c3abd8cd70334fbbdd04695e66fd1a7e898fd68901b4360ffaf6c4d601a57ee60cb2471e8cf1313e71d8f512293c3e5d5f28d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9db4a77b42bc12125e845eb7e2bd7452e8c893737499954a1e1b5251fa90dc93c42fd3f2278bebb834557a5ea7eb897a5ebc0d38c432f2f87f2ceb40b796aa1b5b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ad3f2223fcf68b09abd771f6074d30974a203cea4f849ee060552fe31fbbb5ba614b1f1dc669cb5c9015442ddcc89ed97edabd1e64585ad6281a3ac9c9789d3fcb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfc855f34801356418302e25d8d9330d6f046f55540aa2d26bb2419c3b609bac2ae15305be1065bdd6345c330edcc62d6cdd702b729888178d4d6ca7f71f0bdd7768;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a790ceb94240859f02daf19391f23ce3235963e9a40e4c49e3667dacc3ea7945ba7fdd9d1a51c94da1b054784f1340ee4b2df55a6d00d0f00c29fd080a086a9c0d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136e4155031f3238f8c3bfecef5ab1f008631f00648236ae106ff20d7b234eab710bd4350c678677e385f08b796b08f852b25bd4a2f605a041c1cb6bf3bedbc3f1320;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26942960ece1e4366dadadf24de3470c0417ba258e88b9de0a2cc87ac6615ba16c66a3ea1470e484e4b7d61f4e33a0930ef50f9ef6153909265213440a6c7f0e24d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28c7bab5d1258f1e1716ce0e1acb34a3c36bf911e4f5972c4106ca08bb7435ca75e218e75b7c04f0b1f4037b6931cde4dcd4e75ef4298584403ea098907091284fb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53a9cf98983c655c29ca0390e47ef6daaf590c1bbd5772d95edf9a995f4a061945a0dc6c8076112a77374294b8a8b862b9f8003db9a42cb08bf43ae3644637a8f40f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bf5a9cd178a80d6ffc19c743034e65c8fb32a8c0d0ca50e199a13a722e397d4538cfe00510f50bc0c2f59d4772b5cd15f94085670634f0c061124229aeaf6d8edf3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1292598012b76a6d7c1bb59a37ee29bfad49bf57e3dd1365df905c61ad52e6cedcc469cc732201ee7c57f08d7ff4e3c62a0681646861fecf75c1b3a19d371919954e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cfdb3330857cedb9c8eba91c4a567cb43fc264990c2ee841c82be7c8b3386554386b745e5f1ec7904c8b490e7aaabde1cf92c479af96dd484ac793f0323d998f462;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d10461c0e2e77ba03a02cb6d3c91e055ac482d24a675e3fcd7d830fc305e4a52dbf6a4e4000d5408c86eb04f6fd010aee625f976f583467c670a2acb377a1b423b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136f724bbd38df0e81bf9a70e738c8b1cdb3bcb9963038ebe48887bc73f59716c513363aedda08c66259937eade304accf0fe5c5852fedd6efb2409eec4e92383a2cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dcc2a66a83282be29cd3cd28fbe69be371cc03590bea7ab3e86aeca7859236c470d4e6019795d055e8ebd947c6d5e6335a6da7d05d2ad3076a4bc88e24e8f931013;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d5be13c7efe3d0c84936f22edd4cf17586736a38e546a616b3fa43946179e9262e265501ee9944098c7eea1163514337a84fe991adf913b17c4a76042c7dca9834;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b929b5c3bbaece11cba9209957aca96f49d75eea3d2c07bdcd62d15a9b3c25b803d518dc0c56eab360d57f87ab5f509976460344e57211750862fb2b10510365e7f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59194c361ea2f7dca885a7eac5fd150d1c39ee11a55534a338dc431024060f80d83110d93e0a2804703575cf7df60b695bd3fdf77e28fae41644ec9ddd8f7877ae27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b46bc5d5ebe4b2135e21e906d3dcd46e6e50b9dabc3a1f6f63fc02cedd33ba2b90c660076b477ac8389aa386975a35b012141edf66b2bfbcd245af1ddb43b2985442;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h687eb15ae06dd1649f602b0501ef1615254e77c810de36d6a625016de17cc5de29364b550a1d9272ac681c77a84ec587a5ac4115ec4007c8c958c70b0080fb40ce3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b0d62d9fcf070b5dbd97011906f911218e43aaa5a6c7e05af92de46de3f9be4f25df038d7c45dc641375dac876bfb580325b0047bc5e411ebc86da1ae3f7b4de45d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1345a3922a8c82df895268cbba32440e31ca69c347887b8d0b877ece9967008472fd772b336fdd50cb4c5a41d5c20c6bad953df05f5b40cd07ebe015ce6d22011718f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ff5ed23e53dc8c2a2408c2192abaea99bf0192a72c4d9c8c09777e7b3cab96a7421065f5b59463580942308c9d66888e66c5530757084bde7a7e88c28539d947dcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184aeab0ad07966f2f391b20ff2c1ab0abaac2402bcb7b1816cc449e70059af2cbe644c935dcc81a0966192829f1c4517616df2a55f1c2f1209aa988fce927ae31a4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1746a039c6b98c1c150ae185bc6d7076634d88ee70f7a476b0f3d62236953341b35925629396e20afd3c215e2f914a3d7eb916f6771f14c5fba5dc8059c13a808fe7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce551687f3d298d9dd7ffeb19eedbae590f84ccafeee7474f8761d84235057fe7f45c7a17e5bf1e34326b6e6ee7da302b0c326d66340ddca64cb94af26d8dc7cce2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc77ba3ce452d24331b62f018f79d9d0b431562ea90a60440e0b2083781e4ba9fc1e912bf81d32eef3cda8b651eca31e0968a4b0279686d7f43a9e48bb9608821d1d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171251c8b55a5987a81a3abd4cb33b208657925bb333df58add04ba3f7746e177e94eefaa95fe1cd0654456126f20b822e2b367f360f28aab7d8b78219ed405e517f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2a945c409ff9a4898cb6d077fd0af4a4ebadafc92263dd6fca83857c62658697dc34222816e4a7983b807659c68d371c8ad5e21fe3580f6f24ee4dc4a27b544b3eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1712f4d37d36b63087dd744d0b93a97b0dfc8571a5e2e97123a6f8fd3f900c21d60ee6482ba839b9cac4a10941a46c7d41cbeaf6a88707c947b2bd0253cb71e830c31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a32dc4f2ea9159a5b0bf9ac9bb1a817898c804bd96e05f03d3640ef370cff2d70276ee19d96211e59496b11017a6e511fc2316ee1e33903d7107defeeeae613b0baf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b850281881e7a12355cea72b296279207275d8d39d76510b5ed58264da5d5f3fb5282bcc6faa766247c59d553eecbfb7a6e992c4d277a441fa89395b3cca843e480;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189ae85a367bf130578ae99f2d4df9c6b3c81937894d77affb8325ccb0e1d17fbacca4d96e51e567404ad5abefebf330b34e210fbc211fd7258886455603195da79ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3212bba367fc4b9d88a8160c761916836773d65718841dd42e3a46140d08cdbf53523eb88edb4f1de397f0b41ae1cee057c441ea74159e694e86c14fd227271b177;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1995985467e37aff13352f4ecc12ba003e8cd4a34d7ca521da5afa98785690fd11969c5a8317ad8716c2d20bc25703d9f135fea04c74b4bbcfac92ac482cce8981741;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15571f38cfcbb311b4d3db6fec8c292a325311fb2edb4eb1218d9417e9a73b620763b00bd8ec498033bc77cbcc9b646c3185bdf9f0467143f3c835fc631659debb48b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fb5bfe34c620db8acd8914df2950e3e32157b980926b0fce81e91d9613e5fc2b8be3d86c15873b1920d942d88fa9bde89c8ee8dc5a1e120a92c86e541e9e1e7099f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e6400b2f5aa1239eb8fde8dc312b1f5b099eb7f044f9a62266d79819fb668208c7038775586bc64398c4df9473fc7e1bd5e07c77639dd8ceccadd4f7e5bdf954ed8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ed76a85e6f05545d5494ae62eab28bac563b7d322ffd26c4d6bb6767f98ba583d2fdc6a3f48a215c596950a1b54d45d2290e33589197dcbaa8831c0374578cc5450;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h903ab78ea2e569fa5c2d5ff04a0aa0f177847850150f6b20b82647a6db8fb185d344c80b76da1b3c6cf567a5ebfa914390d7b9418be4c4458b5c67f82ea09a6b8a3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee4880fa9e10d0ef2a5494a0b640be13491a9729fe0109365ceb94661a0731716408b383015509529ea30d9c65379d14943977056edea5285f33ac56c7103ca4350f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37a0130de22e35fc7ef6657b276029b8ca903ebce9ae7e3ac1e0bfd8a98bf51836145333af667633e6fe946fb08f64d0c438c4f35f5847f77651c8cf1ed71e3e3e8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e3e3ce0eec050e1e6a2ed41b1db8f1c7d8771601d867df1c3bf8cb5cf9f77f9d437e31a2d3f54301ec33d21ac862bd6c0d80c52a97e787037f52a92356dc79c3190;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3209fd119f6b102473fcaa0aee3e1fe0ecd76b417a5c1d9c46bd958d7b882546b8b7f8aa2aefb42154faa3f00c7c7834a2bb7231bca416eb5f329c4a455db77c2ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f5c8f20c96aeee2e3d138a847cbf1c6bfee37a841c14a5419751863d3c424c74421e209695493a3d00ede9a9cbf6a8686949c0be1ee4bda6a0e311817e15f9cd106;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa9be7832da8d4f616cad169558cb8a1f295e2403336cdedf0d3d39b37c0c13c7b2d28437be4f4aab55f20ed2ece0ca702a1fe01e23ebb05be801a0113ae1f4c2c61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf08fc5b543bad1c0a25f549c617cc3464aecaba05242d4532ee7fd3bb0417b64276c084d18ac0e65c4a48033adb427d8fcbc351e54325a9d43c6dfacdf92fb8a785;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a70d3afe9bc481581f7439c01c6b8d1eccf44c655b6ae3e88e24c37bd8c421e2a51944c08397da41eaca676b03fe9d8aded7a70ac95cbaab395379d7b91146c9389;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189ea410fc75363d12241705f59a65f24df50188b0e9a4204b70cb6ea3b68071e8e72da94deac22313251fbe325f5676f6f3a4fa0482b03fabca4c3a68b6bd59a6a27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8330261878a2e523e9914b8dd5d2fa1c7ff187a9960ad6b6a3c1b67724c8f5c1c270842bd3e230deca532519a6dd94894b7eeee8102783589f08693cfbb015a1d709;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4483a9fc780a639016345e782ccb022547fc44344c203a6725b0d2197e74c6ef65b5192659302b4a9f5345858ca25365b4ecb552f6426f21070177896647ed0de476;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177e30679b82d30e37c0e6a2c63aec75d4c85c01985c938e6c9163455ec2f5fd2a2a9c83ded8f21258abf875eab2a81f1f3a218fc81a2ce32211047acaf5c8b7a6336;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ce0751eed8031dadf38c3a28432485ae9aec5845ed45b1990c8722d779e63c40f4774b7acdbf39fde5887537b784249fd7f4ccbfb4588f2f2473b7e1ff41109d9b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10549e9d89d25d655f35e4972acad21ffad3dea6bc2cd57c2120a10743e56831c79baf0c80b784c24bc032905508b6cace4dd0d0eb19602a20c09be6b10201c1eb1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f7153681cb870077a0e44a239bb5e52a46d4612f46f07ee7acf7ea81c2322c35a48e24b61965aba48f9d55bb40eaa52efd815ac93b4a56ecbb12c4d70c447c1a33a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de5be731c01fb7e961bfc0bce23b33da8745893ee799a771b305287bc7b34164af1a86099159f2e7bf83e99923bd291186fa34b3542e15b38c4156dddeafbaab55c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he128ac4318df408224c477601fedfdeb1d9a75dc6332b72ca7b4caf5cc6dfadbbb3378db252ad2dd4fd242054e1eef7bc5b75f31ee66b7291cff0a62300feecfd493;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a46585d509cc75d9f3353bb6ffab22c2a6bb8a47718bde1e04390eefd13805eae60067b03e70a96742afc5aa4747d2cbb5c2fb17088f219b3bdc4fd04114688225b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8331c7f545a299dc49626f8e0c68eaf77d914de8816e741ed87ef8aa4abafbb17c30ab106a0d88fba15ff3649f324e4dc81fa96d91f7649321eb9d01b19cd0831011;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2789fcbee7553022416372d7d4ebce5fe2e62be13678f606ff9921f61129d5fd254064dfc761f08a39db4fc832b46cb02795adaf720c07eb52245219c39f6f95aef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h278bd51a58cbe050a70774a38f15b9b62a45fd76381c361fee28264769f17ffd79970307c11ef5e2526f07308620475af0e225c9f3bc257fc64a56650eed8eb37b08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc28e80dce924b8349848bf064d2f96f8248f8517f94440cc6636bb05570eea30656ea10e01ea2203ff67d1b3a11f13378d5890e17984780a472e9e30de7462a63159;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af5f8d37d9e1189357b6bbca50408a1ead6560882e66ae7c23e05a44b8dc25b7790e1c706a5f6a968abd6ac7a66f6749e6d2401d064d5b1b65f8e923bf28065897fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c9b3559cbea2f8a15e630fc0df7dc1c12705e956a6b66a1af18744de845c615dd7d3888f9300bcc07ba6f242ad38b4fb8629f043d8c9a1b16f130223cebbef26fd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfe796a953ec240c8d359e0f7f0b560b79d6078c2f05f98151ed8d8b0c18dcf7ef4f7cfbc9a01b2a5db0788dc262838acc6399671bca151d677d5c12ef0be69a17ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4ba55daa263d004c70a79e07c6edb4db390409dbd73a144678b2eb5fd34f518297697b24e16ffe75b3df66d89c642c8cbb3c68b3e9db8ba817848859772d91660ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142445bc11858f1633334fc6ae995f4c8e7ea7ddc8e3d98e60f7e795860ffaa5ff81186e107491f48174e7b943596940df105248a9232dcde906d87241711155d9140;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fb1b4fecf538499386883dc34fa038258fe3874dc12a88449f52ada6991d5e04b8292ce797072215cce3ccebf065109c673faf1f6d762f318c0bd03f35e2b3ae343;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dfc0a1965bad2f26c92bb6be8ed019c362aefedfa7e244ac6e036d1a71ea60ea5f164c37710c2f0676f88bd5f18942c5cd14d18e2a5673e3e6c881a2f288ec0f112;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168bb5abddb1e6bda605ae44fdcc653a37d797401369a5f05426ce50ff2cec30e4db2de5b49b13f144406a34bee046c022893c33c2753df4ab656ea4509fa102928e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4d615715044624661c677e6a697d1f2ffcaaa42e21376c283c698acc3523306bf83ba0a8d7d0c5c76de198df277eab79a3d21980fa5138126a21efb4b83b989c77c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heac80e626e9198fcdf66aac2dc85515b124210307e44cdc0cd232621904e4a2f04dd5bead389846b4ccc4c21b619c16a35ad49105e2acd661b8f5b145bb8b66477a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9e89d7aa66c992cafdf39d13920bb8bbcd4265e318544585987eed249ebd2d2d9c9bbeec7a2e335677bed588cda1731ef0c0bccf00ef9017320d44960a114b3ac8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c23427ade2dfdca74dd62acfb55410ac6a03f0daf536d8887412858859e60bb337b865f18c11413db0e90ebcf500b28749d7e880eef5d119700b22a2edc8826a2f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h836430450a4bcd00e939dea9575baf564545bbc9b51dae82c70e42dc7948202f3d0022302c81f9cc4e5d7a0511011069ec48af37e492b4bd420e5eb37a5affcc647d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9a20dbd916d86343d63006e26d2d61655613d09a2852ccae951537c09b1fe308f7332aaa6ab6a480c367098d0d3b49a92d2b447eeeea7ecbc4eaedc6848e78c6c47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e698e752009d8e5528aa084e4799ecf7fc3da4590a7efe712a5eae9278537c2494daf4fd47fc7c412b2678195e7d6a836f3106c172ef638efdf2edcc6dac5732e5e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc07b39b504a3fbac371b8932485465efa7f29f63e6127151373f8d528775948aea6cb92066d798cb63a0d135085720d22e9df2ba37dd64615d01a0236b39c948959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5384de36c613cd9572dbee183c312deffd8fabbe016f50b4e124ed4754cfcff06fe1a143ecf452247e4befbcb19ac1452a6afbc7bf6a4dff6a220053a91ae3b417c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfaf3cbf703198b1718ee4e9630b83cdabb612125c67e929652d7bd35c457e726816c5857f141c305c320a9158d1b78a5eb3cb2de32bfe411167c92f5c4b13f4f1138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd6fe267b0ab12e7cdc6e6fa1a4d292307f3b09b86f4eb49ddb6e278097d68b423e29c5cbe94888eb226e1a8f5fabac5173c7143418476b192d130d3a4e65bb627f3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd81f6b7adace3f7a3fed04d341a2a90cfd454ba6e6d52b78a3110e02f570853ff7978d1a6d86489dbb5140cf78060390fe6e53a7f094c1ccfb75a135def3ba249e11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94dae4498f925f26e48a750e3a28195c0e0405a1d4f2ac6c9de41fe07c7b1188b560a8f69024681f36d0d28cd0bc0a9c240f8ef564796c7454bf557ab3d892a0b543;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2062f3cd7e6c4e704f10a0540d6ea16867bb636d1317a7c0a51ca109df6b93d922cd01200007b356da3e20029dbf91f17b522bd486b23235cbfa9ccf93187428206;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c7df8296dce8df0021b1c9c8c37d1e3b6f4c954ee494e17a11feaeb38ac983082f45f97e8b1a50b552817e77275c3db7069a6e19b5fafe143bedd4fe65ee1188189;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3795421741abc504a86f4be2ff2ff1973ff56257cac07c493880b4243231c8ff472a3fd406c51c1f00fe9a09a5b4b4e51057fb273a48040f54ec0515b41151ac5561;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171ff0759ba4925cb264801d43babe2d0aac3aeed7267e9fdcffc9de25fba367bf0e3a222c25c602207293355d085f8ed2fd779bb28aafdc7c2dbbe144e77f2d030d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70690ece46272380b8b6276a00c2193b12b1831825f6c86b41c908e4d97092a3a4d44d9e10b40f0f3e42f854dc93b3ae034ffc9a4532ad1467544bcf0343d4635d01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2369b12cd521c9fae345f568cfb4141779c59ef11d9a3800f0da96f95134ac6eb494813eda4a905196c2f85a21caeea9bdaf7ed572a2485524af349aebb97514b68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d7c729d9518f7ea625cff863bc4dd1d65fa59ecb66842ce60fb13b29fc8cd556912f462adfd0bf2571bc764bc2203d3c85de70d2bc28c4325bf0325465b952d19a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4533aa38d01f7e51736d6408264548ecf2fd9d82ad524355329276960ea3fe6d2411737d388908d9a1ecaa6d341f6778b70c37ff3fd7b1706a1adabc13ffa6f4743;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c09000b2f029fdf1e5e34256fab7b4391b783d0432bb511aa731ec6025a7c3638821d9becfedb2b19a50dcdd1ba97366c2659d90453a5f7f97cdf23923fd91c463c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141c0fe4641c25fe873625efbf574b7a354b115f45d585d79b6168b2eb17dfe3cda35bff3432fa42818bea97daacda088c6c1049e368d748d30bee3160820a8e0ad6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103215d9cd82192114bd5a1324aa2a3bd16767735753b85cc1a73618bddac4ee2731656b155e8cf65eaeb40a2ff5965890a04aa60f498d55d989a3d73a4414f1e2d4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadadc69310dfeb38344d1412f76e22684b93797d03cb40a474758fc92900defba33acd710c79f9efc1520321ea20b8f6b6cc929f0634817ff3c09545f431d0ea89ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10132a41aa989ac555bff4e4cab5fb45288f6e0ce206998dce4e0384c2d09d2d65c21fc48e38f89269fc0f7fb4b8b67482fde2b8cad71ec4364bed69ae6f0b9694b58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h859b15445f7fffdf024fdb06f95a3b6b2223725c675b23f95556fb3dc4bd314a3ea2380aeda149e4d750724561344e528e10ddd58a68594fb39bb29d16367bbf422f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19989afd6e2291a4e6a175b1bd37f6690e57c9b0d672a46b3c65e1cb03db8bf8cec2cfeac3e1fe599ae9a81a353e0c432a2299b1f12d70f83beb3c34a3882ad772123;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c6a0f514db0308ee2bd606e6436aa83e6c4b0e66f3c953528fd65a861031a1c33c7e4193178f25fe1084bcb158920e71e818d64eb904bd0baab7ebb4af77431819b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89bf45b8f3e57a13ce2b38ba73b97aee0dfae25df6143c1d5b9428a3d3fb23930753358d623f3e8d578319c3023eb57871ee62930af4c19e4a8890efb6a7694a2446;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53871f333c94f3709a27c80ffd6e08e33b32330171fcbdd57c42d2d0de72ba3b237d88615af376965ed77fff0a0777d4076951c1c4838ef6372684e0793374b6e08e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fb96bc2d375ebd9043a0249b35a9dd49b5b0e13a2980f73bec7fdce70fef9d8d5ab6fea45e07f938d432a9c35e66e35414c57cdd436506baaac9c5c14380f3a2d6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heacd26b63ca04cb63b2a600af5005d15be229d820833865719e6eb17c01248e2fa5b91ae5e76aac7e1ce81ff0d0e0461e8e1b5e6b300506ad1cb7df9ba3fd4cb7b69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67bbb387df103b66654fa3bbb9a55966173d7a753b4eb26ce338ee031a085404fe98bfc19466ced9fd221290ea7fd4318605266b36df3210390322a440b67371f9a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0a901cbf75d3e013a93a0628ba4ddc1ce3c9eebaf0ee360f971d3c272b67cdc58ca3fb1b0034bb38eaf7f7311ff491ae4673d8ac7a056cec958d35808df54469a9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17efbfe499d3e373ab4f52664af98b9f97537c2dda30da71e962e19658bf826475db3567b795ded6a292fdfe4d8fbaba8987df4cd8c8380b3c1e37b97330703554fbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b79f14540b5e5c720010a66c0b71e6d99054ca6d73b466dc0c94f858bdfec9eb64fa933de366cd6f8686483de59be0127de9e44cda5724daf0d20e8069e4919bcfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26ca33f6e1db086631182b5f5a4f8ecf333f56a326b936bddc2059fa9504da723f73dd1b493fb8be70f4486d12ff20c6634d56ec47ee737f5d5d06334fcd04629cb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b5cbac1e40be44bd1fbb3b6e0607dce70efff6e6fde5d6450d40c1d58d1b5966c6c163d7d603758b60fb7c8a02389c04330409585cff40ae78d37bb39c89c3878b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11be10834fc56f66b961f820512d07c5abc0e7c4230739415c1098d88bb3f6c3cf39996fd0fa0b57a5b456c8e6fa81b69a76dfe81347b0f230da2180e59a7bf303d96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ae9a0574c2ee3a8084da2c724b878b8b4d1c9f08be8d9a0a86d7f348aeaac75ed474f5dc871dc46f24619800eb9ba71dbf0505a6b6962a8ab88d41211892e1befa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180632c8143bc0471367ddf85780219d9d8c235f6df501f385c03ecb4054bfa143b92091686ff08a029bde87c384a12c3efe89c1519e3784c51129027542b19b7cc25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e36abde1c2dc79953fa21e0273499e7a88f871a62d751f7e389df8ffa9b00809e8a0f717053c4f31277a5c9d9a504f5e81c8582d77dd44e045e41bdd666006a2c87c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h860ea3c82d0f23571ed86649b6bec381bc4df53ceed70d5e5d09497b6aaf612806710c0e3aa13af06562c722ceef72dec65dfe89ca510f466982b0b5b6ab49ccc9cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fcc4044dd34e9798f65136398bf70a601eb157fc48f52cf895063bd33f96edab8df771456da06a9ed08580c3f4116f0b671ddb0c223a56ecc7ca717fd569ea569f48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f861e4dec80701a7102826e797048c93cbe28c5c08c7ae547ce649ec3902c24c62a7ebd82c61ed87822a8b3098339153e7856825e9ae139e38d232bf94800a4b320;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fd2bd31a8e04a86cc1c1b76c6a051d45e08eed07b02e8ac6d5984e79151fb429f70938fb921cfb93bc2a5162af772269eab813a75c9e3a448df7bec25fafdabcce8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafb19ccecaf6f7e130639705e3c74ae55730eb0afcd88e65ad0d970ff433082084e9617adf9be2e271eaa68491a5285bcd7cc8735b6842523e1de0fefbded8b76f6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h450a9924c210e4cc7ee206a62f98b3704b5484d5857d2d979a72b123a38f503f7fd3cecbaa48a2a69ea9e0d1c59611c9e89925ebcbf4bbfa32183aae19f7b7822e09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4900f6caa7b901b0a8acb2f40a1dce3a9298734bf88fd9a9a982f77afa47d300872243d8f26eccec1530015bd8e002b56ff8f8db26f774dc574b883c77720904f0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfaf73b2e77e0b6169322de4b4dbe1b3ffe7b26158e7d58c4d6310b404efda4933f068583c568124d0579dadc79a2535467b777c264aad645a02379f6075ba109f419;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47ad87e745276871e3dd3061f4e1d64cb1b7c640f3dae2b8749af069975971cffb9e63cd093cf8edd4e00dad2fea8130d34f27df09522782b5b4ee74e7e27671d002;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h768642062c82cdb2feba82eb3bf256155a8f52ba27de4ce4454ecf8a6504b51d8aec3f05298071d78fd1e4ae9af600d8891d46825bb70242fc77c1c5f85e41c90546;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h227bee8d4dc1d7ee9872b1916f317f6da17540bbcafbb337ce45729213a74eff0d496052c704a0afb3ba6a7b5bb2f83b2071f8ea96ffff48e8a48a6f0b143a295039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5a934dd6a696707322167f96108ba91ef89d84860552762a0a51482973b9fca4b45a6f3731bd7c328d2cec63401e7a36cb9a03678203312bb61ed1bd79a84f055f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180b05ee6c3b62766bda7b426402c74cc1b41fd530602dfa02782627852fef3b9a39e70ea36a730251999c94f3116949171310e5ce83c50a94663154f85270881e78a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f860e14b055dee873cb87791ead9a1933450cfde11a0556c5a3eaf91f4db55c0b402de353cae0ce8ff0f85473c444d767b8cb0c01885aebe120367e858f71a833dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13edfc19df39a15b4feea6992cbea267e7424ef571043b780fc6cb5c17feeafef4717d32155690487f3394b1a85314dfb03352c2ca17a3b31bf1d1c52191d72d39fa2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f81951edf7749398e471fb44a15e24c30907b053399dc7acfede758a6866f9e1bb5f82c664d2c2178cf7a8b97e36b8e0e3e145ff20caf3bb9920ec4f3c4b2b762673;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cedd02c784b0bafd4a592e8d1074148ce5173ac47a76c12ba173ac14b782b3865a620d01b83a423a09cda75b8da04a40de9b9f41418aa2cfab34b1165e68f212799;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h750b98c2e3c6f202af4aae3e19560be9c8add7876e23379b883c602be4d9d2b07446681869d43f2fe026531a299406dc2e20620ffc0ef5882581b2ec9087d5cc4255;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18234ffe899967308c416fc96161cf72e793ab4c57c85e040a08d147c07b66fde1d45d531c7fe7f797a1b1630d0ffe4ade5b2075a60f8166a7676f29877e9914453ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dfc879088ccb255ec1d2a8d9b44e963bca44eb5809b65cf35dc949b5bedfccc68a7414b86227d8a1b92eb6ba2db3797d2347b740ec1513296e1cd90d32cd0153193;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4bc652931c4e9c42df1c1912cf4fdafaa5e48c9c466250bf85ac0920acda7c8cc431717595be94f473b4593cbed3c737cdda27891df368369060c3c21598e7d95bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24c5de7c2d3dc9bd613e6442a4a12c79b5fdae8eb40d12dfc4e6542ecdfaffd5af3814cecf90b15e03d968060c31e18f5439b0c8e226253836e0de2b4c3196dccbb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ea41b2ae5842bf3bf0652ce90e2d10ed0157afe0f02e1eb81c6ca78b07ab1478ee958e0e736cd5292bcdb4badfcfaef7f0fb878a74cf91d9646c456f859ef2bd88e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb29584f187ec6ccc66cce7db0609d0b2d3b2068573efbc03b8f5e2a3ef43f4b9c83d6ae8f23401322bf58bdecac94f6121dc880925a2869817083267bc0d82841efe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15811be8e2f70ee855e6ddde645f554a48b4f62db6be4bd725f5373f5f440744a81c745e5c701e171e7eb4ac1656b3c6c3b16dbf031d851c9846493b35c30e72a3d36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e12f7fbf9de3b3e8a033fa83ee960b6385bd348086eb82b8ce3c70cd649e644d93e0d090ded86c36995fb573ae1506bfb4c62d9919bf08d4e16f1c5e5e594975b5ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6eff644f25e0c39ce830247739e97720876dbf941a5063ad54ed24590fe421651f9c3734d0ce425de198f81c01c2df1ac5888988c1dea54b87d141d4bf58291a7039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1790ac28715a5f4589cff1e8206311f44bd7c001bf002dca053a33e5cbbfafa13d9858f083fa2b976a0378f00d66f15b91cc07ef51b394d9bb805dba5857177f84fe5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1d62c0584372ac76edc33d4b9ee129eecef0c1dd43744715c8a41cfd595f3a3ea3f5fd6940a3e01f97260216deae413edda78d8f46368431c426d364c9e1e7e796e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h626d7a19c4b73a4ed5d558d932e56839aefdf38e8d6cf83e4ae274045308939bf189edc1534c5463d0487328cf760f8453a34786663d57338219d0405bf167b1cf97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b48faf895e5be343972015c7dfd90a3afb7994896981c77ed2e9aad65f947bbefb652b2a3b4868ad73d6198ec5892809211d803a0c22d5642c692d525603d71efab5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba2b07971cacb55b3b1fdf9292d586422475302a7220e853df8417804d20fb3eab3f570ba3d005a33279f4829f965bd669e9673a47c7a9d0492c4e259c87155e3d82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bc6cdd5b172db8c6065519921753bd120327d246c082d8d96f4b9a9c90767470c003a4d549c14a380df24995f686b6bc7a856b09f49ec6cb3eebc1baccc69d6f21d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106ed0ebde8210c024f001a1c659dfe65694500b3f94259e6822db1ae1c44ea991594a1d2b8689be92bf50621206b24d8645a1a9ef25f31803dc728fd991d0ffa731;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3c1b2a62189dabbcc6237c139b431c5ccca8350f57fbbc93b5641ac59458bb822cd48d497b1f6ce69ed9c6ba139787f86063a0f285a0c3ca11d0e69b38e25bb215f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ef2213bc3b95c6c2733c8db6eca8a6a01e6e08ff1d068e176e98cf881cc2d4ff61532c709b63907f7c67f07c9338ddcbc267449effa4c6510a620880f2c3aed5ca4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73d87d369ab7e8dd8ea2c502ca3cbb724f72f8ed4f62adb4698f2ac59575dfd3abf843423e04715467d4d1895baeb79b981fc01ea28513ce800d0ca2acf4bc0c2d01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1946b6b1074ac9db53dbf03653cf381036185f34aa83928c98e3dce2a7154a9362bf6e5fb056fbdc3be8c9f227edd4f4e2b7fc063baaa861458a74bd3e8cd91407c94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d2e75839648eaf071e373944073be71f59141484ebbeb85689781f80a1cdd0c373be387bc3fc331afbe48170073d32a008f9c0ba78aed9dcf90d5ded7628b2c475e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51b907a711e4772b26f65ac42250aa48e71c6c66af6d354635792c927e0e5ac04988baeb01b5ea5d7a5eb70d583536a861a044d16c80aa9104ecc10f8a7e3701cb2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ab979ce3e9b40b31d04d2d9149c279bac92d2c8d50cac5ab999b3ec135c748f11dcccdc1af80bbcc67b1df3ffff2482c0ae5c638063f584e3dfb69613ae5d877132;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b6240d1f4e2cc8ec6d083a273b6fe086de42291563021e3564d0dbaf754dd52fa803d64694fb0dc5426db28c9ad2eac19fd20881bd7132d768f9396a9c9f2b01618;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7b6a648c5f49dff2b1ac9bdbc4505334810aa37388f37185b3d343ab6f84de15b9705fcd17a42544d9972a70a72c5b76c2080eda326b2743b611bc2a502a6276caf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66119b92567beee685b3fff4a1847d069067964717a39d85d81fd27a11d99d1655556a23650a16f2c9573c8d5e8cf4011bcec709879309cfcab1d106013304208040;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d7b11aca85411383ca09b4bb17a8806b172c76a26e2c3b803e6dc55e2a6d37b9a6b4dbc0ea2db6d46ca01dac5cbdcd1b876bd3050f21a1920e0292c4bf9250d5742;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68393365d4b058583a01e4b38b544f92d3caf5a4e7ace67113e36bf8ca9ece54bef1a9c77ed28fd79b65806310ad8b380d1b062df3852b4b3ff78e26ebc751961095;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b66b1cb289355e9865e88ca133fc6c27c4acf4421651bb84dc5563d62ccf4535f19f1f16ad2fac14984156ec120831dc989a45b4a5f5a0db6bedd946c36a31d696e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1b173ca2d7ccfce5245ce18e91e9d8447fc29e3512c167d57fb5449aa99d55e520aefeaac59fcb42fc845270a5ef0d22635827289a9bc7589bc03b925c6bc374a9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab71c8addc6aabbb2a137a253c2aabba86f7488b9dd99e1c6cc86edd3da81287e07001d6b707d71553dd7b6cfecdb26f590a0a13b1e2d76d72a53a00075feee30540;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16454faa3172dc04034f8559c297f377602ab8d23e40dc31285d5f3279cf5110078b14e13117e7e7e6e8e0608c4ebf12c5c78516a2d21d5fd9d751413f379ae12aaae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164da962de651c654c553d5ea56e01e0c7632679b14a4551d01f644e9f19fccf13b2af610bad1846e5d316bc710dc8f7562c5108d04f8d318d4cc2566d717150e271;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe0c4ae00f5e24e7e08e3d37ee65cde09023eea668b216a43e0a0bfbebfd1a25453db090271be44a0937408274a7ccc8c2d074c70796ad8db024d9a6292d4d4d8e0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9ea2b84a00f2d4b897220a4ec6ff731d612c8630b8741f22c093cd50ba705eb4aeeafd0f3a70fc3f3723ef7b4c767715cb1a9db4048f2cb6c165bfc2884ae9c0068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42978a76e7e73e9fe4d149c01de4e18b2b7ae23790c2edb28ee30c029ead59300d15e07688df7402d252a65ea8933dc041d19aba1ed99e277640aefb3419e17eca1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f42099408138841213f154566651021965ef6a3c20ac487967fcd3cd20067543b9da49cdbe72b32b1cc5f5dc09356bdd40548283ec3bec5a01fa24301d7879d093fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c5ab7afa7c2007c206c06b7184a760fa37fa32e6e925eb57fad7631c433d44e5b76a172bf5c8fbe2eb92e8fe927e3bdcb0e91763055c7a94f1f6270a673073fa73f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9499b814c1fccb90c0e3d3b8a03adb6a05ccbef99499c291c3c2d4dd9c4843987bbbc40b2ad17977798f3913575c19e58dd4c0605909e7c8aac95bccfac605ecae74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf56fcf250992e267d2711508ecaca358d499162a0578914b05283816b9af11f32a61125a14dd4d12f43d9bef7f395e341825a7f7b036b03b466b7393dfdf780708ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65b1522293cfdcb474447d1cea4d09e3d35ee5888e9e5b9e8250761c2a49172b484f4a8f934d4eea4702275f5b0fe60ad398a214ce99a24149d8f884290e3e7e52f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10aa68a6e8267a02e0a1bcdf43063974593e1a4ce9c3e7cc0136bbdb9be54cb0bf1588d4a58b6193dd82629aa39dca39ba8ced7728a782208a75c48e5f445d0e2f520;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbed799d15966a99e507034a65557c2e2a4716425720257bdde3695f98976824b2bc2e8c3ace667a5c928b81c12d49b636559c57de2514d13d74e408aed9655724d29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h754b773c93870b515fc461cbd7e443c852a139af56ec3378591ee353eb37803a78c29a74e45d666a8fd9ed6782e1b4a9dd519f3363a47be7ab1ea961acf382c3d792;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1507d188fd787493220c2793f69779b48aac4f9cfef5d4d9c45228ef2852e6b25e00595e62fc46cc5e67f932cdb37795a6d23e53f825e9f623c6bde445f71a69fc861;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c3306e0beeb8cdda6cbdfa6f261e4ba4d82184bb05a1ceb2375a1406f5b6a3c70d0767f86a5b09f6bf365d5e3bc3e55a49b30ecd139226e84de74770d78e0b67667;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c99098d74faf7d3f267330461ec54425fbb19d9b47d6d4b9e911a11540914f47760f775f1ad4a192eafc8e0ded73fde25f8dc9393959e464a618b9b435cf629af06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6d9cc3bb9cf555e75f1ebe56a2936650efc1f193a38f0ba032a17062eb4d64bf715406344a4d1caec5973fddf60eae4e2fda452fb682f3322af1cbd7d7b7cc0cb91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5f3adf8eb7acad4268972e80d594655b0d5b0df6551881afca84ee854c80ad6dd3ac261ed1c7bf4efaba749b624b133f522981d8be5530263f9b4fc85b6242625e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67d7b1b33d16f33a3a0a15ec13d1170008286a8ed2d020bad869ab47ab56a4fa836c858a9f9d7f5be6ead32b8b28080f4f2efd8bb6e9c617e5633da32c6687895fa5;
        #1
        $finish();
    end
endmodule
