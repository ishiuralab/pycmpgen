module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [19:0] src21;
    reg [18:0] src22;
    reg [17:0] src23;
    reg [16:0] src24;
    reg [15:0] src25;
    reg [14:0] src26;
    reg [13:0] src27;
    reg [12:0] src28;
    reg [11:0] src29;
    reg [10:0] src30;
    reg [9:0] src31;
    reg [8:0] src32;
    reg [7:0] src33;
    reg [6:0] src34;
    reg [5:0] src35;
    reg [4:0] src36;
    reg [3:0] src37;
    reg [2:0] src38;
    reg [1:0] src39;
    reg [0:0] src40;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [41:0] srcsum;
    wire [41:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3])<<37) + ((src38[0] + src38[1] + src38[2])<<38) + ((src39[0] + src39[1])<<39) + ((src40[0])<<40);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h840a13f4419bc056293f946151704dbeb4ca54cc84d35a2bd648ad52fc865e44bef1d62def5303e5d314e5a88e62bff0569d866c7d406c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2dfe7573efa3da85f71d966e9c36b82358bd6ad358586a19b806a5d746880db485a513eb3762ba0d4dab9ad22d3c964b96e4163ab6479;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h952c049c0e2916ed02d2f18cf6490c8fbb8d0f5af4d1c6716f6c3bea280dedfa9ab0764a43cf18628fcba9fd87e37170ef07edc01d28fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf1a3b9a679f4bb8e866e5840750bc646111076f5e5a8153519fc01e530933a3ec62304b4990acdb2d85d92168e5102be09bfe3a11830b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55085f2e2ed7b101aaa2345a7ae27e836109020b5a7c5bdf9f0d58c64540586da8b854c58bc5acc07f723f3496ae6d3bc20867222fe335;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197c8e017d58dcd4dd54090131c21254278e2ecc5e14cfe6af4221bb1424bb4d5a4fc15600c13d6b0e7f82fb06a52c02274d09ac0693b23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c3df62b3d16f0b7a72511d7c905fe39ef33c02562aeb5b001d52eb7ad36de6f250ede613f2d5ba656d18aae9abca1620b0d673c7b9604;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1926651eff1ee94af5f00bbc9482d8ac58ea1806da0770962bf1bfc1a1690254dc3146fbeb895844a43562a36e2f8e793388dd0ad8b541e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb41bad07b0772a777e0d830db42303837b52dae8fd189842f7fe4322c59e0359b30f0e3dc94c4d88643c80e79839055eda7c0f79cbdac5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110c0984fb78d46b0b920dbea0c36c1cc8041ced32f783e921f5146ee1c62e04fabc5a4a9a3972739413bee78f3529d492fad1100c42a37;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1568d7e1cf85e48d69c26ff99159751cd81df6363a8a3be220ad23e294f78803a9766e7001b27b1d4bf1b33b77c93a9fa288453db77daf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h316ca905b0d2b9f2464b6dedb4a7b4d78733b7392f7aac9b6cbb96d3f994992c499640facab823797c6496772b5ee31aadd6808132e7d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bb3a5898bb9b91eee3ab89efda7eb603bec8a6fdd771e4080395e4430accdf8c0a2a4b4217bde173e4ef9a6a3fd803d705af4ada6bdaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac9289a063ed7077110843da6bafa4170d65e3d678a0e62971842c90b47d52eec6a43217b918530585d631e17cd4da79a1d07ac68b467a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69f3a725dae10054fe441d31896c5f4ce7886e6ba4739bee419113314ffc5f591fe0944d029a877a5f8944d8c4a521a8f34d1d5a1bbcc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77dc73121020949d3da62574b6c190bec8a8b1cf1e860c901d01286529feccb637a4526d2ae5bbefeb90710b99297d419d6aec14021d85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf340c06ac9cb4b61c7361c266c3fe04c86d30c34f589312684bec44d2275b151cf027ead924b505ac2421837f56a54e801abd34a76f4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1663fb594de842c053375bad9e53ad3d854b4de1027dba1260a064fe6fccad7d4a26579ad0d738936bbe15dec4ae4caddb30fa556d465d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1579906eb76d3b1c971ec1e392a5672a3c17c08d5ed7c2b3e1621cc0bfc32ebbd2b948ac7ae15633a02d43c2eaa4552f33b9043dab4123c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13763a36f6c78a56948ca452353de48ba5500721d0ad96496b76fc04f6a424b6079970d6e64e3b082d493adb91aa06b02c997b0dd1d8a24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6b4db3c7dbb99ef00bfa03d5986b10ed36d957b58d6166c4354e8628bb1ad000c75f0ef871ac67c0e6b3d3f96811777759b171cce5434;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h209c0d291ce53d2b9140fbfd8c9af41810f2bec590bff2e1cd99857e2c3c886d8901723bb08dd20dc4fc8fcf7a99fd353407e996b63d8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75aea0f364a7e6d45cfc2280e2bcb287222ea5a8b1c753b906fe772770aa486101027ef6838b258516099108e22180881c711554a74d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8bbbf0261d91060956e3f4536ccff35050bb465e0b222ae5dccaf54219ddb1f31144ff0f356aed7bcfc5c528e407e819c98c0ef11ff991;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f8c3701802acca15c76d02ca30c7e86179e95fae84ffbb65c5218691065bae0461e8ce6ed3741b3d63d84564521d178f719fefee6cb4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96c111b229289e4b8743a539bf346a4508ee75513d8871203b4cc6e15898653c6316a54320ccd149b756bd786607855b0d94244abfccf0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f92adeb6a74e5f1978e2c052acff3a5ac1420311ab82ba531b48ea07bf2159f1e09746c8b25e390f6c594f8dd1b5a509b3b33eaf8e3a2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h870f50470229040a84fbcd2359f4171a1437dfd05b4e96634138689a52435101d6bcf0176e71b980219e2968259ba1578679e21b4857a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c75a115311acbb6599662b3c12648070d5d02c69220f969e34a08ebb0107020126690c9b0df4071d24ff2f2ea071ee67cf692b68992401;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c5c5ea0fa5a47323f09ce8a274c18338257b67afa4aaff84ee709e98da7fcf2c7b93ae026b7edb0a4860616586f3c547ee72538d4c6dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h933299a6fe34ecdedd3496b962d252c4b101305f16fa2cfcb46e0b1533ea7ada1632f42d0923a26128b5de64e702036802ea076a2925ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c55e96b5bd57d35857e8bcfe5ef938e5bbc1aebf5727b3a50f75ab82b690f5d7fa67e8c4d3f05860077c4f5b2ed8b26bd3f32537ca59eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3a7a389e9913747983ae0fee4b062f8faf2ad1282af59b5e5dc069592bdbada0e9806399b0f4d1d1cfb30e203e9c8e1bf787de28297a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6eee2b94343c753e9c1345d0fefe2a9fcc88afe70fe4385fedfc15f2b3bd8eaca7916a1d683dc182cdb2a389daece5df433c21d383da87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102487161454d9ae80a708dd60f62a3a8131203e033eaaedc1561c2155be0b52d86fa4daf9f56039f8b988bd8b72baf53f31e98e9934b00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a079c85815c28a61093408c3cd9b6630f1eb9aa21e74f61e0708c420c371952300b88f18240ecff8db5ce349f9d70eb1270265935bdffe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2a91dd8f37756866dca4a03fe31e86bdd5b778c423ee7f432f547c37ffccaf0425e9a58d45603ec3789565d9ab0079b04462f53847bb9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc828ee12f171919e94d480118eb0106fbb9d6d30aff5a00b8c7a2e66189e45c87cfc262c3c7a18f89ac4a4fbd2eeab7ab83800a944bf5e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h160cc4e6e647b9060954b6df500b946cd69b28999d7d1ed6f10d2858d74cb6320a39b5cae6a09ea9a9bb43bd0610528c1cd040935628d63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54b0687f40ed915e581db91cea33c2105c4d964d3734b8af94e3392304197918e7f901654d65d365fcc2536a3c5406856565d058ef6ff0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19d4d2944b5052c8d67f58dd5acc6dab8399a6ceceb42068677099afe816608b58cb6dddbc09f3adff88514fbeaff8e4e70366b5afc7b76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h352e52301afbc7fe3b213f1ef9e4fee813fd5ec2c35466bea5f460fabfee1b1bba84f362e95a63df0663bb26c7a8e18022936fa04db744;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141b6ded3a117d2b357474699919d7b76435d8fa0ff5d6a6ce20bfdd1d4bcc72315b6702c5e80063b5020cde3c139191d32be0595c100e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8da26689ea71a8e5647077fec5684ef938be0ae31b7d0b58ac5faf91605496eadb3b6083311d338b7e24ddcf2bcdbb6f22381bdfad1f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d01c241c61d988b07489187d0598a28d6de3235ad0f1e2263c41ed638810f3d02a8ba4bca6de745b7f29a790973054f905dac05c0c479;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c98e0f071c9420e7cb0c5d439b067fc8a0ccb7f007cf629de14c94c5badef79c1e1445ff9bc4994b8b28d3ca547c56a65415a524e97958;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha16c610f2c926de691e4c81ddec0f7bcf538cee89bd421d4d89b81cccc471bdbf9de385eedc636a1c7260c4e5689a127adac88769b704d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8b29b0310a2938bd8c9dfa9320687b9b01c7c5f71e53cc3dc40904b0a6c99b6ee33ac69cd375617a0a4feb35fca4a7bfc79aab1d99c4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69127dcb0d6eb5e2690c0e15d203380f1dd53d3d23291e5d17d72ed8dcc462261075a013191af106dcd9d3fa7ddd57317dbbfc454f9e74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd882785926e9de055082265b03d8ea177d71c70283bc52630b1285b58625bbd3aa14fe9b2d33311af36cf45f7d70c6f1d527dcd24ed79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18fb8f479d49bc4f4a3821670b947e23c08d36fa3fcf71dbed7b612bca9efcc912ef9854932500f69397ac52ca51e71eaa6378acfbca0a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e3f80d4f3b7d177f33d5129c712883600f4922dfb423644d84c87813661fe1a26a55a983055d03746171f2f64c228cffeb91e90cbddf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17564da2f04a3da51e79b6f5a84233a8d6512348e9007901ddab806df2991f301eb0c972ca8fcb5a9be68aa0f86b22e44c724dd167d2921;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f43798a6a1fc3affb1f63dcf14012b588348e1b93550d6ac94ca8191942ad481ff608b03a5f205880ffe2bffbdda0fc648ae8e0fdf153a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haff1119e7cd2bca105554963fd7ef3099af716a06c15666999de5098db4edf9168969c34d31968b7a66d9195fcdda12e5a525cd3ba0fe6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181972223ee03660400e1630ae1f84f629c6dbddeddb7bd03e292a600661012d8a0314a7d33b6ffc67bd5606d801e3178d725b5726437fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41005486398af8311e0f6994b360afbb9dfd93cbc452d89599b22fe9e933a27cf68b14c63c21092c875d53f10a29b131d90be9083e5818;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92ca50228b0363e761685c65208adf74057aa3c36ff957a3988c3a06c7841ad5874d0906d0d2195bbe8d3ed4b1997a3538e3bc8dfbdee2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf8f0cc108205f15aa0db3c24ddb12b71512dca32c14bcae22fcb4897199c3175d34800356d9136cf9fdb4707c22b00b3f8844a78d0181;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140b5795caa3812ca647830fdcd5cbf2aeda392646fc597cf7023a75f5b3996e94b76baab0374b31304f5635c1819ac99bac403b617e79e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1deb9032c64771373aa063978d9e56915e1c9515c313d844b8738f48e8a91bad20662ae1aa4b807184d67fdad1b7ec90e6dc25ebf4c8d33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1950822d69e62cb9d47741a45276fb1fe28a37696622ad55fbfba5799c3719099689be418be8a46db88b6845ec9603d46ca82be1ccab27a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a5d13d7c81a2c8820b49aca4c7edb57fd78ca67a0ec4c7333382a85cbb2e488ab549e7c1ae580b30f60fd41e4268061018b4f0fb920c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e83c16bc7b23e7f09f7399ba1bbf7b881191262b2ac5b22dc7f6e242e5ba5ce303630828df22191798d1fa93aa40733b2aaf447f63810;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186d00ca2b0621b0575169def68a6edde4799f668cbaad818d59e5b9ea96820be89648900b937aea112e9f1d822fee6b73674c64f0c10c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e7fd6a4f1bca7cb30f8c00aba75f270b6ae19d21016aeb484c37b15e9a3b7314c944c07fdd3d232b56fb98c8ac09646b9d7e69021240;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0e9b625eb7c904d88640653593c99efdf64a843c1a5446b014f6eed14ac20fa4cb18e83d99a2bc6f58b044cf6f618906b70d9bdb0d515;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f2e9eeacc7e646d2979d5c052cab921a7d5f878105f376216646d8773c515a56627b317fa17cb5b4be49b30c3da7e23bbcbcf07d475ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10036bf5d350dee29b935a52e2ab1af100ae76c99692c3391f49d79051eac8d4a983d0fb4ec715da38f8da864ab572d64977d6f5e3bb181;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c16c3f368c5c0f5325aa4fec96d4eec2d0717c7e3fbd28a4d446912f95715df95f4a8e860564c8088045a624de35a05151c7baa704555b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20330705782922eaaaed63247d4badd8858ddacc28fe29bf02d31849f8f0c3952e3eaadeff0ac8ed94be29edfea2ddbad682417037c172;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7da86542fc1ee551869e080f6e2f5eba107631c8f4e471b410a433b989182b7b7a0e6b7b3b0891f5a54d5e804cb94fb541265d7a1be9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4f8817364051d35c820ce8cf13413fc783ea51003cc9c7276e40e2dfbb01441dfb9bded1b372c4ebbb37ae99cf89041db43bb7f81a5b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f3a1a5d50c7845a940e466da5dee7482f534bb92291f211f5eddacefc46fc88356a498bbbaed49bb7096884d3b58669cda0056437dd0f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b781712a6f0bf0980c09309b680e598be0fb4d74e197e723b7ac0996c109758f63bb4fd148738c34c14349db0ae1e9c9f5b39f0f5f138;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64cbd756aadfc044e5abf84c17b75398d9be1fb969d5cd16d25e1e18b3fbec725e25c76133146abe624039743eb270866f35c31767d561;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151f6dfbafd3aac9fe8a3567bd8d5576821acfe3dee4bc7addd4a09e625d4e5c6d94be4aca3d523a371690b421e185304a6e5c1fc7931d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fced5f49e7b96f0fe7ae53bb40e694a6608c48802b433b23cf0f455f0321309b2b1bfc62319e70b2dc9b97378f3077ec54042c1075d026;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f7a5db380addc6df8d9323be979fb6939d5da5bb9f04c2e4d87094deb73c1377887a225b77ba618bc7bb7b7b77c4c16a20ce2747143ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130749a1f2f2dcc59a930afbe2a223936bdf21e93491e06052e15911eb86e7e1db4003d46967f9cd62e249c5c6eeaf7a7eaf52ff538428b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b1052f32577d1d74c6ee676bee3cd69f3e1866512979525eb19a8f8e2b25177cdd6a7f9688e746a1bda29b83a1b6e71475ca1752477af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fbdc804a8740578a2833f8cbe3366bbab6cba3a167ecd9db8926ea25fbba178a899f3fca5e76d271d209e731443ce3e43d5c8b75f6236;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a474d1c01d8828a6415e1c80c903f932269c4017d5db6dc00cd13cd3bee5002fcd8b8dafbf05a6d4e5f8def4295c7292368266593af09c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d93227e0f6b630d3fc36851592252fabbfa3f5a28efc317b318d60b166a472870f64cc2a0448fbcbebe5080096bae67ebf9c4d2d97d06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed8dc69ecff03a58e05123e9828a526d183d45a5d476fb0587f676c0f6721b42d6a93662f04405f1f8f6af467a01ebece61aad57846ae7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b5b4709ed8513d6da8b4ea0cb1a06d147c101455436f7c3854e393776dd8ec08b36a0b5dbbea745246dd521a117b46f5e9bedfdd04a0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165352a88285909562681b101f20e36fc5fcb96e8a766061b7b9a4ed3f4b890ed85d8c7e4c11d728626b1940973878f4315004dd40557a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba6142ed0a18449a8798d4bf1083b0ef240d1360db1286c13b68f98cf47e8866e4af43c7962d5f392aa48db969a1e43c7d39f94786c5b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6974a78d944156a0f4c7f18ce85eecea5d974428c50679573ee84042e659b319bfbdc7153e28d43a84ef133885ff75736c8a921d59b67b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d35fe575fa0b531af6c8d7fdf3e88f31038ae37d104963675e44ea6cb4c579dedaa6894a42c48f550ae458c6c77bdbadfc9868e9001af1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8f638a0a53a57137a52f28436dee19740cf7155e6ca627139e64c6a605871ac899e52fd3b175eb7f54b8cf05cf21bd7980acc21c8008;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1414a542b2f33febf835805470e33c93adf860aad413cfee649fb1b4d8e60d3b77b220d6462d92c6ff1204f6f3032f9191c256261955ed2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d02a7812862411e7cfe9abf96826b054177341a3262902a06f946abbffeff533d1f91325f75155f03c28b1d3af05dfa2768521ea742c11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h409e6db019686ebb17e1be49581cca25ac90f18f1361a70154e70d11dcfe126d041d8a9182c2d81e9e3f001fe324ee2a197bc5868c4eef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90cdbb611f671aa99adac08d679221684daf3c3be9cee70bd3d32da6682ef096c13cfb742b073a56d6e76ac6ffa5b5ad7951efd230bec7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c503a43335b85d56992eee96d13c1177fbc8f2eb1106e562a4ed23a1d4f03798a99897066e918803818700b56f03d598c91c512c0bcb95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd55e77bcf8edbf14773c044b3462db8879b9ad779a431eab334c124aa5c4cd899130e708433691a1806a8f6654605c2fdd5e4bc50b6296;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65d53ab65c2542efc16468c1a94bbd34050b300209744405b83652fd1dba5cc4b191e9cc2699dd51005534648ebfd1b98d94eee0f1bb02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f2de55197824c7d6368aeeb13f7763dcbf22ea1abe3defc2a3c96696c553b97403b887c18cd518232bd96d300aadda7c0790f5022b78f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f0c44c624cac14ff06b4d24fa6ea8efd1c262e27511bafaa3e8428f43b4984a7163083dc7f39edff22be6f15ac83801f1b420a1788bd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8fd5ecf2d2f8e58e4a2445c1d0fc746940d600862ab96b314f613505cde7fe03f7ec4743738ecc21c4b0f72c1ecd68f67c7381ed0b9eeb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153f48a8c8ef2894a92c202137d5b78505ed85e2b2127dca5fb8a08ce3b61e6063555919909449023f27fd89416f05296198ba0dbea688c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22580056b4884c61086d8d73e2bcff2bdd2759ba3a9a98861dd3db94c1778c3274e4796ca2b885ceb24ad787eb2a6978b6fae633a4bd5d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c244bf9edce2c1511dd75fb45d4ad8bc07d9a2b11a67f308291b6b9a244fbed5a49fa8881ee1cbb6f14228e1c448d76209be3a904b954;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ccd9b5a9f8571684ee71645688ea6c1cb79b71db6537d9bce8ef2d5e04713850cae337a7b9b567f14ae5b818e92425e2ac75a817e89d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ccbaa490762955aa780a538fc7df748d0e9538aea43b17d2c06688d2c824661b187d288e3fce80d3b8fa43bf748609ca49d6474d89740;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h167df50653e20a2bf18089c9432a9898b970a9684c9c6e7c8127150b87cd79c51412507182ee4fee8ed26af5093f55302f6c5ac9475c731;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad83059472281f618604da5deaa78ac214e64eb83c573fc1acedc1839d6d075b0f9a7a7fc2cc9c3863b32e47c66c56e01ce3b617cc88dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e78ecb9611c57e7f2c30cffe54150bd5c7faa68b5dd18dae567833cc5674df097034efb9e08dd141e5d857dcae6a73e21b93713b51fca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d8a12a4d2ba10a402d7097ce744f44d63502023eca7813c7767a46d53fb5c03a0a527bc37c38d99d28ac1416d9b078caa036412ef97ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heaa13fa28d73ca5f47f8e15930c7ebba464eab1f4b97328e641f1f7b7751fb2fe77933715ef915875d8688f62dea7c4f198f4a907cf82e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h371a9377d6cae13af5ce50f2338e9ac0dfcff5839de61b1e59cd311f4846292f6f058a7acf7e0ab65c68b408bfe4d0c1b1431214ef5db5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c6569eb963e2eaa503419ff5ed52413b172cb05f8f603b1144d9180fb86b9fc691b72120d1c62caf36ea3ef84787b765fa637462aa784;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bedd7b51586e630bdde083a1fb89e5d513e26240d95ed1e425e92de15e2a4115388982264b213e3f5a1f9c8582a8811096d7bfe3714050;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfccc2f96c2845705a6f5b88e55e38793e71bce2376579588415172cd0c951279c20100af7ea2b750b701be0140dbfa6db33ca1f9a670cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2500d3798970a91adc828475068cc8b6f296ade04156a0fc428a20799a8f284d5170e78c49f9960b27fde27df012a67897a9cc6a1b5ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h143e9207e3651b31aff7338f72e4db5c9a2f276d9ac051dde92f0fd753db71baefd2e9047f1486ebd59c3f8eb3424ec8784f35aa671c7b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3198395c9db591cee163f9ee16039f36c69ed772b333b55bcd840b6deb126854cf79be1d45c2652ef8bbf37876a65d1ecc60f4d0c945f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d2427aaf2616d324b4205858daf1dd17a366c4295cf38ef4e1dea57bfe1badd51fe6f718679e51c79fb5c399c4a6ef27324e22e56b589;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc04c96b746fba73ae1fa3b6f65d0f3aa9739211ff48ca546a7381ed03d1c1e2371d9c0b558139c410aad7bfc4afa3ce33895916c54ec6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a176961330a32b3b1c214a94d20dfdbcaeda4999eb1187ecddfa6e1a499ca345e090e79e4e387d75aea75ae0fcd87f46d203e9587e0725;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf467065797eebdba340044801bc0135a07a6616ae76110d5f45c39d60bc9f8e25687877b0dd577500c7b4665ab5e5b1ffc85c4a17a9e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h614dfd84ad7b67a865e1c734f4ec2334b48a7ef3f6d277128f82ad62b0dfb61ef50ea187b16f1f56d1d420038b0f4c9f42b5b10a47e8f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c38c68203fadf0cbe283b920172e2c798f69678eec2bf47c8e8c55c337eb279cfc3b23896f9c17d647d4ca229af9c92c283949f218a6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc37357ad54538fe36a49d1b64fb231d649ab488c14909b1d73728ed7b9ed3194a4dac051834caf58539323024eacf9bbcb4e5bc316e98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa9f5a502c79d6c470cc4e14520d211e6c09ca8e5d97242d26bc406c19712c213a1c03437e04d15b7dddbfbe68f33d5f4f121f63aa95f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef42ecf8926bb68ba2621e6bcb8dfc31a54670bd6d2062712d5e7821623d97bef3fd0d3ae48133a31e998eb6004dc30c4ba85671bbea78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54f2548d9d6768391e9ad74ebf034bded8d51f1aa9329cef1dbd3b15bf2752ef879a4eaf91236b5744a1b882958b410d802e0d6bc7d89d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c6ee4640762e76b53bd1a83ad3b2e53e58d63faf1e0577fd63e8690a4e8ecf17e8ad8cc33423a4814fc7097877d2c4b3023090592bca0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d073fafa3520cedbf6cb97999b6e2ad2e5effea3dabb90d4f4ce1f2a55e2afce848aaba5d2a62e1b2f25a5b3743fd72c3bcf5eb52dd09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc784a2302e73eb5321addfef23cce05016cad1a525f4447b44f7041a768dbce83df20a8b4430fcf444310183d7a50fda82eb1800d334b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca75f10f2b3a146d5cf5d13954ca922042107b1d15bdbdca3cce504be9d95f1f672a725f74c5d860e3e13cb33d2778dc98741e7a6551a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ec6cda4d7c93d176844d7dc91e55acbec2939d9553d947d8c5cca7acf81dd4e57d6c497ec0b53fa23625a82c7110cc838ad1398117320;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6005bd92a5e3e8c737333c30f8b59719f7c76f8bfccc5a4979b34d7b0ed722cec6b42680a41326f3ab61af7d18c598de7bdc40d03956d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8873d458325a413d7640134a9d3275bf82520f760d900ca7e4bf8cba133274031bd4e6ec8f303f6b222431d27753944a367e5b699a9c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13550285beb29486fa97ef2ab98cf4e1ca2d1e2902b0392e41b5431a4785662e3bee98f2859acca13a7e1c49c774fbb3001eb12b5af5e73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6fb621ef216b8a69278e88ef807ac770900fbcbb5d271037ceecff82a200205cb4d2a218f4a8202af1ff3eaa5615ecfa738dc85d1ab29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc992ffb083e7b61a8d3f873c97cc0b61d05877f062a7bd03b53c17166c5ee75e1c5fcd6ab0adf577b54dcda474cc954279700a807957c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12cc49d2a49eb1c4830f07a6e7bc6788826909aee139b8c195bb233def3927d7ece849f231c49a2d816e8d26ae3626444082b2fbd9a2a06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126caf4fc8d15eac786e1aed26e25afd994c4e217ca12fb94a97b58b00f217fbffe810c8b37aef71eae3cfd207fed7d2bb1b9257591badb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb588d0491a8968024951bc7b615d45daa55b2be253f881e405db256a2d5f96efc8ce04981c1de29a25752784f9387c8724d06e88ffd56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81e5fb6325531a3300aa8c93831636c5942adc9817c908e14ce4859f62ccdaec01f5a460dc627c7dc3110dab91ac040d31c21ff4026505;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8a67f0623d46cefae5bf96902e073a72d0dfcba85731482c4cfb4bba88b4508fa57f21abb0fc990901fbdff2e683af5027b3ab3b3f612;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1574ff840391295959b94c1589cc50a45f4897837bb8312914214a05b969726949695642c7b6ee8cd9c19403de0af3485f971b230732e4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d21f59bcdff7bedb69cf0232067f78ba290815c1aff8b40844e1bb30e673f1111ce8fb9660cad74aabd8d03be13fc7addf6ab0edcd0087;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14742da37fc38b6a6c5c7f417ef87a58bb2ec927faffe936608d3142bf77d60009279dd47f94ae626c2a32b3505a71e881052fb7da5bd38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e9e8bf5b694697eb8de42b86f59278131fae3348cdbbdd20d6e9f004d8a3fbd1316547bed053cf11a794611e0181a542ff96da944d1edb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ace8c57c111a681d630647c4345c2c7a28b7e46fa8d8caaba80c8e1996fb815c414155d501b3d5016cbc73443efb811480fd01fe77598;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h272f99c6d59b8a1eb59de24539963852b34684edec3540fdcab471401ab0de8a7bacc84d5743367e6933302b2980d860a7456522d233ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he31528214d9ce56b0b7bccca4ca42cb08316075fda4aa6a1f303a48d6e946c4e799da967c3499c83b6162e21ab1bd58d35c1850760a5e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9153396052e0014bd886335e2a6d74f7f4b883de0ca9f4b112083f3c3993ef08037d058fd36bd1f39b74582c8fe6a7f6d755062a54607;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ac4822476183e729cec2d85bd7aa955ddc492ed2245a693ef1fb119f789ca1faa4fc87d001719d6467cf1f562eabf013103c40573bc33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce54078c27fd7fe94641c5612e1643ee43895ceae94e984a873a69db981f36d6756d35b8fd4ea0d72692441f73ee5d421dcd043cb8c224;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afd0e6a358b241bdd0a57a3373f7934ad9311285adbb7c90fe66007b32810fca6e013601b4b9e330f8b0dc1a9e2ff1ccd78f7ab2e883df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haffcb7222f1af8e15d2649ab8be626062c10259c0b58330f58cf735bbc873d82bb3c160f5e5901d884686399380b014c22c8511ddd1022;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h755186d75755a98214ebd0ad5308f7828c3c16dc9be2d851f1980aaf2f4ce3334bdb1e994566fe840a8cd97bf087e3a3f775771482f316;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70e8f3af122ab09db7de577a355cda509dd6d62a8e95835a1c3cd0d2dc8f12b2fe04bd76f90392831d4f2f3f558af15e518a10ba4267d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cef934c182fef4f3c0fab802f8dd5eed1c811731916830ead6fd70c78eacf44002f88d74bb5d0ba1735009cec758a205143d0847c6506;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8eaa4366c43d9552b28a93ba789cbf8ec90ab5905e567180e4a3343860f41d8899ba8bbe09e62d119700296d247b787e64ce1015d33076;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2ca7437e62f8346e143467694f4ca7929b1514f257790233a17f4ed7fbeba4c7fe31b491cf95ca1b18ad6448eb41cc8af39fdf3b02eec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3eee1bb74d6edca06b7b6ade42f36637b1b6932ba34f413071a6d70faf6260b8fa1e875dc7bd9895d3ebacda4e74a625d79e9f6f744d2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1182201d9c22960bcb02d6be95cc4a724277c1db055a4d8dec455e45aee39b11471526154992413b89f4f04ba8d7f3ec8374d66ddc10afe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a2a7246d99c885b9ffcc799c3219035ef23f9dea8c1d75a86ad8295cb045e0cbaa7c08cb1d109b96321c321bb0990589ca0b95ecff9a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f025ef6fa97c9cd759537160dc66085b0f66370f1997b726a9ac1bb72fe214250a0ee41bdfd2005ad7a44c4cc97ceda271de8c9aedff8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2bceccc7af8a2892e87f6c863e0e18b80d2391e72e55092d175bf781393f0403d96a526bdf6d920b371305b49789e7009ef8725d226fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd65a6054da19e94e912c15ff3b3d95f96f5851201f307758b7f26dd2915faec5a97f68b967e2770a16c9091e054d381180104a9885ed8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171f981659615c6a53d6ec342f555dd67938c78749d74055b7305b2a513bc1000433d6db72fae46ab9288b1c7facf61c435cee7de6d8935;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92eaff1705ad82979fd2d1c05cd0ae9e5bb9ff635519e0445d41eabc42b666f99f48b6bcf026dee7df044cb74182e81ab2911e4dc964ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd10a8cc23d6badd63b1616168d787a04ac266a6069b801c9243dda756d37b9bc230982106fe11bbab44a76616f97c309fa084458e2c9d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a7f874a4500a3abfd81dd89af01829c313686d3aa5d887936a5377f4aa9b4f7612156e1d865fdb8091b7357e2f9b33f166ee4dfd63085;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c31727438fd2f3e6f991cf545bb6e2d029f946b730e0f31899338dac95c49ef3efc7755db138f0b8c818c26e4279532acd4afccf445bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea376e3c47cff075b77c2cc76b02028313ef21d30c4601d3e835ee47b019b13570b0c5ed12198ae27e60ad8fca307960da7fdf9e096da7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d7b864d569994e7093e98285e43d2579b9d65409a6030ae7512175ac4825760319579672c92e7abdb6a51c592420c7973eb5c84fa3ff5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h642dd2996a23fedb9a2350bfb3c22bd117f078730f8656da9567ce0b6ac82d8bfec6e00b5805ff90fe850c1f5939b337934a6f28b14714;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h403048e20cd918ed2973c208679a642cf2eb436252bd3d05f128d2b1732e0479d7ca1a4cd327640b3ff9ed73093981adc57f92fafd68dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeac90c6a620628c3a2002bd9ea5e3c70e52573ac2ffd907c6f2a866e5f4cd9aa27f90d62a88b7c5053db5443117bcf7379bf7acd4d1eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5c5d758693581824db6cb21c877fd38fd98c77a082ea9da57cb92efded5381263bb65799217fff2fd15e584f9b7a7c9074197ca8eeb8d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10915696d4894e013e5db3c643a107009cea0aaa87072a1f3128bc443d8e9d27384dbf2c3797e631d2781882def4560d3ac7463dd2dcca2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha265c58b87a58eebef619675078589dc87a689ced11581cab5e668eb949a4231a71f4d420db769058993c48bc2b384303a95c2a5e3539f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21d854457ca34c40c7085cea9ce03167e46879618f29f1ff07ca25fac45e600a51330547fb1f3cdf4c5b5fb25362aa5d3e75b067a36edf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f97d67c09eabc0491554010e7f4d3e13d7bb6de78fab0b7f836b819b613e6203e55e4cb74814f1d4bda0c1f5755c744fcc00caa3002693;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17116f23812871a8bc82a351d0394d4b7311d31cd2b681addfb3e37c837f9f677afaa91dd3b42764ec31b4fd1a0b15cc46ba0007f7d436e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbf2ea91882b1132a881104dc960e00bfc4ff7730835329ffe74c56414f094a629466fcb64fb658bccda0b3e09dd7f3d331e44000ed252;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c60be59ececf5a4b7a488d27c03a8519679034d1b4e53d337a63515b65657c5330f7bdf729d88978e6b56fe1eb757059c7739e213850b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b71613bb6872a7bfbf40d104c1ea35f607af5888a3163c19e7de244153e63bf3a9a35ee01a50904f0461ad0b25a773cff8c238712dd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123be7657bb4243d769c8c570a7e70b457cf3ca6c58179e15041ba2dec2a97035514339f512da6d86aff5f20b887311a8ad18507af7fab5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e74c18bc9f40a04e83cb9ceda55d1f4a5f43c133336843b0e10ae8122360b0d0f5847c02140b1faebb60fc758f9d00575002de0065781;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1f054d9a8811eecb285e78e40d28336a3057abdc467189f1786c34125e88fc22058095f1f1c1a003a272ba5af699ea6f04fbeb1e0aff6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e4a1ccb4377b7ee78ea1c158c06bda146c161d83d905551c363de4d78045ada03704af3143805b403320afe28e6a90b304dd99c8862dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f14e0620f9ea3d75938e98a83d8df8f304f0db057361269328ffef11c0017b2103204acd74edbce87f268a6d4ceba58d89f70bf7d39be7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h743c38dd159812bfdc775e18d3698e2f7af39a6b7cb0706eee42346c2c364f6304408be24b75474416a7d5e2e3de25064b36d1c82c7a3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5c640e9a414f740fde3f03b29434d2d6fcc1d8bbea7e34975f535ec90527cdd99c72bfab362bc8ec22f22c181767195b1102e033d5de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7d8f32a27cf4d816ed343a96d5cc71cdd529e567139f32188b9f2d0f85a180d81e8b9bf1e248ee9e27888fc396d6829ea7a193693bad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d98307a1b3e99b3bf8aa9b45d4f90fdac13d139566e5909e6271dd5ae0aa16c3ae32c0fbfd8d6b4b2f8d823dcd74c981921442930f663;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1517667cb3ed21267fe3c695401c4df04e42e6bb65f5835f5479361c7ef786bc161b50b620ac4a393671e1ed23b46bdd75bf6b606851943;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h731d75504847cd1f345d4900f95ecd2d415837d5d20eb42fb919e8098ba3e915d9d6afe091ebe33464265fb02d59b1d62f44d8e3da7cb5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b05b5abe240177f318b85b19dabeb98dec1b573557d9f38f3bdfe0c895edcaf017429313654ea1b24640faf655b5315b4fb781df3953e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc897c1759afa6654fc8c8c3b9c0904e8084b51b2b5273af32610b6a9d2d88a95224e4d56186e29efec70d40fbd87515d59720e75f5b3c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf555a756c25b8c959fc1f1ad9cd0df814b05920df0a4643c92e49d53de539c74ffb5ecec1dafe8bb8fecb2ad7af6d7f586cc2d198080a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3bc1c40c46acb1bc4391ae2d6a11757cb22f39cf56655ce688e11fa6ec494a560aaea2d4b903f72ebac12f1ff9759940e7c7137771d7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108063c3895537ecbb3b0ff9f1d825f1f9ec2c6d5ecf9dca2011b75352c623ced7ec16fcbec96830d5f87a8cd65cd7a91de6ebc42830203;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35968862ef02cf2b387c80638499b7f76f79ca98b85c2708b06b107d11dbec00d1a947e37f2d3255e4f8497617f803e9eae3cbfc215300;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140565b08970bed4eae4751181ab48568dc5426a0562b4e98f3463b91838865e0a6731f717f25fb352c9e4a792396ea8c9540d2e72ee177;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9afa1a415683fb71455d17eb5e8fb7f6d9767a85dba4b84399eaa878cc3ddc05a65909d71649b7ec55c0a5476f1b845f5c06d757130582;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d6e95dbdf9e98a156ab6b5ec1203f8b1a64ccea2fe69c09827c591e4e522b3220bfc1eec84af0d10083b2458c7415a9db2e54e661c8e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea7cdcbab257919b592beb87f6380cfc2547c5c8f9de50a77e3b894ee808fefbd07e82361305dab360f6a0d0baf88301fa50a4b3112101;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71a7d108065c155ac0b2ffe68b5bab05ddcd871bf54b3a73a152f075f6ddd1b4d5f6f22262b8dd69b91d578b7618a3bda1102099b9bcbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h266b833190593d8f4302b0cf1c7f566f183650bb9a5fa0846333f1de4adca4faa17cc05ce4776f50e75041b34cbdcaa5108e3fda5aa6e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd4120d1ed104f50134b34ed3429a1f25b96568e15dcf26a424a56f46dcbe885013df5ea9a3e6b38bd7cd479d3b62a0a4d8b6437bbf0fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb08dfc3b430cc84bc972ea8d9b08b674e112b452fdabcdad3f73e7c4ffc36677fa384467f91a70719f7f8fb4d72fde72fd4ae328f307d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e01347a526c93eaf70b6ffd630c0c5c1b516ac08761b0cbb7195f5d6b9c93e145df3412c853884cbe5f702dbe1d80307506330c58d690;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1069e7b93a922bdd37facc6037247973b72e227d32d77240873a2a9d9740cc7d976d4136f2602724a029fc1eac334580b47185b63516fe4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb664f4a057ba9699aa24e14a666338eea9aa1e49b72cdd1055ebd9ddd617f3865a014e2c70b20500a7d0f06a81450e646835a9f9ecbf6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4a30c63c6b3ac04aec8b05a495dc30fe22104c59368217493b571c8b2a0988d3015437225d7d9fb230ede5cdc187f297e63fe42816b95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130078f559230785367aab4faa9ca93a18dcb880728316c147abd039513ec7b956acee502625e67faea2a502b3797513e325e39683e4edf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5eed212a2c14851b49bf03e1c16a2d01f4c471125867700580fe457b90dd33f433d3b9fc22bbac01ca83d703f23d1dcf25565dcaaadaaf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a0a18f62c53c03ee2d895319d3c63d039f846560b93639501b5158cdc39f4f57a85d254f92baa9c0c7dd8c9837c9791e6c22e022cfe68;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae99387145e788db7ea3e173754f9e27a31afabb2eb24b51330fcc80bce505ef5018538ac6c71f9789fbf50b936dbd87b2dd102d291bca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a77f30aa8602c1d99828fe304e506ce5e60ec6772ede2aa9ff43944dc31ec7b9d667cb959e7ab4f642d3bd4d88ac738dc4d14a358efe0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb7cde291ad6e725ee234475eac647b6919cc7ef3141208cfaaf11e9e9c66476b0eff0e4b3f5834bbd4515ca90a07e4e871d252006a229;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1aa50cecf33b2676cb044c6ff4c4045681b2b9bcd4ab658abd192305ee3fc82f7ed47b5122a71a87c26b63025cd60b9d956ff411c31ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92ceb0fbe747a7bacb6dcf84b9228294db0a301704074f4a32d7768987f4a8aa0a87594fe85cc9d00dc92d6eec5d1e36ff5d7cff8452b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1431fe9430319531d82275e2e3ca211272181b95f1f5e5f6e74f72a21bd11d5362df74872bc2d1ea4478eb01d449ce884db4a551bf12eee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e903f029643507618792036ac42f6d6b93348b93060d17373f39d36bde03f9c7123e644fdcb082b40631bf3e9a694ad6ff4b634287f953;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e738a50a2fb0521d1d49eecca1a513c616b9fb729b01a120e1ab908ee4a394d1044a31d6b22f013bf1b2198df8036d5d490f564addd5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bbf057828d43f545fd21ca4ae60f5e4e1672568410483d98671659f8150c61d423e65e0bb299feea01285b5d11516d9bd51b2ed3a54f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2c3fc635fa075dd47cd02a8cd1d142ccd3adbb9b9420dded93c5e14ca561b6d4ed8570fa333fb4d5be9c6378e3a91f72bb8fa938d1b04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b515e7288a8fcc7dafb8c2db9c7bdfc4f4d68b94152bbb4da9100465815a1a2638a301c81b1cd7465055dab3928272b79386a8bb4451;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb591e8b96d05a123c2e08e7fc613503846f91d93d2807e38a4c5ca823080d78b3bd15f5f9202e0e6d37f02293e1ed77da30d0e9b8dd97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19713a728663b3901379b8e03ef3d7ed5c15a24fd3b81bbd7658eb959e47fab72260498c54f3b0814a2dcd03815b4d9012d51efe4839c0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17834442bd8bfe8e163f4a2a4defc8e2cdf91d8c1042221b027e21f2a1a4a54955f344fae275eee6dd4639fb72fa5cd2c83cc4997a4a7d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3d78b17b7b47e11fa7e0c6cdac1b90ee5233bf14f79f6bafcefd4bb6189db98ad0281028066f84b26d8affe42bc6d6ecf47c6a26fa7de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f122be8120aff175554765fb0934c62b87028e47df5d95bc9ef7fc68780f890d07e045e70115db21bc91a0dcabdc8561620f8f29a12c09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9bb7540581608050f0efaeb82ea96c332973d7c2c75e966dc367d0b9972da1bf7f55df420811c365460ff8c6bd1d506151481b1885361;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc21d4d9150fd6f52a2f2420bf081bae21ad05f3fe066d55a1f8c346e5f0b95767005393718179320afc88480d93bb0ca689fe177ce96ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9807675141535ac4c9f5786568140cc86d12521540555bd943b52e6215bb211bcee747d24a5e7460c320ccb3d70a008b95afd724a6e88b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d881face149957677797270fe4f9056ce2e8fc6837771fe70283af4298ad13de9c9113324c2bfde2d3a67f2ba3b4a543fc57c0e904712;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d90432cea4e0b7e1d0b888e6213aea4a3e21f2a3ff89af2cb88fa8085d85b1d1edcad36f0c9886ad4abed1ba2754e186b377289725438;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149fd34ccf7c85f1c4c2476be0d58763c4f24f9c7bbfb0582620d550ac3b4b3ed8650680f47cd5600ae25878cc650d2a065b90c4dec93d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e23431eb695fd82f885070aeb2558b46d103616ee6a2bdf0043e0b5d633044a06fede875e2d569d49cc352c38906da7f467d8ab449818;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea58a1a13f13c14b26ae6122aa7be0934e98e43526c06cc89a4090f0d39d62a23991e6832ef63d27e3f8ed0c400a91096712eca7489a94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16939486d43c2ab9578b12db768ae1d1dc5e70813ad84e211fec4e546cfd08594a1b63c4206a5f53ef60ff7345ec61f15c663ec2c6550b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h814f08a2ee0aa0dfa6a8a1c4ddf88cb2967f0c4b162fbfd579994b1a60f620c114dde7a27a382d6c0f1b60539aa7806ca89233c2d2557d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56c530fd0725b4fb9baf6662e8d68f4f6c0b77d76a2807e2c95472f77b418ada4064ae0cb92ee6a645ada6ea0bf4408f2c5bfbb6d02db7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2a8ca59823e0226d4c52c4a2c77957614e972a071edf90266d68e9d81d90e34beeb5e10f5fdae1fb0efb329053081d3c02e93a66d0fdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a56695c3f48735856db4cf4cbb24dda3a8723672c6445d7dd0e8dbc18d9ad12ac5e1babe77f50033a821e11a4ca79e07ca34bd51012374;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe05e16513e02d978755c4e2ec7e30a3ad139c60db61b45ceac1ac817209653218415f3dafb7931b89980c4b6ce5a2c6a6ac8142f9391b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c17afab4646e2763c8ff2e351b28fffae770c0aac4308c68784001972b0cec94a9f59a75cb8215bb6983ebfce533b1b6a5db66df9ac28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175e26b00068e3f0f35a67e9c21f8abf6e00ae5082cf04521e06869637c7a266a88cf87d0e0f9a985fdc48bf1dda44fba345f6ecd914d5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8db63d0c00e6d91c9aad4b1be78d8fc6d8deaf36bdc346a1d67bc2f78739ff2776990de9806d62bb9ffcbfb48d0712814d56b3f710e1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h265227fa9a550db045a131189cc77743c091394656abea145126a0acc93480caf1cb759f704f1b12270ce295fbdb8424739f5fe00f6e80;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e99eaece514859516bb332873b00819cb869045543332bb52130fce13d02d604d175ceae3364a2d3a507016285d4197a785d8713cc958;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h279c1b429f4c18099d5d5ad879c9a68d3b1957bd9a00a8ef2bc0d3315c33154810ced1daef8de6b72aca29b6a5c5ac2d08ec851a7dc0b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b04d238dacc04036c08207c67b55e5a271b17ae3df5e378a2d4c01cf66de9c618d370ca18b80c2a46c205537a906e06ea6eb8b3ae78314;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd926827f19dbaf363fd3de281324d4fc164841189c3774e386395572495056344dec9c3b169e916cba24fcbe4b586e49db8edcf0a00e84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bd756066764be6dd950d07a1ea6a530f2cfbc90bd09dcf17b9a8c9c893b0e8919cbea5377903a30729c290f3f179e8a826a933a87f164;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a0743e0a2704de6b0b300ea6e51ac7a15e0840493087edda6dd4802a0989641c3002e0614ed73881c033ecd3681c4a44ea8cfaad2799e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b296a440823aa70e7d286bada13f4e85a518e3b5b3a719d3ec3472a9e6959141b01a551f58d43f591a82dfcc9c1cf90960866c4ab73830;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8dfa88298efce0d6384004eef4b02cb3d548f25e698f610032814d42af83f938bcd59db87c1e708db42502883c08b5495850ab1276c7b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd76b1c6c763471d848a38f94fa07c26ef3a1e40932cb64a0506432464f6ceb35608e7d76ff43a772996150440641ae7b56be44147ffc3d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfdd0460f20e619bd392bab0ec8da1751bbce55ace3998b62b0b9bf32ac46f111b600751c3385b51de745e262b8aaa6876cec386d2f329e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0370c10d41845c04c5a13f465111120a913509a4a60662cb1a2f31be4f7836d51a560d13f5381aa3233883316852d932e7ea136cf43b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112b54a6f95229ea53c1a02c3214859bdc814d40d4c7bb4f7a29f89749f3a56014902e63286fb8465b08f2cfe94c9a953acfac93d0c3ec5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5655450e5a38f1d369d983f133eae357286fcc482bc247eecd911efdc0060d8b02f7696e3cb0998ad4a45ed7b5b2b8484324b8a9eb347d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f323033d157513b52764620572eda5cd8ba0032edef0c99232a30e9930784f71a618a623bcf4feb010bc8022eb121561dd705116766758;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h884448d3b8cb253f1fa75ea10f154f1a76a75806cdffde2b66e484eff953aaf4eaf4838578096b530bcb81ebc800a16d646f9b0099c692;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha632e80dba0d775e744ab2491e45bd2ff3b25b80c7e8657f15819ab945168537246639c3189f29b06472c30f767bc1a1961f049f49723c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4f1fd27e6b2a1b31b9f51a7004e7d31fa14e6eb7572a86d1c8a0ba2604c58eab507a2829562344b084fd0cd4785b8a638c1f0cf7b8abd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha39b9042aa22f1fb0ef25b5be6f5ae131d78a7c62531a10d6dc91b9ae2b44d035176d547549be4f87e571afe688e69c0b344fbdeb849e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee687329b163f276e8854a059184bf5053cda4bb1347a4152f68d1a0d5cc20e94f00800473794fd8e44d5a95a089abfba92d7e6a26bdfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b116ce59854d80ba41408c2b3953a0adbb225c3911c29bc770a165652363e9daac31c2af734030ffdde283be34907a9f52dee2ff53e13a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f6e8d4f644d46f01899664ac5b37ad2e4055273a691cefbc7afd4aa5efc32e652962800f0b8faafbeffdd6048a2db87340183cf57e3a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f5daef2f100af9e20d71f61e2937fd96d352ee46df87b043752d3b7616d197384cddfdafbbf91f65d8e5230bac6a9877800e4880bcb31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h822421758abf4e9c77b738b391481fed6e750b3ea01cb04515a01bb808f0f8d0dd9a527a14d5ac13fdd198fc01bdbc7011cee2be02f9ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e073d6718b8fc051276f0ca31e2721c201c5a4a52f32c5542f29421f217c9a295833e877ba5f6aa141ef487667eb8173fcafa2cf551a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1740dc90666c5ac49888643bdc0db4e8de89f812aea3cb5faaeb9f0395b31c105706bd022f1bb6b571f3fd048af0ac65a336615ef5f621;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2dabdc4439a1e1872e568a2d9bc8714618232e498aba02565bb48c6a7037f9fb0beb399e7447dcb2cc9b700c6ffbebe3c5249c23ad6a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1217ab6d7a19059cb3394fa6d5e9eb84e8a0d12086f3ab94684030f3100fbada26d6d7bd5809620b41f9b0460a098dbd7e0c5ffa494d744;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183301af9c5bcc504e9710c5ef43f781e14441db4536799dce5052103524eee30f81bc3338f3265568982867ed2864cc729bd3060a26b1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffc4457092404c66f708baaccf6d3292a26a56cdcaa5ffc5505c5110f128d857f2aae01f2775533ec4386c85688afcdb203590970ec220;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1695bb048cf25e53b3b4fafe22836941001a02ef5f978ea07ffe86d9a97561285cfbfccdc6d75ca8167bc109e541d2cb319a81c039366af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6759e45762efef79fe626164612bc989b9a899db9382f5f2eaf4f0cdc4b599b39b27049d350d015d66fc0ad606fac0031cc61c670d9b1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fc093f28753bf865d294ea21fcad43a8c4f26e9824d760f5605b4e89a17b39b972f4ebb3fd5e06c98aa111fd862b280ea657b8680f7fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1775e30527a7e6ce7aa6e196da18d68216ea22a51ab4f208bcde125accf04c391081446d36e52339e0e64584f2219b42cddd33bbfd0fdd3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0a12448639f90ee9efddea8d27f6008ab7305e6439c6a12b5d35e579c97ee46f598e234a061241a298675928f749bbe8ebdd09b6fe427;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h515b3b16fdb467e69b29c6ea7d89d33d3381958ac91d9ddff42a7624a31e1c3bebfcad37896454865232957009e2a74a93795784200332;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a780d7a340a14a7c31bcd3a1eff85e989702ff506259953b7408e5b7c33cd1e6c458ed7f20d17eeebc4cf13cc16ea0c329bf264b87605d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha71764337ad1710777d30bd40ee6263f495a922f0f6d99de32a4d768cbc47a6c7a05c13f71276bd3229dd6a94d75d048c1c5a8e2bb55b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d1383a15d7bbdbc7eba97094fa21f53206dc04c3f5e0b6e95fc31b6244d73bd385bd37802b062857195d217c9261f4f5aad34ba275ab1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e911fb1f0ee9d1aef0e4fc3087fc8970b2d4866bcfba72ed8657e5e93e32b4691b43807cc05cd2388c6eb91a5a103d7723ad0be411d0a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ae50cb8864d833dbb26529e2584bd426219a50b5a76ba95ecde1c6cd0ab1f04ee96deb5811c2ed32ac616b5e55ab49bd429122158f291;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9562810514509d9889b7036a54b0436fc478a6fe6949d5d1bdf4e333cc86accb47818944957177016fad6a488f15c59280db5cb06ca65e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c64f1a18abd9f38ca3b6a48c20689a43839b9d9423329cb1f5dcbc5ea6d7be4df9faaacd4d1b0e0bfa68be3c37df2e63477e2c05ef27d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf5fe4d6d4ea255def10af2e17fac3fcaab43f434196e01fe0bc4de6bc27e08b38eb6315cf85d2131638e9e776afebf426a8e4ef66946e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc976f4fc4645af23aa7228edc1ae62b9103ac695412941bfcfae7bdeca260c0c7576a05585d6b36c5a87f55b8cdfc3703286a471b4c827;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18dda8b1ef7e8a64f98566cf6b754a775bc683ae93f07730cb71d8a3f852996784e4c79335f3589e76c454175d909710cd321a640b295da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb53773a0b770a24cf30768326ff25987d003996f2d1b8d0592860da7728a655ab612c9b50960818f20a55c5b95760e813d582b939113a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1193f620b9d186221d31fa0a1254aa670c11318269d25fd2087d54f119b8c622fbef5d7b3216647d837e3748b14fa94307d6b46a09fc3e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d0e4aa9b636c467e6a4db8b11c5768fdfe36a1af2fc3fe629f807265c0abf9705e43424e01d634082b6bbba62a3e55a184464a8252820;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1dfb5022c7b306e68448a65f9afcc2f10375d02534ce9885577444c00db7a98b9818f589c2bbe099ed3fb5ae6607428b19ad79661e362;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f937ee63d61f14f110bfdf4e31f2d73f21994a2e7a2571096ba6be278f801b47a82072ad34eaef6be36f7e55c36f882c66734992f9465;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3992ab599bb81abee3bf4a8a2dc0762b47fdb4b69caee7bb05d9fa7d3fd229137d6818585188fd8e2ef9262082fe71bb884fc78ce729b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha78cb388f18255efdaaf445a460ae6b9cb52575ea57788e0f69cbd41c507f85483711fd83c9a5d34aeb55a24019e6b2bd2b366566a41e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99b76b4c634920459402617b8b2b998c7c97477432e137787104d9919fa23672e1daf66b393c5a16d2fe90bc88a4c950717c0e47c17bb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130f45014baad5037b2017f4276516283e78d70dd402c78d32a3a9e4e08bc15f641b0528c4b381c9954cbea0a3f41840b0e58a49e096ad2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89784908dc0b697160fd2bb9bdd2aed4f3d12dc5291bce3409bf2f418fee0b08eaa7194c22884afb21f2eea8f928c572caf448622c7f5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca47b8893fdf8fa7817acb4e8aa28fa4d70738a2c18b0071ff6a8d5c3d64ee085855ae5d4e536011451e655b2e8f5c02205f4cc625b300;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df017dfa7ac83ce803b9ff81d2bc4190ede7f9458cb9f4c71c890adeb28f4b07e33f4a865c7082d7473cf0af56fe7e8abc32691dfbe0d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39b25236fdb9821f088e962a38d83288d3ec7e555eb0e571ccabaa7fa3d62193fd714c2241b666e8b28648a6377cccb34debb22e0c8784;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0e71e0bb937aa1fce5ec9b9f0d892088dac72f6b92a653a66281f31da426ee421e5f8dba9a28d90ff9150443294f4f0e4058862470057;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h383ea1563ff902d64ad019a00c76974ac2aa3e9eebe177bcdd2730b3c0f136a8546daf823d9cefe9cf993e945ff2125aa4d2a13bdd65e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182238b59ff89cf7d4235ce9255dd9462154eb43f0aed78baad35e03aab923ea24926ebe3596b4b8f4211f708e729439313afac9855c602;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e277f64ed843ba8ef5ebee22b7aa196073871d37060ebc3850c46e615a7d3479a6c1ee9938e97c9027e894d3e805c962f8899a1f2a5e60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109f5606b077aef755ce82ecf428f5bdaa7960bbd8dd6b1e5d9cfe724b05f39039deabc673202e75efe54fb0a98a9b617d59abb6ebfbb49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168344c15c51a3f374f05d03b634f24d994405165d7e7eeb2b5da1cbb5ef619bfc70788a4e9fe7bd96c5a8bc07d2d81d3325b37dd5da25f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11482ccdfba3e5fe8df56a2654337aeedf7cd5b747c169fa7befbba2e2f53739d562340ceeb3f1fc1c84a16c7abc17b67079bc6dc18ebe1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9040934cf8be283ac8657bd8a2f6fc5a746fcd0878c0198de91be184b77c5c9403295d64075529efad968f8b6de2be9f0d5ee66e607d29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16805dbd5da7527ef1be052064acbca290944566ec64fbdd941902b1b3110407d17dffecbda6d1be28780eaba48f2b71e844c19fb454424;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h628ba4d17ccef12cedc8feed7b50d71276fc657263de49755a2304259cf8d6f84dc294221ef1393e45649c0528fbcfe06bc3037b04ed3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153475aa016bf7ecff7284d50498a8dbe270a0645d919b60afdc34be0c04ee61be166ac43f30c0be69761d0af6c217a482ee343842138d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h963471efaf06022ab79d34d2566814de251f20e269d75a456002afc5a1ebbbda842c91956a00e8a297cf8242a26066d2108095bed2af28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17eb9779c69f68f1140baf9ac206c8739ead9421bcfbb0c5be4ea12e7ee273c276ba47234cb2d0679faabe7743ca52cd75880d4814538c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156d06402bb4689d1afbe7d0d9f7113337d14ddcdd86ee6254cc2ef4224d3ba1867095d43f7e43bd01f6338c9ac1e84f9e9204163db0e4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6458d9a4ec958b669b85c63d5fbd7a2fc835361bfeefea6d12011872d49019872e03e9c221dbc8ab3771b43531ecf43df6a1617148eb4f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116a13157df3ebb954cd7e866d46c870336cea0e25e90a88fbc919b2c801598361dce7579673ac2c4698fc628d9ea44d57f71f795343b98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1657b1577500470588672b8c5547ecb49b24dae7c3b6f78ca58ef5697e91382c6c89611beadf077def3488a53175054e5d919be3624dcc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f15a12bb5ae440b9b79496069c0222669e4a59438ad25a1a5f25f17b5b01e43194c53955375bf034a195902de31a3791d9b9ab0da716f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4110298cbf603065f25c76ed53c339b924afc3f959b2a8748e9a006f094e3dcb79b69f5039f15ab642d0d76dc5974928084d7441fe5443;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e579d0e9e611689536c4f2b5038d2772c5299cb2a3d7d3ab9fc3b35951b80a1570b4a9fdc0fd99313124b23ef5a3ca0003bb943e59326;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha18308d00fdb2080916dfe0859feeb93a1f1527f4bb81ae0d9e1401f1495fbba13f39fccb2aee0e6b84202c1e1ddbfd0858465d2f4acdd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2125c1b1e1eb2c82e655768df3ecee94ada54add75bae0ed66fefa8ef96bf9aa1d06c4db30ebc204a5b534e65b1b8aeec699174dbbc1e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1256585221aa1db1a523a1c8029a2beb8325dcc18807fbe3894eed3acd2593c2008dafe54921b653c80d079344c10e56e1ddf1bce4f8b2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2767a78258aaaad763839c79cd30030900fdb94e518f3fdedea3e52ab1c8d892cea5111044bb04eecec944e8df3c6e2909d92ddbfffa6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a9dc30f3e4a5414cc511f3c0de387a72e2c2c449c70e9a366cf78612d13dfaf2ae83d17944cb56761e48ffe89eb83ecdcc964d886bb54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a05a11f2939cfc1e50966c54c497969d3df0caefa1b0e7ba28dfda5ee42f6d67993977656f94d48d95f8a9ee3033cba8347bf4aed316ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h969c4ba361e0525fbf46a023c2c4eef7cdd739bbd4ce9b337f25a23fec139716688efd9c85974402d9bacf99392940f9019d982148078c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c158cae3f1ec531b3a876375dc62caa454411f050cc2a36d88442b352c7156f7579cd580bbf2d3d3632b988e4475b9d626dda90db62d38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffcb8db3957c8eb646a9f9e52ffa5bac0a144be24361f59433237b739ac72ec1dc76407cf6bda6eb8ff9df631b9937d8acbcfe06f1a72d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b34c78c7deff6cab843ab4cd7adbcc955851b00fd5e915d61e0520c0b5d17e5eb7db131cf6eb033130be15674ce30f0f313b5b2e6a5e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcca7f1d48d4884d2feeac7b5fc6a85b59ffe9dcb5cf8106ab721c7efaeedcd2f71c79dda499085bdcc61fe3b9e4a929edc1b6ed0a8b6fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1b3bfe47a56f499f174d15a81eb5611bd6a9149ee099070417e479a2ea60695d4c94340b00c1f47cd3d24a8da56168e27877486f69131;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd8178ebd2a27e08b5326dc7304667e1858d0de394b32126e30189d9c18f3d1bd80b9c8af9b2da8450f6e82452ed3bc8cedf2ec4a4df05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17043be97b830a7431ce1f6fbc116024efca6983264cb7bbdd44f24d16eb26504948f66b680b89b66f48c197d98f26251b2e95efb8db3a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5745d011261c206b124a9fc44cff20e6b848a367f09058be9505b466d51cae832ef77d85d6acbe81b1fbbd8585afcf7e53f77f36dc5751;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14262d920c530251079103372cfbc45fc79af2e43ea74b60f71fc1f6183e15a19f99472397b0b07bd68a7cbd79df62a74e0934e3f3ae8ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14393f7d41e2d5ae2879f4411bf727da47f48eaea00c28a9a463bea6fe50c90dc94c2617a4b64a7b8d3640981dd8523ccc9af9a36921b6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf0eb788edfee8be8a395fb48711ee386f24df08b889adb542c6996256e44c2993e637e6a5cfeaef2d9b5900a45f1c6954f8193b7859c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff01874abf1f32c7256c62f7e51e2fbee21442c5d013c3646ec0a9e8a3946391867bdd9514e41945d9db35fc159de313be8964025d3976;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1852094ec8e2aee1243780d3ba40be8baed2cda723ef3efd5ae73ca0f85cb9a6c33e8d7c2f12a1168a15fd5f2d0d5577ac38eb9fec7045a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db575a23d42af735f392cd7f18c35a28a289de3b1d45897e93066f1356634d30beb4a962421cb964570ac9f4a87d610f40fb309791fd31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e5cb515c9da1fbfa6e9c2dce8a53158d0d9b7d8a95c3d0956641974c10c5df4bde44610b9e6a84290643e5ab114a85ab83c93784f3890;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4579513089b9e6ed7ff961cfdbc33c8a85204e2d346b60ddfc7542f06b86377f4097ed127ecfaa9ae58456a913e0bd0d3c75ae93dbacd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17af4ba9d3ca4227bd930f87cc0ef0b8511ee43ed7792d09d2b50d65a3af14aea95a299fd7664fbd685a0635ddf25c80f327ef756e4d455;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec83aa51960e189f207c62160eae9674204311b292778a882b7363f3ba467f9b66d80c8c18fbf4ca44183911d15155469c9a8fa93dfb60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd1b97e7e97ddad68a2f9c7e184d58cbe40bdaf89f7c7bb035ef376c403b75ccf60febe4496530b4d82c2ee915fea4dbaba5295d734fe1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7dae2755959b5b9ff3abba12e41e15645bab660ca3438fcac6d280598f917b133f36cf8db534ad230ce7ac2eecf4eaca2d4886fe3fe424;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1879a17ba09563db4b62137e4e5bed6e9e377a49ba40751c5af163f2f7386cf30167b3bdd576a47540ca2889aed14a05d2021f9d4faf377;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b8d75fe1700d0117b1e5ec1ff83208453669ace98e2715ddace26b4f5355f8948eb364f4437873534d5eac1f0fdcd078a40987ecced3d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152f672738e7f774a1bbf13459e313e144f65cfd489babd057cfeb7fce5dbe7f5acb6464afdededd8bb64a1c3687585dcbda66cc0037550;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168d89b6be920f00dc6b7e6f9e8db46d09dde7180b616d750501c9d7c4170963d85602affbdc70baab3dbd0d79f5d766aac396468a4c9cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e3b4ce7b3679513247cfebfd31745df57fd349cc0b7adf21644bb23ee1e9eeb53dcd227d57bcc2ec1271233d2a6e69c1c1784388c0461;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16bbd3a483eebafcd01df256d5ff510c9bffd4b1093dd7c3e595b85855c271da0c19dd96b24dd0174e5a77d138e33cf1b3da1f5bd1d85a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181c751ceb72e155a790e2ab903c3786aa3788385028f41430be295ff43beaf7b7083f67afd05f981f947ae1e429cc24e60acc55a7ae8b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h160aed30468a2b7b7dfaeeb9c72e060f5b0a7325d798d7e0fd5cefc48a4a0d53f1e27b034b53ef00170ec366dd8de351c3c67d8a4bb6555;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h466ec94d2e107c471e2af0326d8c461e0570e327fd6ac8460f9e76127aeefdc76b1f83fc7f02b5f7831ec0ba9d543358d4b4be5f3202ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91293b7bcba767011cd111a35fe2f3d87cae5db5e3f63a9aec272dc5747e48b9401b8393c2dcbc291bc205de23596679a9f0388b8f059a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5ff327a8ed62aa609cb81fd1cccf1bd92ff5f31b89e5c54b911c2fe3a2d3ed9bd8aba646b1ac52003e6299926a2307ff3ec2471a87ded;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h944b15fbabe0d6d0054793b2afc302ddc39a7afad680af26f2de6b860b00038412f9e939c42fb021769fb26bc8b5fcaf762951a52dda4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0a3e1223e958b9f4b343a51fcad6372d527ec3340e26cdaa14dca0b56efe9fb12852c92e17db9d29eb0393b525a3fb8b3ff8bb68a3948;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127f42537f4ee47d050bccacc8ba125906ee03d47bbae2d5305fe5d0ffd63302efac8f74fe4448dfd1913721b12601ac98c3454209cfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5426c80473458a780f961985feb28ec0bc659174ce0bdc875b0c51c2abb1eb236bbf25745355a052e308633f12889cfb94c23c4391de4e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd7a8d495e4ab7300193eb966ca28037b5cc3fccb4ab151823f7924e88c4ddcb6e67d88fd0f3111b9922706f0273ca1fcf109cd4688a3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0abba4a9633e1eb79a7f76fa9e9529fa5ff5e06fb06b04a18ea03e50de92be25905de673d00400b994f9880c16b39b3619952d09362a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f9691e3f31535b75d9b1f4308f2fc792b73ad54801e7ad61f8144aa413f63bef32b1ba092f02c2566f3341b6c71035f76c61215b2cff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123abb4808c18361e7d40415fa4ea4c39f841fba631280a749b84486081315b75fb965d6bb3c4d4bd8dd9955224f0f0946276b338ffbb54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f30e5df4a313979382210baffe5079eb8e00ac703f615f1c63db72b0671b50c298771a193fc50d9d639983ee163a1f48decc0b42761e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9fd43c1b508cf47e4a2e0eb213ccfb7a85d35916c6fce38b1375fb885d413753607ef156272d9a0e3fb5963945c7de73542755f316973;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14105dcf16564840c168f527c97d0032ce7ddb8004bccd5400c1f75889b9af4ca4d33710dee72891104c156e52d51bf44731dadcd7339b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f08a3f2b3c98140d1bd0db65bf91565f4df3d32454fecda9185240ddb9aa68e686f40157a68f806c5e1266a618374cc80fcea50ef12ee2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b684435bd0026eefd5e7cce020f175cef5c29ab62ef715e8a37c74e591059d8655dae3081204b0c0271f348c5a02cc04fd58cb7da1ae77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3760dc945aaa5ca1f6e9dea6491d35864ba36c85a3833d976624ae170e5b0a5206c83c330c426f468e5ee6ef6e30846e9ed2d96b80f8a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128e8e64c2b0586c3c6ce1f566aa0ab05de81c258c6d6bca2e6165d26f148da51ac30d99d43cd947099b48a9776b3b0b183eb46c307240;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35f2d3cdc75dad21a44fbb89159686de1b5ec35ac8032d5a9c0114209f800c9d7cfd6470d712589def311e32b010bdfc3fdb41bd6a2777;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ec84b868e8718a66b29ec6aae056bdbd4e69de1a4efea6963c5398d84474fba318eb7240b3cfab8c84286fe58d634a40cbe863175887a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193b550082d56709db4f1284f08e9d1ec15cb1090b836e7b6c168aa9afeaae406746860b361845b7b2ae343ecc54705a84a7d3b04e799c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ce6b8b06fffb5c80bd12bbfebed1279002913f7ba0c46b8a21565059720343e3cfcf2ee0d71ba305272cb9d7e1379d82a95c293699b31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b689fd64a030fd760370646c27a9c0579f739a38e59d6380f26e68f2456a2e38deadaa784a7c9a1820f30f1ff53318ff4452c9bcdba2c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11efe5e9f3b1104a4612970319f259c829f6bd3eddbafc49d41d5e37a991a09e43fc672eb8ee3877c68145e16a0313b8047d2f4f907a2cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5c18b2e2fd11b663ebf6bff1232f19e6953a2f32e24e7ec37f592910ea5e586fd2db507b403d550fb91518e0b1c3325fa294c19a2ce0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8b7289581f64a845e8d438343d95e10f3f38f506f91c93ec8a8200e74f2b8ed07acff844b009de6fac7c5f416989aa140c0f1d713af3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107d7a0aed0770a23dbdd684c606a465eec9ffcddde5d07ae7c0ae9455468af76912e78905d523b3cb9719de6fbd0448a1ce404eae1e859;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ed80fe93b04ff6cd211b3f3cd579f440b8dd4349cde9f199904e7ee079108a85f971ab29f39f23fa5b05effd3fe2fe20b83869a83528a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h983d203a41b9b3bf411277a7d50bedbcdbd8ddb22a6b5ab7ba21e0d3ad1a330414c83743a41d26dba58ac692c64b9893bfca056e7f1420;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha07258f5685d9a6ba769415e09bb87d57876f4b12963063e3e499d8daf8780b39ce411ace91fafe4ac736a787cc9c19c88b095f3b96afc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb8730161b82b8b32456a68e414e0b56651be6e50819d65129869bd436eff4d2d9c5fbe5bec7bbc9c4a687167d5c63d62fb5ebb5735c57;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d43144603d0ddfb879f6f17261fb410e86ddc16b476c308736d605ff93d1b16b19d160dde3ba1534c11ae5a87f3374177476d6bff27490;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3baf0776c0a6a797bbdb060e779874e5ae11b057d527193e33a41f9ab95eb492114f50123a089c929a9b405bd7a3f9a75452fb1b72b6ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc88619fc2b4834a28d73b407f6eb62db514597667cc12143f61d4acc171610d9da741e9058cb12f16b4a4ab849ad46b697a882ca208a11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce8c2159f78102144c7c855504561b870a0de83b1d808a59a3bbb4887803cd0e1468e4ab270419474cab275bc833a800e0ae3840b69960;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa3230e08461b5352a34a11d5597ddd29e9be59303cf1caada51ab703ba9d1e1ffb03cafeff4be7e5c3665cd95fd634fe9ae363016cdf0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be3d8786122c56b5e664308f8c048d14aaea74f6e8ff38c62e07098a11b0008451c4c230f30f836fc625872aec220a1e9cb571dfd74c13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8184d193ab658f8327c6a411a34436a2c4e3b1a5bc016f650030e6ff2809d828aa49079df38b45a2eea3965c71b429d0c2b5baf6aea863;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ce47c20f58a31d752efeeac04af247dac5a4b600ecee15ba15a350ce6f5adc752b2e826c80456222612b96deaa8843c8d9cd13a8b6df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c48fb4ada2cf60690f8373d63a04ec6f000dda61b0927266d36177675209d5da52b8b7fc2f9d0fcd114140ed07e7d43439875c55d68fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186174cd218558d964eb344526bb6d2176bf4fbccfbc53b83f24cccd2814820905cebf22a5afd00e78a20b53766aae58e12b2630ce678fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102132c925e793c730ed7516bd149fdb62ce5aabe0e52eee72a80b51118905276cf5f1c2ac5de639fa5f4122df53f74165bc15d5f4fc861;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd3a36ec5fe7434050ff86a3dec55ef4f59fedee45cfc21eb92814b594e0776e9748e3c5269c915f939c0ed4f4f93ffa93b2c283b033ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h143100958d2b2dbf74de91ee87c3e15afce421f2d17041f6c4437ae90cdf44b11548df1cc1cc2fb9a2a1562f2b6cd56e56fd6a642121e26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8a85a04a4928cb88e73b554195a65bcdd378f0ee6c5ed02cba46b727e55250898824e26daecb390a0eb54f5397d40dfeacfef0bec2563;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af876e837f20bbac8d243a3288edc20905b1b23d179fde3b14db1578f59b2aaf7e595ab57baa156045f74026b480168fe9758d4d2a190c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85b3cf0072db2fdf2b0853614cfba38feb616a1825ef1bb7ccc85d0732009b48c6a2bf2a5a4be740b515315eab47a13299661f83e67f0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3d721713c7e892e6a29fce33ab741a4599bb59a347017da9b08a5c5f646017bb5bdcecda11caef4372f0bd7521db6646b9cc870fd8d86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125c4511f2e7f0c3cabb345ac4d30d81e077fb6f2e32b6ddb2b19198c31a1161ffaa0a229fe9f05acd1a7b1f40f155e80f1f26e9d543899;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hace14d67d02019c1245afc314687497ee3aa56c482c57fc5c73d50416a0be411daa511a82c69c661934392977aea1c636b085a4de62c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d423da23dc302225b81f3cf723bdb1817edb5aebd5c789392091d0459475fea149cff13cf476ec370b6c608297843584781a6fe00c632c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99cb7e66ec5dc1e87bb19deed7ac589901c755d6664cceef4e34a6b7cf274db9be6252bd2bce2155ba790962c1ef7309185b69058acc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a631fe60d2fd49591ebba0c41b6c401180e66de86eac89e1d63e21119f4755c5ab382436f1b22a2d6122e620f20767a1c0fb5dd9f82d78;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcb30f48378ad935ef7d14905f75ed8d7ae2f4887e1dc5312fde17d744886c7e97af265d186ef7f2deef0e070fbfbb26e64572edc19cab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149375794098bef7b32c15c3f7a80311da447dd8ee3ed2c29d3c640af9afe5ec89c3aabccf1c66b77826630a6b9c13c6bba702202a8cc6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf990e13e6eb14938ab9aa4ff2318e67a7c3c2eb9762fad258af9d96cf7dd24ade7f08a94cb0c890ea0f101f09df6580608b2c725e320a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7f4025559ea051d19f2b443b59bdd67c9fdeae6e7cd9a80413a30350762887a6a37e2d39b847ab455f5a2b719d1a8b4be0f724e786dd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1072cda6a6ae5c671e812f9fa0713e917699fd8fd7e21a14861965821df85e7646a788dd21977a895e6d2f1a1ec69b327a4eb60914c9484;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf361ec3bb281acd55b909c6d62352174ec6b2f9e82e1e1ba316a988599ff7d580e3f58fd823534359111e0944f30af21205827cdb4dd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1237f3406d266753fb21dcf8bc5c9c5358b568d0594051610d4a8bc235e8167ee7a107efd6feb581a61a4839e6a9f2a015012f10283fb9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c2872e2533bbc8375f27b854a5d69266018896d6aedc962536b74c6a5c6c5f166017320920d16df24be78a547dbb396c591825669b406;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17df132c126ffc43fa78a6d5dd45303a211e6ad88edd591420eff9e540f91aa0186bc1fd9edc7e04696c664c4fc02de521e82d6b97f13d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4e64b8edd7f24bf6e44120db0f00ce3d2ca9ffdbcd15f4b0200d4397782c5efa05cb555633cbb73102b783e02c1a900abdc604e6aa75b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1010ff26d895bccf910bd3fd81c90527ac9540aa1e9cbd204576b4ca912d445125ee3257b339940a7f67736a84c96e047921120717547bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1710229a67ae9401750dd5590d2b19fdcf56b505519aec1f92c6033c86ae432a57a7b4c15c0e7b766c771b0e36b016724be788b244d136b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103087047477348c5e2ff31885312e93e58a63ba142e37964e275c74a322460197cbcbd0255241c7d39910de1a2470d35c2a82e880bedc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca420d1e229cdd842422afd55bcae0619404038f4d7945e61a4eeff66703b85c7378b9ab3a3da7203a8d251d10b93badb8d2564ead06b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3500e7082b5025cb954965da4b748616e9992b350a2eee37e93bc94a2795a28d5070481c3dd6ab743181b5f2236bd1d14b5e684d88ee08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c807309fd56613cc7e4377b4815d6f8fc3320b5818bccb93d5b25da74d8c127cd62a5685ed7e6e2c996c1275fbbf7b82466a302fada9fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h381f9fc8a385c6b74c868100512887d40dec266c6bcb31e2a1bb89df0e7063a655560fa1465dcc500b013de1abeacd62a9557dc3103e2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1950b57134704d1db399702fd5ab37402befa2b2d82d6d9b5ee75f5a33d30c2d30c2f3ebc26ace5a7b00543ded49ee0ee85b84bfe3f26a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ad2be8e239c89cb16a9378f99c3c816f06064eb15d9d8248681dcbb92bcc1238ab1cef72e834c737c6dbc4cedef2903ad05f2d4087bd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb0d18b4635c871b7997dfc6c1404d29a177d39bfd690891ed64e3d44ca6fb8c7a96819cc4d0e0e77d3ff7cd8c3fd54939d97375bcd38e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef3139d1450557bb32512d2704c329c084324ee0f8e591f7cf1a0cf27811ea93f71db27f4c581fd4929de78c1e20e082204c3ba7b3ca14;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c9eccd2f843f8807c145022aa2343cbcb8dd562e8f6355c185491e3bab643f2634ad7ad5a91a144b1f7d3079bdd4a0d09a1f0a68808d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h320d0bae15f24ff6a846b9a8a3d0d08ba3c2b6d6e887950f6621cc77efbf418885dd37921d8af68d3ba19560313f2072554d107336eca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18562dde068a4e579ba52c037b917cb9e1f068838915deec58aacc5b1c7ee1eb68e354da842c0d299fc804a61605ae83d8c8824857ee29f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8d038fe84f28f767364eb3e009457de49907b188a5d12f4de2cc33af4c3aa4ad67e3578327badbca124fb223eb72e7fc822149a649e7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd091bbaf48e2a8e53d365364b17f51dbfb854af25f3f51eade37c6d3e09cd50f14226c7eca6120e399410ab0889e7c8c0a13bf78a0cae6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1221fa42778f5bd6a7e45dffcc6f5f8051c962e11237fb4ef18183b3fff5401992f0d867a9fd28777dbc760817cf8900683fe62ce5cbfd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138ff055d4b3a36a7d2e2eeecf3525a88f282e7c7df79fc14419530b7fdc67d6b9b585434b636bac058a4d769c71e81a64055680028d55b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82a79b03a5d7ed4bb48008babd7c03c5e2284df0a2a92b404be6b50d4de2354921534bdb9a9b5d545904f5f26426e0fc02412fc2d0a141;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h979ff8477c026e62af8b071f79b7a2b082b3a5e42704dc02cf9298c1289502de0e119bb6a7e11511a2d1744b708f7b11ed6c47851a5edc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2d897764a96529fa87843ef10bc2d4a2c2c343993e7d1618e39e906b7e824fa094fad4a7f03334187a40f00be6124006cd87c1f5c5c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e63ad30febcacffa4df8e272601ecb901d2cf098a6c9b7237993ab6f60d08323cace0164bb779d273da4b76dc40f9c9e98cb8825f5a180;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10dfae972870de6f7d89aa406162e6fa7e1e8649650b4b50d32ff2d78943a08e59021b3a0077d184a40e7ee5e3d53e4a4fb4a41977f50a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h711672212d7cbe5090237f650d4afdb4078f5a6fdc5a099ae21681af0fada1725d7c4ec9a17ab1f5b6ce065d52b0470e8c661451441f34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6393deda66785b9cf754f8eb2d5f1810bd01a143ccc407313c16a976ac5ba75577d028bae3d106bb74625c45fa34b33684dc5fa4101937;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c20ae67599b4eb0737d383f5a53c2fc81795911ab295c9f155068be4179efc511c9af14afe444f23e9825f01b35a9e4a5024c72f2cb500;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191f4f61007957e4b5a24589b54f5acdd7f4c20a7bc15373f41fcf5dc3346bccf8cedcc529db5b7c0130ed1786f68c4b311d55a9329316;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182845554880bd30de468aa8d2ca32b8c95894ee688c3adea6e05650f0e78fe624719e7fd31018f5298eea3f11d4bac2a65391cb5023c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111bfc579f3e8e7f5fde972f9f2261004e0b6e9a8aef9f386be84f9d7f151fafcef84a54e7f36762037c202dd6197c98b6ea5c9ab88457d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86032eb13d0aedd92a875a814008182e333d2b209a04196de457b6445c87cf5d4898dccbee32bd92d2a048fdb37c3b1311406955c5023e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h313eea81c4595fc3e0eb7d35259d7751ebf5a2dd1a421fa084570d08e0cc2068fd964beb17d925e88c03d578284a6384dc4911eca4bdd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87e64aa61828c50b9b180dd3c488e19094fa813ecd24e1876c66292b7b91b0fc812e0240e107e8fc3004e0166ef50b2ecbc8296052579b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8f707c80f6ba845cb7d8b339dada9ed1257be1314c501dcd9921d0bfedfcb23bf0c7b8ee2f47a7a1255193f22e3adc7bf612f42833b85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18dbdf6fd6ea6d81c4e7ed172fa186a3a26ce248ff32b71ae67c0ccf0a145a4dd8f04226ab583b5de3d4642e2ab05479f23c0edccb5c08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bce1a68b24d2e5c640aaa8b0144c334c078317cabfbbaedaa5c385f447964711d3ec32c9b60adf0ebc14a058d5c0d969efae82c02dc782;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3decf8ef6ff9e386aeeeb56736b9b8ea57c10634e48d1bd9d181379576a65c576dd28278d4531ef734096dcfa8c26e18a419550485011;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9b206f2ef11c849d0c1aa9258f0f7e55159fbb7538bf2fbfe2436082e89f82ccf5d8b0ce48793f7a4de56d1e191e2025c4de3bc8ce688;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198d96ee993f6bed1317e0676a73fbeb82dfaf5e1e32a3163419b5706af70a0f7c85f2a6893b2a1bad1de8da082af99481326326fa791be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h205c207f32f9774e79bced751450ae766852919acd60cfd986d65210d5b609e40c1ad4f6a04c651321c2de58db1d237caa4fe5af042473;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39bf6e4ded4279656bf686a43556c097b9e643ef12ce279359b5b41658d94051ee44be53e98ad135c64dafcfca2f4ceba8dc61589d6247;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haea533e19642be9d10a1b14fd469bc42857aa0fcd884a047c0eeb3a44cb7e90f1d8da139fb7e09df892912edc779bd8be02c68c5a7d12f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee58624cdfbed9851ac71fda84dfe8b26d9f38cf5dad2ab9c8359dfaeea35220d84e0b14b6c44b6023fff6fe46b07d3ff1ded751badbae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140034572066ae2656ae80ff103c812fed3f2ecf69585d8862ff4fc799026f8e859551d614b2ae5e4ac3e42d80b868bc0bbacaa776ef644;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc36ca34ae7de98906af14843a97cfae48214cc955c6c65e0d8528adce76de5e51f9c46447c50e7aa4aca1ccf0ee83407a3c1ac6e725b6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eecfdc196bf968f22fd61ebaaf062e2190f975aac04af806374d0c973c003e81035a7690e5c0fe2250c357557aaf885e37ad469c1696a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e918c0b1843046c7cceb59c06743879258f37501e6e5408f365b6d664fe0960ff0e834aa92b19dbfa93e5c4993e8d6b14409406b53a66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155c51c811a227e300f266ab6e2a4a4cd4241c2e9f6a3839262b664320d279d46ee4586aa9676512e39b6d4e28e4c8111789ffe53d46a4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b116d62a65eefbf2dc9d6b073cbec5da74e9d7a8de4d3d7e5758decdc5af2d6070a8fe691d1e6c3c7836ba79a3fcb84c03b3edfb573576;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9031f96e6aa1a4d43e11b808f2ad1bfe4b042610b55a60367f23eaea11c24ce143c6b9a16b753292f1ed006003ccde1ad275fef39256b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81926efedde530e255bf3bfb9207b292dd6014da8ab66daa66fa3f9ae7aaf2cda5711a9a5b25681412fd79c0613d2258ebef1b957a27c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3792152800d69879ad62b718ace77b5d9fa1aacec0f93ac495a21a0b2e27fa772f7cd428a90ae67c4f64afa9ca5da967ae33dcf47d874;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e790484ba8eb4cb1a22136aeb9a2f48b74c7928bd05c3a4a1d0e77132b693fccbf0f308dc947e00e1740aa9a28a4fe9716dd803a47664;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd436f232559a6dc52b2afc2d033c886dfb66fb8d948cece7b6c2a7e428910c814d37471a3879000ea267ac1e7df0e6d102112f7a89df1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a5358e3d97a2beb744dcd19e725a608726678c1dcb01476b5a9fadeadd64ae54ad444ec2638a848b02b3717e52773a038a8e510ae8ef8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec7fe1471a0feccbeb94331e2c0d296252c33bea359b628b71054c2beceff7e7eaacded1c061cde06281c182ff328821c0f8c7d36c7430;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0cdb4db0142174a50be2f3fc136d1ecc5c05029dc389f083037190a254b308db5b38de70d68137affb0a18c06df903d1073cb2b81ec73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34a56f4daf961111be38b482552c138cd5432b203e23e71ab2dc55275b89c8946f2d31a4965d11a71a6ff42b4b932592d158a0eeeb83af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4dcfb8f11038bd9b5dfa8ad5079887dc0cb1296e6f1088fd24b0c2375cbcafbd95266d27c36358f9b49b8930bb4c70e5fc17a0a4c0019;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h741cf0150ff275bda8511109d3be323fc10f8f79e228a2d92a084099a8a5c8ada0e1ff1f227ce3b398dab77a6c5c5560f366d7b875855c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a65c2ab4a7fe830d13323c632dc9aee36df9abd2aadfe7ebe5b5859389f16c4bbcf70c2f493f0f7d0c8258b2cf61dc2ef94eb1e55cc447;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee666d8c8eb713295fdfc3c4379d246d318245c89e872fe578b26cc3f77c5de92ad46dbf3995ea3f461f0c9d553e061e5c81977e8bc1be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c13ce9307e565720f9ab6d376d42f21de587b2fec3231096ca64b2f726ad5bf9ef33f5743fb0977ce16a24abe4dfea9fca8992e91431;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcddd09049cf2ce60379aa442292499d8d26d4ff39bf0d1877427dfedce099140c3d8e146afbee9d4bba76e88e9af62f86b8387121827;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f9bc41ca4aa2724261b607673cb6179fa30833bbf5621154ea8e0b623da4cd0151e93c67baa8df3a47137b373db88cd55f063f0a99fca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a0631500321c2b432e39613340ac619e4431951a06730ec9936c53c09d81721bb13c9e4e6041d37ab7f7fb8d3ce178bbf644338685bdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c9610e7b847e673abc212df59875178b3f26847e6ccbd0502293029c37aa303c472e36f3eb082dec2c3af25f636f05ec02fd72370ebc6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h777549c03e13563731afd1431b8a4a9af6dbd25ca1b068703b9a9c1419d0dff48bc21439af54fb5ccafd3b9d031b7cc36047f6a3849733;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a3fbcd0c19d32c9cc02d4b15c16d3f4c2080a27c5f84c1aad1e1bf37415ce1637b6c7019c4de34086a3322133153d2402fee8b96c13c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h807f43b6e18eb1b4c016505d1449eabb490fcbc7cab6a3ea6d183feb75c9c916c923edf46f7e2146e031d205c1e8280039aeb188131eb8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c20e27982765b293add783e5341adb7f5a4abe97d908bc6ea5b6407ea85cf65b2c2a2d61eff40a5a09fb42ad4072abef77170e8359e79f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc2a28e0537be7ffa49f570253baa582c6b95d4350e7d891f1dcaf53f39b1ac4cbbdd14ec68f217801d1b1452009b22069685fc4f44d51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0d3b1620593836e1c1f8c60f2041b23bb0420ba547d84da32326e05dbb0074c9ada9a021457428ed545dc480575eab75764e9ee96028e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc25070dd18844f5a02e2bf17f70d494d1f0426341f4a0a1d0fc4ec5e9acb7d11e4c7efd93e4574cd41da594e8a77086e89397da2de767f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199853a2d20571305b1eb5850e12d1c25123bbfcc6559b7bda45a4bcbfa8d073a63e41fd4cb0b9b4839745e9adf9169a0e3df071c2f2e3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h970d1c24bca4a34e14a3ce6f3416f0571f77e8d2b6a9f8e63256b553a7731de83c7cfc295ffe75d0762938e2589588861fa9f15b5e8cf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b82fec53eaff1a64b87863b40f5c3c4a7887485ed8870712edf25a745207e79a2d4463d4b33412d4c4dbd16b7bdaf1344ca2c49988d73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cc0121137830eaaa1c5c2326299e0bd0fdb590283ed6bc641ecb8b8649a31449df75c96a7711b028549f058e2ad7ea63c1a280feea8ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e82a949db249e1d0fa4dbea3166d3a597fde0fed705a9b61a03508d726e613189f504dcf2196ab1e4821c0b00357352693ac55539fdf7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1589637bde664b6171a7f02b7bf5ceb367080e62dbbefad814a56503a4e6804e235d3fb92b148e5603923a2148d4e12068655cd8cf13c66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd326e3123209c6e965a3d764630ab52de65be8975d4fb13b9fed197a9cc82c0547535a381d51b305f4b6287c3b5997447d294c87c4f8cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c4a67f2d6a923dea6a95345b69f090b872ec0a5daf102b0980dcce49d1ea2233d2e776290288393a92a9de69fd85ba1a1305f5b5dac27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d4f6444605fc04c0d0274431ec3187c4b9bf8161b6f2854b1273ed6e40259ca03094e0ff85c40a7656bae686f4387a2cdfdb634ea4485;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e961f5c7bf9113ca754fd909ee9faa428c01beb8304a8fcf1b8c6b94e02a1480a73839019d84e2929c7421d20b08f5729fec3b4c4d1783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103a7d9ac699e2c5b4e1901fb4e182f2e5ecda33c53c1ef1e6008619a1c4c9f353d60a53915906ad53af61d38ac5d83d4492872f68473f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98de35cf94ba7244ca6d6d7c4ec6719b7f846eb92d795c61f65270ad3c75b4e3787f69114e4bcb19b834578699e7616f4f86d27ad4d19c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a01bbc9b1c9e86b7e3d5ff8ea4646b2e0f27e6a8ee439264212c2a486f3305bba05895d8b849af51e1fce90e9e3682721a4a6252e2a97e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4b3ed360f2fcc9fa924f792d16315a0fef5190573bea8b6f784ee334cd5572d7f325709cc8ca6aee93ce778fc9b1c31d9665b80248800;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1db5cfee19c7e612c3e04bed77fcaf4b182dec1da4e5517e4a235293ec50ba5bfa8db408699e2909a98805bd603ffdc6031374b497852;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fdfa8f46236ca6d14dc00fa9e99adcc4b64aad668918b081ca1c4d6b628b9d0bb1131750ece7dc06916a96110a486c646ae2deaacb7dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h412ac652a2153fb4acca48e9934f86f5d34d11fa8d3e756b4110327ada9ce11a91c3fa264557e793c787838a0cd03212329ccbb3ed2ac9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacb69d9168a91f5a80f0822eb02fe0ebbad1812a246cf541b4f63986ae7a76e870cbdf15e38dcd7785b3501f595c814379e1037b15ef89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141d7dc3be1daca32b8821cc94898caf2d76d0a38fb4094839bda1f3785a7e6f793f6502935ed3baf7b2906321805817cca4f7e9d0455c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87900f460cd333db88238202712f2afe06b3c55de5bea65ca1c15cbf4ca618396cedef79c65a5d664fb8b183858f42f28cd253352a41b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe6766fb2a49ada5889165d8c7f582668367ee837ce3f8833e792b5918880bea44644b16cd2c7c386b08e8078c05a4eb6e42656e0e7a52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166e3429a4b6eb1f66219403805fb23c0815604544c1d9d1b34d592ac07b8f37a6186813ce2ceaaf8f45c0c2af95959b100ee154183e724;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6b8641a933c478a0f6688b8186a0741abb4bb491d45efb9755687c98f5b0b716778ceffa31f88bb0f12f84bf5e4cc468e9bd2138e202d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53c6fea8e2eab47b4946fe99be1fb01acb06c8db8e0a254cbaf7e1db84676f58dbc6a039fb9657a3c0c27df11cd78818e8eee809120311;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab8fafa0fb081c6ebf19a8fcf995261c336a7bf2013b042b39cfc48f0cdc9d73afb869970f9686fe9459c50d4b68048331dd2bd25391a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h737c031422375f75c521e994d15c8ef7ac419062beda1578e3d7f87e6414e9950d908b42c9048a7f8697b5f16d4b558d45e3d2c5dc527a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c7bfb0f33e59dde637add9e2a4b059419f47aaae368d76ae96aa75baffee0e422c3ae61a82746f5088afb83244d413503b8ea5c8159d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h359e0410d67af608c5935fe1f5db278c224009bae29cd521395708d15f4918006f26fce17a7cc5fdcaa6b2a053a27feb637266129ba08f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fb9648db036c87cb5e2e96d96b77538d037537966ccb0cf5f08a9824b38fc79f36bf385b97e38ffc1a727629fe1d7aa6cf51cc810fb28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193d5ce3b3176d683a15b14f0609ffb67bb1918e451b7857b0e2cae085712812981920645331af3836cd29e83d72b397ce4526b8d323015;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a769fc991e1fae2916c06794bbb4875da7d38913b2ac5f0c45387e1956c1766476d6f9e7e65199b40822d6d41bdb0e1d0f355213d899c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18328218be7129d90eb629af47733c1937720bdd2aa8095559eea4a714b9650cebe692986962024b8fd35bf6f0c59ceb6f677886bd9caf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac4b5111c1898c3b55cf7a718839a39adf6fe264bca39ce366d8ad571d295e2bf5a19b52b68d675559481cb330608f4b2b760302268817;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fae835899b6d96a578a059482120ef76a1cfbfb75c20a4fe9738674b296d024a4a5a12053f8cc2e0bb77c298d84f1b6ebf7ccddcadbd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f52fc433d0599c61022eada99b57ac89d103ebbbc523de969f9b621911a733dc784ff1e9f1d49ff94338c9ea531a714f935600e6df700f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bda7a6ab0ed9b9e0995e563a263444fc75b9f71e010ab1be812bf76dc988ca9805ebeafd537d50c927e9416a51727f7efde9d036266191;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d92f7d6f74bf23073e10f8fafff4a134ea060477519c976b6907be5ffec2930152295b4270969e38df02de8394439de37f68e9e103e91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8b969b578fe1a80a4978b81accd832a36b884d5ad9962ca6a06fa8b193b73ddc3127cf8e237dbeabbe1a98259731fa62587cd03381460;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8bd5de69e881a5c896bf0d156ba47bc1c522af498a4c6844b47c5fc16e6b34009a5fa41fef75b3fb7566c7655dce8e4de8cee82617aa0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9f6918f4c99102667358741c5a8b9ad0b44c4893b0d837b9ba5debeb0b0b362cc20af32ee2a305b17a1997aef742f7bb851d6c379f96f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c9243d772e713fb70cab395e64e77c779fe2e040769aa968a35120f973deba812efe8ec47bd6c765a51a928663cc5771937d940cc95ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd428a1c986ee68f8ac2d9dd78ebc1964d81d5d69bd0510f56cdce164b41dc9f1d659860f7b131efe760d207c244bf265fff9787f4a0a90;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ead6cfa8c563f9dc7466de5018fea260bd37a77abb33af694974bf3e840a8d5ec6f445017420128f80214b15bf9417ff5240144507b5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190a55aa4f9df6a92074680299982802795770bc138ae8400e8eb90580bfecfedadef390ce7354050f6b3b18f3b00af9503d369ad635d08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1577aa6782b513fb21d62fab49035e8a1c44f374321ec0fdbdc0d01db145887a7de876ee9618a86fa4d92b096fc28e1fc3e26a29922945e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h318b63ab3cca63172a2818b810c1893a95ff99d322e1b2bed13f3d65c3d28b3c7752736c9865f65fc10ac134354f5343e24d4deaac8558;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7fd6f6e49cd96725f09ff7a72c76c48bf9878a29f2b93eba00d6899b19333eb684782e7a33887ed2a26d16c4ece2b210db99539bf99c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181882882b4904bc44899ef8db031bd99540e8de7ac19b3d17573dacaa574939061b59d8d8ec136b2faa18fe68caf2c0c47d2d1c127de7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e8d51b59b65689d92750217c195f8ddc2484478985440ddf55b2520a79ae73f1f24150407eb2f02de5560921935a1dba2a8b6bd053034;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156336b8cd14dba10e249f3455cc0b19aded2aa84ce91151d4e13508118c5612cd0af19759bc58c3c47749c89a350ddb8eaa372408b8e39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52eb5520d173f2a34a64f8fe9f5a7e8acc09195cbb4715879c61e1608cc3b785280039e234be1fa9f4d9639fd20a6b7a21e3be4c1bbc17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf41be7c961f45a2914bb7397b003b683d19ffeca344408756c5f7d6bf7a73e78cfb0b918a0c2f13c25b13a1b92210d008a44bf87c073ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he64c7658984dda91866bb9deacc25523df9e950bdaefe1f6ce1fad91596509a4991866692eeec9161a9118e892c3522434f966a7b6d5bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae0d123f409b37d995533dc5b2232a41ee4cbf02b9d5974a741326cc47924d9f9b63e4302a8ffdbfe03cea65776656b4bd04524832f9f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122cc5ea2c6bc9b7972fcf8d6345fd670d08bdd5e2f5ff6bc01ae759a0b3d8a110ba5dffbcd6ac282b10f17cc05b36a0f020b21eb0ea296;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9febffed9810d3a4184f3b4145e21ee415c4dce65661f37204202dae055140792c5226d29317ecbf8bfb72a5bee1c34f57f44a03ffd58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1588fa231a93a1a5597f3fc1986eab835ba030890a619bf97b326bfeb91e5ed3b64c6017346fc77adf021871842f1bfbdbe0f77dc615163;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be4ebbff302c45461ffbc381c88628bb7f2044ad958940f8c060c38648074b21fcecd5aad9675680ca3d2678060188e201ef2e7eef7020;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf545aee1235681f371ffbfe09a75b033529de3ef9579d9e078ab3d7f40ad1ca2df62d3c88b524479ff25677974e4c087252275f93e100b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8bb040829f614dc8857a49e401783b105cf488401c5515eaf5a9b2e9d1f90e42a2af86687bc9c2c4ed4db02c14fde6994fda4fcc47994c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc3348ef1c5c53556bea1d1a360d7f4ca0f703a7a721acdd38a9b79e008e718de1ff3382647fca979900db275e904d77cf7900bc6160b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7001e65d27866f89b4362138bf0319908803e73ca5bddf93b786422da380c05e2acc4f82426f71d4dc9e3b8b014480534315a737196869;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ced2ec0204edbe765aa937e0edee7c1af16c4b6c757a2bf8bad4e2486e988e599c872ddd7cfe59a72b042c0992bb7707e8cf64dc44cc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58cb9abfc7752a7a94a82795049f07ee9b51303fa0e78d0dec0935ef9fe01f437959aa51dc5bc10c3371118f1146c3f67890cad1bdfad9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48d13308ffb7d4e69023e1b7c1b254362e1def58ea2353d32bf64297b2caee76f9afd91ad092ed59cf0deff40e8e9702c75f1df0f92bb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h652a7e0464845ba42bb2f80bb4094e9019405904972578e1f1f7905e8fe9b1a9ed1bbca3444c23e57970cdc0afbff6a6b9c85806edf7a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa74f4ce5ffb64b269c22c2a72cf060c0dc5b71d9e727ee24a504eec4ee46f3454a9930c425773c9e186fe44122e49fd0285d2ae8b8297;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdee7bdfc818d947ed5526b7d35ed99b3557d1157b86f673049f84ce627a62a3135e5dfb06c221dd52f5efda3e3fb3f9ad4810b929d0d86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b6160aaa86f79b957b3db33cb65e775116d4060f6bc4e1ecd65a1edcc0d55e78605d85f4671b34c3c84340efeeabd23c2a8a7de901ba2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1056338542b759ff4e2aa77be14958822c7c5c96545e99f643e6fae8e8f5ce10dec92fcc115c9deaadc82d46e2e8d4f82232bf7c2790f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfc0dd5663c6e9bbc5fd83ea9cf653edb636c22efe0c27baf17f24f9d3acd7d08991cdee62004b883faee646637335c9828ec0cb974264;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7ddc6484acf5a3156bc0ab4eb861fb625f41b655dc808f165ae1837304acad367409b2e5e6d49794e218ab0753fd8056d02a0c4b4374b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5dd9c6a7ca3832cfa70f796874ecd5a5f3469e21a657b9736fb8a0f29451a679980bafe068a5fdb3e2ff03ce4d1862dba0a1c10e8932c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h960278ec7192488433a6e5913b0f80b2b490a00e09d7b7156322c9c156b7eae8366f4436d63e53d8e2470fd620673de9f0d04a8065be1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b6e2648f1c77feb3cb35d20645b7b3950d2343562a57dc8cc3f3b64e219f18a9d779a04024012fa850f23785ef68640b88b48cda0448a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2ed14544d5fda45ffa27e07011c828d9414edb12e18994efcaa57d62d1d9cc384cf9f6809ed3c4925b03d255837af7a08e5ae8128cff8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1810d41bbb9fedf71c3bfdbf83923db7e11e2d452a568ed67176fdaca39deba344e0da374f15a054d9215bd6e35b96fc4982bc5dd9a338;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31f1e93e9b8ce1b78cf705468fc868c606ec4abdb90c32a8d7bfe66ff4b3f668a58ed4653aedb9357ebc5c5a71f7f7a6cf81892057fb47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7358a6249589eb0b0f4c2e0497bb83fcfadaefdc758ac65f848f41cd51e35cbc787ccff5a1bb34b59f3449e5aed5026b26ea9a9240a776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53366e7c07ccd1513ae22df01641f2173110c1b0a80074a4e367b403395f4d58e4a297f7aa912d520d794c5388a3fb567604d11e87dfda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118c49e67fdcc665b188f0ece8aaeab0f034784394a9ee7a2f597e88b69e3b0bfab6224fefe5814af7b6b2dc0982b9a052c283ecb33feb5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha92a4461967c11a0f6a5e950a6ea25b1e1c735720781351839b065698e3b1ea69cd1dacd97c2abc403561c9cb5284f80bea021f0a90481;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4bf3b4338e2bfffa1b518313307c282cf532954447c169fc7339ae39f6c19948fce0ceb79943baec6d55c1ac3fc80f9e8d073235db63b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198025408fd31c3321dd430cb8c6312003aae2fad0360cfbd501c8587cba6c66e5d16d754e3d2b3f5f2d613dab605d77381c8d88f06d97d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2185cf5f0268785f96648c197dea6ad03245d6eb0a03474a2c878d2edfd1b460583f44c7db6f0145c9eff53237d2ee0dba4ff31af58b24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e76768f33b32f9e1a1a56a2cbddbca981321e36eceed2e0f510d0937884e4ab5762bf2fb16aad49825b28fcae9b455748c1a32aa91837;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138cca0af0b16faeded664b1d18af1290f965b6a6faaedcfc76202e541cc7064837074ace4c571492a7e8599b8331ea8d0d32022edd748c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ec65af7f2c4479cb3940e5c4e6fbaaa16bd6a33f6071ebcfb762e22870dff3d86b474137dc8ee962cd5f6dce25f4a6576f8ee2706c72a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb04b27112ac32c2f7fb1d67c56024337edf2f1dffef745f5329dbf9a8b72bc64bfb7716f7a8ad6818ccab0d5b9218a26a0e4189f917963;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h444aaf5c70209b37a38fac885466830ff3ac7018f4323a0604dff095a7cfd07a895fa464979741bc65d8a1788e0a673310de14fbca93ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11443f912195534e3760c96b3aec1f42f596413cc21ba5d4cd97072f59ab6c1e9607ce12a5b61fd12060321fdad125ee9216454000d4dec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abfcea4367d419f9f7703ab8f6fa77572b5ec2261972fc3e3208c65260dd57c54883d791b19f5efd4f93a816382c1869215e4dd1d68f07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2e560395d83e56e0afbb976b7e11b15c8ec8ea0a6cba333fa48ed04cc017ac973ea5a698eb876075677cf6e58d743b6741a885996326f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9c9462c11e1697228c018856c13878a860b017b65788aee090b733ca04431e023e8d51a92784bbd0084b98abff4297b1f973c55b7310b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18fa5af24fdc71a5868f10bbeca65da7d31e957f1b051b0269256a93fe1466525ade521778e428676466f620c898c1c98c5ae2cdfc954bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9dfe53c464e455c6cd6c0c1dd6c7de8e227511e17736f98850673e98dd8291dfdeea718ef7c3c5d603dd4dc5273d182bd0f84376f522a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h355f366a81797d87954384a4e8fe4868052127b4d82deca16a04b65e8e77b461ef76e1f5e495e09d3fbb9e4fdc81ff7a38661306f29837;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12df30c01dec516f8e999a1dab323cef189b96bdb4420296752566dabf10e0d8f13246683557ab4ab708e20beadee3054a34a00ffb1d24e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8b8ee3f9777951d4881680a87e5c42166b687279bb3feec9487deeb89c8ac1f4c7e226d3395998bcb0d90ac3f8aeff309a8cef3dbc6c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11dbe21b346b48c876114669451b04d0a1c87e4671057aa3bac8d69ffab5b30b0806255a164026db92a4e4ff1fb61ac0bf608e4af3a1205;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c9f9490412970055488809877e643b47692b7f238cce0af3563188084c30663feba4003e4bda106a487a565937018605d1ef37be5cde;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c5479aea571deadecdfc2dae33427c0cf91af8f0e7ff14a37bc9f430651a0fa3bcca6c9b4d0e90b27d27c2afcddd58cd82298820587f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccb38678b46b28e31e951c4233f5e14e703cb994aa52cbc57681c43f3965a9175e7b6f41dd17482e148bdc24646bb18e951f2e0e6d8c06;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15884f78b83e829bd449db862104006cd3e6936d69c320782d628e6c51813b2cf69f70e195cb23014d08a17ca9c49d2fa0f96962f49aea4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acde596529f4cc51ee62ed03eff5295111316e4b139a423de8f7bd98f3ebed04fb0307dcf6b6d86a906768dfe03256c93afc5e1c85bc75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcea4048b7635b4a55e8d1458e5a7032e08f882b7eedc1ee921e2a5c96efcff5ae633dcf76d5621774384ca00f0b19aa66c7b08438eea63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104a4c284150d92650df0e52a9e537acaf7ff99684818329da24b40fd2a6af9a5c59ef83f5b5310025984d63c1e47e4376f40713c9ea3bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ff25ac2ad22db19ca6142562bc7c69111cf9c3b67c44c8e513a871c609a18dae752d8cd89ef47b821033c26d2f81e7e3ba40e0410a451;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd92b78db27da77d136ab876a33bd4acb5098a89ee57a1b48231f86a72f1b1c56653d6e9ff127b1ec4e7d83a66b17b580ed8adb62fd306;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h728d37435728162828a0263f710ba5b543210c6d087f2277f9610b2dabaf8ec689d6c2db65c52f83fc7af9086adee31d43459123a2bf9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddedc19904f1734fbd501fbfb7ed03b77b7e6151678686875994886048dbd3a5060323684d78c1ba1b5d26c688b8fa0d812a586b5d61aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e1fea51c93290a7eb615c349f6b4dcd11028f520c4c2e13e2f7a57e5739489f875d5f5f4450556d1973c9d1991f8e4b2498ab20367685;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4cab5acdb47429d9079ddb36afa6f7a5df806dd6e136c5e315e5c2bcc529b6e5a65fc49ef35dfc7a83043ff0242814c8a7736ef84fe2c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18573a387a8e42863dd51cbb94f89ed48bed34c48ef94504067299b21f713ef2cb34856d3493e4dd7425e9dff84a1ff80a43c1ae6bc7b87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9d630ac9d3dd18c421a7b1a48c374e669bb1062313199209b5fb00e8c3c122fdd2a159a76e1c021741d5d3d39440eee9c1baafe32e1c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40770f2dd27c7677cd21a3ac9ed6f0627d15d9ad6ab6804af6c90179ffd25ed2ac90529c16fe63e5d8facfd55ddfdf54e51f0718293d00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a662cf6ae9dba718ac2c7bfa15849bb2e291093d134392e12e0871f15f2e5b01f9072226d5967b2667ba7b0d92df62f28a07df173ea516;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19aaa7195d8dca01b0076c115957cc4465e57fed644ea42c2afbada37b4a8d39005cf908c8dee4914b98d07a28556ea837bb9c081b53880;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d81256f3b48bc6751b539807e7b85ffe1b84c60ff1c19584b44224c8db8019a3c4d4e7b8138c804b0a117e11a568968e14c05a2524b086;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0e4a7cc5e18a6deb1771beb690d8c87d30809377d8364c6a4ef41e144fbdc6253460d2c731baaac4b0a21f7d3cee3713e42789f74206d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5da90176bfb02940deb6a9a6b2ca9b61135f01b6d5aaaf4e3ff85e4630739c8ea79b93246abf020b5360e28966313e068dccbff7fa8150;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h659e5e952c39cdffa384cebcf1d9859df7af12e0721a7717ebbec86f0ef5bf52457a9613c4eefb0ecd6eb6d2abd840a4557f462eb001b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1450e1c3122b5bb1f60fbe1e088d0885448ba8d34e684bf8820e482d17c71309d53bceec41b5f61143150f84ad054e502e3f80177a0f38d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haba453b024c973264d6821dae9c9c0bf3d04e81661b127aa6486782ba94b891c6835c4f201861e794b1f17f0d962868ea79b63a03bf326;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h68e038f8f0ccec93df2e29de9516949b71ca9a908c38b79699c8a4f7791f314ae99ebbf3a2415af15f16bba52f434e6228dab5034416dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13530c7e4f1e98e79b6c0308ff3c8f860f29b4099192290d15ecb9316841d444c72e8a07906e355d3170363306ad463d4afc5d3ab3c85bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f46dfbbea192c795df58e71ba15c0be75ffb09fab9f444264dac55c64af60bfbc00aa875d10e86a1b8edf51a0cf50e1c53e86c55fae7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1004f8aba1179322022506bc9b16a3b0140318b73b39574d474141d09830b314187196abdb901642ce1f29649a9f881337ced14628423fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56f9e9f4437816e02011b36064293d66be21d9099e194c41d5d50ad97047c792c8e90ebee8dccc3c47bcb64524914a53a2711c1adba35a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h725ae88bdce494bca96d31bcc49bff1082dff1e13cbea46f0a8cb08f7ed32bb5e24d33c2fdefb32814be6d19889a70677341a9f2042c8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111a1e6d972ed5881f7315ce7cae6f8cfc4d50673b1ee0c006b7f986fc0d6d982940ad6bd4095bf826b424df8e0c618a8979aa491055f6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe93f6e1d11265fb838ce1753b403b7915605881c454c19ec8b9b9ee30a7bd8e3b2c3d7c696906344ebf066c2fbaf89c3a642b70548970;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33bcdec3a87f653c18c4ef593ebfd460253b14ac32c3f56aa3e8dbf64f53fcdfdc981b50a2bca42cf5aaf0c254dbfbf8c518cf627a4475;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110d8a855faf642ded92cf667c0a8c86686a365ace2a54dafe3d057a75a7a5ca0d12e36f2ea04b553d79b98f8809a0bdcf193810ea245ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h154e7cf2db250e9311b11eb351c6bbf5bb5617ac4ad6941c9b458a59d85020b51950d2e444013dfc1397b94e91a54b61c81c62b66c993b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17611941f557b4c4e0f4dd590f1a9f0ab8fe5f81f8e031aac1b49f0c4eae48758059cf48365ee8d4b5e00c62978fe3d30f6494d06c6e9f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9be99d8908f4ed5fa9c88c26f9299d014d6e7ab7fd549e478cbaecb33ce859cf654b5ac2e8369a5ab2daf0fd8c3442c5a09993b8308d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f1122bd55b9db8e5a3f1d4379d411a3cb0acf9cdd815b486af9f7503edce486f3e28a7218ee1b3368379ca64d9b23b29400e9ba5f7f89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16bda82eabb4ebddb4fe6c240c57e96af6987bb6df7de0305550db87f765b4f05d17147af7191a39df2c59a8f286f9fcf234f4ef779b67e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a01a59bd0a4f6ebaf7f9ef24fa49122adb5759bac83d2290d7cea88f36c3e8f0767621e9c6c442c8bce1c0726fb4cbce48d25f6a8fe0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9f78cd3e4eccfa792c42159e1207be0db720828380abb9de6bc59a145688321df2fff8f8734ed056fb6f65464fb785c349962cccf9eaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51d714574797e7321a951a0e0590576dc859be75c6be0dda26cc197672be07e8b947c05e5073741bf77014aa69853f1aba532604fa57b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9bfa1fc0218676751ce0c726d758cf43609088795ce89bffbe66001ec6104feeb39fc186340a6e7de19ca831a1db605de9c8029775b1c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171515bbf1bee8912edafc5874c63eb54603864818e024ee9acda0aa583be3b5eae55dd6468480ebd294c9b1e48fde1b9cffee7aa1cc3c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1faa110ea8bdc62b3ab15b83d7fb2a3ebf1497502e0fcd4a3b4e141adcad54762aa949e57c1320f7c05e7a030465d1762e117e8467c9f70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hedae676236ffbb187973cd939bbf84f659b1ac9010214b679f131b56512f7fc759a8fc0777aec942ed0de9fac2855847a5a6ed605f1135;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3294a6634bdca8f086fee431a3f4a48c78f7ef95e0d2604ac7148bb177382efd07d101deadfdd21dfef83f69ef05047450a6a294c81e77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b1914a7de8ec457ac67471466c08ae3c13d6f66855afe86b1aea0415fbe5e91c547e7a786143d888a8bd71756a97ca8281d3c0c758c43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h641a62e081560314995e95d81a3d7425affce1b838bf05026014a53c464808d87e00824be75487acf8c38546d2352b7e1be9eb6c4594eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134c1811291eea8215502c5d6b4859289db256c3721191cd6fbffbae4091e0707a95c36664c25e7e71c72a363b824a829a58a89252adee6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbaea27f241d47bff2df3250741c6ab8f87318f0ee250fbe94fb5b65bcda1e0323cbb94874094e296dde564ea3d537fda50aba0bfb5b125;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b720cf3b2e3a121c1962348e19d4e32a913dbe2bad57ef854518ec25622a14c43296213c566f33f45e1658ab17a2dd517db7b2345e7dc2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97227a8d3cd97589fe7eb2d7e1c6a8ef047f8d33e90f73751ef97c03c9de97cd3463e2fb2f3dd2d0d107242b30b181475b2ecf7acf3bb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15000ed4b9cf83fefe3cbe867b13835f228f2b40449d3ca123a2c8f801107f39ec321fd1836a3c57f0c04663e0d0bd1c2e3057641d4b11e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1778216765a904006870bad6d2b52ae3e49055d6a6c8a82a4d31985402ec1d463f8cdf002b94a2c60c2a87020705e40b7303f2d327c0962;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e5b9634040b46a51ee7065f50f1bc3551e943f3a9813f1ebc312d88efcd752bebd6f1479c5821c16015e9b6e14922c95622c3cc03710b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf04032a7a579119cbf8f49b2805d813dc3d523867bc176330f9c62d8b287e0dbedc94f11be17ed63e7308c01aafe3c8056813ab80173ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8be37622a2f94bccb80a22f36f79ee05e97d88af4e4e6b7c8972ef1027bed0c9c1db0c197c8cb0121ef9e919692aff6e6d877dcacfee3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2633166371062edee6f9e4a9ad7f64b6d5eba5dc174e1112e723ca374b8a8f90df30be87511d05e1e59a800a8a64e95d453c4da78c0f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1552b1d184888ddf9d8f1a7dd3beeaaaf12d1272145b9ecf2c0113f4e554df09e851b518a68f7ef6079e3fb5dbd00aacf289941b84d8fab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12162f555f740dccf0afbf0e698a1ffa3382fbad00110f583447b051220412e73c34d7a849c10bb7abd1d44a3b0bc00dbf61d5b4cb75aa9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1b225a8fb9cf89824f95c30e2bfab1d9165e8a6b826c97ae2f5bf3c22435b534d07257d2e1e35faa84d15a5df1cbf47703192cbe6f826;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdebb6d50d0f6ce5e1676bf3b060fab427ef83d0ccf210d03cf9a970df87809bb7aa1f3cb307f9c407384530c01eacca155c8487c7a215f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bed1db12a62cce60a3c2ffb04a75cbb7868db552b48069cd047624c61b57fa3ef07e1e35de409f21ac01ee5f190ab16cbe2124f0686fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e10b9662a04e42706b82771938392d14130e94db27bb9cf3b5ebfbf6a7fe391154a5de5d76fd71a3062ca0aaaa9a62194558762e6b54f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd77adbf7e98cedd4118667dbe4c40a6a4913548b8537c4c6e3d19a70d2fe655a53f4deabcdd47de15d36696810d1d394ebff3b27aa3b43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h367639ac6372b5c26e0bff30aa089ac7f535d7e2336ea9d369f852923f5d3c0ef4a5713a03a868369907f6a41b0acd2aac5b8a09a536c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcae0ab753a88ec914d16fff33a36fbefe37c78512df595995fd8bb7f4ea87154e714d54ba4a502bdfaf871ec74d28be11c4d94f08f76d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce1426cd3f63aa16c8d3a914a7c18e0f9d68827ca5e9cd3cceb7e6ee4ed72d6a2018d0e132c5846e7d81946fa64529bf6c6835a7027a00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5a554693a0cb06dfe3a5cafddc51f8cfa2aa156ab8a4c55167e2119d0a1f26d13745627e198a23f652b05417e1ef53411d48e7949d6eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1557c196c6dff2d2d3374a297a864ceb9b32405d4f1eb5e3a4cd8ab4ae6c8dc44601908c72d6c359aa3e570887542880e88cff2ce0a35ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13429c30a9a9b1cd53c573796895bd3c29c3f2f19b72bbb3f02ca027fea38fe23112eaaac8f9719ae756f55325ee384ceae6acbbab68f75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134d32dcd4cfcad9a0325a3c3112528697988a1072678eec034089b8bff223a58aa3167ca3f861a6e609bf8aaf6df57cb2fa81a2bdc926f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192d9a197ee00664e0e0c731805d6cd868c10e6873a5a95cc811df0267aa0f876a06b822360d7b4d66be8d21960ea53d6dc54e7c66ff33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113c85a251e2cfa01a766c93d9acb2fa1947d306d58931f3cfd5a15f59cdaa76f28362ddef49885061762900dd267ece8b3b1f0399c6c9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f2b41fbfb5ccdc596ddc31722af449907bbb670f46ed7de1149c3acc12da0d0b4e007c5055e181dc126ce20e8694ac28666a189ab6d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc54089d8de9894f64683426ec0b4ac54b8366865e6bf558b9e6aaff096905ad6aea5e3906657efaaad17323674fd0cff3304d4ca9b31f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd80d215eb1b6e1efcb244341011b0456ed06d74312cdc6ef50dc364f2e2197df09d922540cd954a0ca4ea9f8d01470283a213e2f4fca2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41664a5680c1b3e59369e326b849ac0eaee5a626e9dd14adaa998088c5289a826299f2b7413d5e350de0feddab0e4d522a650188af11ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95393fd390117f1b291a4daaa63154f1afab943215f7ea2ee959d8f87885fd60c5f7d67fcc8d0ce85dc62694402c4745aab27fc80ec056;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2d1982659e1caaafb7b9c6529efb3d43a2f36d263b7c163a6097db72f75b267cf433222360268088efc6237c0ab78312015097dcd720f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36c45e6c2acb4070bfe42e5cdd509edf66ae7168ab3f23e9db92a8d9ab95bae24099d0af08d9d0afe54c109139ae1de45adb41c10fa04e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1f145ef9da6f72bbc2a21b9cba26dc7c2700f52bf9052d80c5cf91c00cf1930168af0ea29e1535a3bfe750349dc8d95c37c413b7c9659;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2b4e1494b8ff6375d0fc669c0658b489be4ab8565b8f582741ac7a85deaa503d2893a22ccf803a5e8e1e6bf6376e95d3bbdc982bdcbac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf909b8729f913c1f731b0745eaeb8169d2c3e0c29460c055e8888302dff6da2d032c6cf0e123184b1ea387dc2f74be1b0f43cf654a655;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c8bdab4687dfa6760144c86dbb7c0800957ff5df49425de1a7edbe8e199a934e3ef83ed92915bc86752633b2bca992002f77b18735b63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14df43c15f6b870fe73c4d26690a7536ad0beeeaf00390030ecf4278b6436ce66dc7f95c26136c6bd6fea672d58fe0bd60508f4bd498a86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b4b426ebaccca4d6fd7d91e273daec1f23224eae9a01f7a42042afea3baa3a0665480aaa167ae58d8f9e007af0cb327f72594c40a4693;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5cc19cc786845d9dfe4838a5d1de290709bc56e82b70e3eeecbec094ac1d13a900dd59035365dfbba9b4dfb8b5729d733d86e6d43b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c757731cd0090b161f7b4d56bb57342a648360f6f6f9f42b8b0e45c4405565f5782b98bce08fdec4ba0620774b7d4fd934ab1c4e824191;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ecd898875565c7138be630357234962f5cc60dc803bb1e9f3aac64b1d1168d00a0875ffc6fba8e1d17529c65e19109bc37960b702378e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43321b2ed11a78bc085a92f4b471e8e1d97d5e2b421e63f5801e12b73b3cef54ec4c32a9b0a9f13fde7fa40760f96bc88fb8bc6fbd50d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c92542072d1cf142c00f77606eabb2290b2aefc27b51bd93553893e00711d56cd43cd0ab25ade3e0087f40b9844d96ba06607af8e6ef3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a263d4e3c25fb53fa29cbe5d022b5dac796b2e638a10b7a023eab9a5cf3ef997c0cb048de25feea8a00f588e8c926a51f973437fdb118;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf843437331a79a025eeed3c8ebd18cb027f71db3600640cde54fe749b782e9d7f5c7ba5b3c4e30036cbbc41016c46ebd26492b7a5118f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cac623b2ffd9ea39974163776b3217fb3c9fd5d033bc533b5e47737629f51426eda8c34023601393e77fee46dfc801b32001439df6c52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c067af084053f97d1303c8b2088afe4d0df57929b9fffb4249380f16c02225e30eee160c6458a790a28442d0774a8d877c46912daa532;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4253ea692d0c8936d0c85c0045f79a77718c935e34d1802d3b5a9fa9a4c329813a11121f5ca9897578d8e3849fbe6b3b101a9333b43b19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfbbc927984443bbf6d920522d758f45f7bfab9550bbf20d13b47d2dd048d2614d1f838e39c538eef0c263fcaba7c0c27adc1f980b27ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc9226f31019464aca3666a494c23249bee85fc09c232a5409e8e472a46a4b309aa2124c5707bf53698990d630eb46b884159bbb3786;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74a076fbad3915087eb84d8c6cea1ddd39134a9844bd75fedef8ba499cc0f46885be77f3f63d870021dea0028d4e0558b195b429038ff6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de0965190d92097fa1c369bc3178f4a04813c281d209bb8e6701301a8f5ea1eaec3e180b2780efd76437626dc5d3d01d4b0e32c4931096;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bcefbaefea580a4240af67dbc10e1ed877cac44d18c8c5167706a6740dabd0a26787f1e6088706522b0038983e4d7504679eb517e2d9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h280c8f8079d0f2b0cdde70dc4fbdde1c8c4a2372bd0eee6d43456cac2b2a42a906409cb486c7ed0fba09bf03302ce4f8194baafe72281d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1400efd36dfd13af61c9eb43ed00e3b5ccc637ad88ad5463a4a33c67e5a09da9304e1b22f96cdcd6cc7e6434e4728f8b94bc23978a1c9af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1135ded5ce38336be57e6e5b8d2ffb2a0a388743a9457bf0e7e094999d544828ed58e5dfcd8bab91ca45dd0e7f8155e39de3ca9a240b98d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9fc0093c7254c7e0f9c352261869ef026295674fce933ac206b477576883661d76817ffe39df11fb22b591e7afb096821fc98c6115c3c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b442b8129bc7af462595db29327f19c74f2467255382e69bbf2ac9ac54b79a73482d2a7438712ef5c7a952f117af754b60ac45795798a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6281beb159cec8cf1eb226992c0b4b57a04ba53ac7387c667ecf62ad3d24eb4b616ecc29ce4b2aeacb0bd7e62b725287edf8ca1257a1ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb44501477f966c81110f96ec48a8bf7bbd1064cd376d9a761e623567627f878d8729aecb3fa277cffd9bfa4ad1e052e4486453cebe039;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0ae3bc55590e3e0c948c90aee741d24d7c451dc266f40fd332a7e9b54f568b95171bc4f8776edfcae9186178d21494cf6ffb6cfae5197;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163c36f2f7f57c921918654df3d4b5260a0a1cfa3c945695df32f064140d042217d7c2a3a11f245c0f8fcaf35c5883bddbf9f1acaa4c339;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66503e3eac8748c65f293a2bfce9d1d504b7ce97a9005a412a66a0badd096136d3331f7d9b6761f756f774a4bf39587b0d10673317c589;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdfc752ae064099307190987a407f5d633dd8ce3cf79099ed23ee1f3b7b34401b48f2a28ea45a238df8812d46ff27d0e030e80d2ad8ff9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10906263b5f5bc27690f63fc5ea476054405eea333e02efa7455fbb7117ac0a1e1a917b651652c0f5ac6a1eb9ba8cc506978ec8a357edc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d4f3030b81fcda00e5c61d1481878bc4e6b5864238fbe39befc858535e3c5cdb9f4f0e33d1b1a10bccdb6fed16c02eada0f6acfe5ddf1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h706115551b56c34a761650e420741334b9b403d4dc6d998d79891a7c725d400fd114548f5b6e05ec241419cbeb3e560d08879afd78e036;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cd56f4ca0c437a80723608bc1ca4315cea9d2abbe1936558fbe4096bf48ba2a80313c2c2cc0e06545a041943607262dd6104d084aab72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d53918bc5f99621410821af3d987d93e99fee12c6596e927b4536a177214fd2a78db5c6b814f12e7072ce4fe2866c9ee95db98ec91cbc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d1535ea59ff67225c216c4b1e1114a9ed6724f860a2ae59fc0c8178840d6639e1b1746b1a6427252686547596d1f67e4187f172e13544;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166d62fd91a7a0c8b1c3e0fc332abe0cd77ba5ce26329a7ac55f80f721823d118bc12ec6fed85be38594c890962162e21372aa819609410;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15fc8c89bb7417c2ecd537e411a195c3e99520ec8501234322d6d63f4f4b0bf0972f167834d37cda556606b3db4d0df3f231345c0e6ba7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b0fb16287025742457d061a9233cba204076e5c383e8dbf441956170277f8e466a5c52ab219b1c88b71bd895b7a26545ceabac2a57262;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7a84b0842d63a6c3934fa2ff1df0d07b6c6ea866b88abe304148a9ef6b3441101a5f2c32e6d9b444df55b34a1125ead391ad43ac40d2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dfa5b37b09f46a20fc409b5e43a079af7321d68cc78916b9a781b69af3733ca1c87ac255822f17446acbebd562900e00d7f09f11606d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf194ffda3d8cff1c0cac2db1ddf80f1283dbf7943fd1a954aa47607c23dedc4ec25309f1aabd2ca2f1130010a968ffbd6f28431fd7fd81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb0ccf03f70784fea3eccd399fb512cbc6a51eaada02e24d7819bfb581f9e3ce0372db80ee428892ca987515e5508a004170d48d5248ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c0e4d660d5d1944f10cd7fd641a0b31c4694f0f021f2a385163ab54587d5707c92b9ee5d3d6313c9ff78ec423d7a76dad109f35e70855;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1fa0448c8aadfa5c8cbda2db7081eef5f19f57a7c380b3e2060a932aca038c5a7cacc48a4f14fa4982dd8666aadaad1e3249ea3f2412b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10496e6d011ae2e3547bfd68b06d164fc1ecf30f1840eb758142cf84784e0b188943a574c8b38242b2603e23a292a49bbd04fc5c67efa73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c90ea1a1fa22cf04ceb613a55c1e993728e33758aa8cf58beb7feb5f85e439c5f7e4fa54507c2f38f444276596516ed2a5a75032eda35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1869add36abf66bd39cdf7f11e64029f397705671d7b819ea795d2dc2130b72d2ebe9d938d48263aae595d08cef0c481abf8ba4d278b41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h316071c6796c965b363895a0b59e4f52708dd5728e121b0d738c4a03063e15912c68bac04d6e4ba0de9c37a1650a546c8b4b0cd341ee01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e47047dd11fe01fc497123dc7c98296ae3c060f3fc363efa12612b0715e192cd47f0c105206c89ed8c3b5e78f3d7bd2e50b716fad7164;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8f38231a998a6ab647f7c19ca54ceaba3339600f36e0e7813afd5f67cb4c27b4fc1419d3f539726274b9585952093b12baec157dd37c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18984f7a474a7c4b12219644276b486304e291cfc7e61758e7b2e4f9884ea8accca62388ee752625a0a32b88b216debc33dcf74b1dbd53e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddcef00b7cad65c8c025fd37b2e0cd952ccdf19edc8e7fecaf14f4f0b300ef2a90fe76e6dce9b22157b0d236a99c9506c91c22b920f826;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha594f4b979738f2c201557db1db096c0b52e10dced11dc099058264162c12bbaaaaa170a0a1fdd8b14f8e00be01da92336f63b8f49303d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bcf050fbf31a68da24883b6bb343144c1a5a12a9dcb8f434a59410e17608558e1e530201ef262fcdecd928b75167a2ef8f25692025ec5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1276348eb8db6b2d084042d83758752712619c65c1a38519f62519abe82e7e5590c4ec9d1ea39b1b2841fb5169e7947af1674adb6c47ba4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4074d0c7e4010f73b61e1a3d9ab8f43f4199595de4fed2afba6e92ff1410f37d10936079e539239bc7b03288228168466a8fb7c8420b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d97f665614936bf159d2951ed2ecca8b8930bc26ce80fa7155c4a49ff39216a43ca95ba1b9de037ae3aca7007cf6786c53cb6b9d7b76e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2d0a791369dd521716c582f7c6bfedafc2476e0010cd772ba1aaa0843ca562a5e5e2546e6c73027ac2271b3641b8c619f8c63d166ed90;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccc7ed3fc472a0329ef12cb0a5177b07447b6c6568a17c5e3b6d3d920115112ffdcf9df4016e94e80d2f62f31ece09ca6ef39fd7690cac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5b3c1d2bfa59512d7fd184f65865188fb8cc1dfa980b8e0870223a84a83d0b9009370931f0891efff7adc06199aa9cba4f015d98c49f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b676a343cfd7b06b3766e413c2e9040de6c0769cf866894b6427df60a7a6cb1dbd5726b764a1ca46362ead53a5b2f8d68ae94a7c1bf3df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a04d83c88b2a76644e0c62094053f7fed720ea4fe20ae00090149d3fddbe91ffd567b0be76ca2cad530eba0b5893600091528caa8f6ab3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bd9da444300b89b2534952b0b8a3758e64e2af797c2c8c31574acc2a64d657fa4cb50392ba42aaec323a65ec1a20cd4f8568f7d9889e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8bd3796852d3060855a898a786c37d69450d4dc2c90df50eeeb918a59f1dd6af870e6d9452a314776759654a75166d0e4be30d9fd7587;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ae9b1f407b4c359b9362717d1f2f2fc7454f3735826d687ca8fe9f7d8b96e81fe57af433b7e143e7dabc36b3f280a34e1eff726517054;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53bf8a911ddc891ee8984140c66f987aada2bf42a64dd42dfe9375fc19f63c8331d25c35a99521b5b57a07e55628926ec9c5209d4f7744;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e75b921fa36be8cdce8d349c667484bf99e11501fb296396f520a3ff2fd29f8c7e8aa0287918f802d4fe8627af2c82badafbc8ddc25a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a09b014cc216aff7908b962dac04f094c3866b4d732622be7f20a014c6d5c0855fb6982053eaebf04c9f9170b2b2454ad79088c517fa1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h779981e4c5b40b96645f948293d996e25ad8f33a884b5cc5bdb060049c2dda6fe01b4ea24b3f7f1c30042b052f63afa46bad6244ad8d60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8de9064d9ae5418af422a704dd7334a0ddf091a3873a0c99d612f11aff0892b7c42f48578bff3199c8d82466528297e60b7c4c4aca3fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16127030afa71939fb0b45651e2b913d3b594a3da2f667e1f777a7302d7ce575381be2bc0666c7508c782787b6b844daeba115a6a738acb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb533b9ab41ed46b039e42dc7f9c1f119c6b4f3811a746f48e38140039939fe25db54139d787dae64b246b5536a24d8e6e441d620963f0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97602877af107400a090df29f01f6ca5dbd77dcd01419eb2baee3115bbc5106d4eada708ef85e076273ee9f417f9f2d8f708ac63ac4c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e89d6a1cde3b36d6607fc036559d82567e3be2d4b32d212186b0a8e8e4589b05700a281fee53f520d48574014fced746b4d404ab3ed5e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eac5795f3fd56c4618ced276205b69cfcd6263be5fd6c859e4bcb9c264bbc20feaac2c2fca93ec2d7e55f96d1cf17cf3b0e381ea600144;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1e3cb2c2081b43ef09120beec979aa6a5344e6a11b838fdba2751e7cc33572e786596b60bf23364a22ddb85f63fbf3d96c218274b1bfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h245e7081bce11b3897ce45fc990bb639a79fb83f8489534084e5e4e484fb6cfa103bb2a0b8f996acf8a70922a292298d0ec1b280d300e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9fdd7dfc59c9bd9a5a17b9fbb39c448914812aa25e04f6f0a815050975363a0a47a024c6e99c715aa75a981d97db8bc22faac265a7466;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b71a6a67aff41235fcaaf9054adb3857a82db0832d94e5a8e9fcd02bbfa28a853715ec0ddeb1bbd33d8272e627953b6a626164cb890fdb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b16449aa7b2b5165f32a8fb71519591f265c9d78608ec4cc10101184e057dbeeab49ebf43ec53b7886a03c611d296b7f09512f316d6ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc464a175c449c733bed2f8f3fe6a28b5320a4e029c17769111100d11fb729db6ae18580034989af199af5761c461befd49c22902909ad4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc099e8a2aff7bea26621373977ac80789e17c5a933554bd17696993515f2a5ff3893a4080bdea8a221c35abb84fa7237be379e7e6ee48a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11198b0823b9aea5db192052cd98ba4e09197730a8e7fd0f75272c449b8acd15f0f570efcf9cd9a15335a0e8845063a903f0f7c20991719;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40da733904c065397304d02f3e5835c67f54efa8dabfa9957c4a1aecebf6b86e748d609e62a5800559a072181bb90e7cbc188e2b508b4e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd36010f2030b0c99f7c75b9d420c1b02193c03a1352f4a4147c2cc739c32c2453fb782091a949a44d293b3837b881ed71d24f88f237a2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142eea4a50a4102ee2ea278a7a1e89a4dac007377683ad3709c5a7340a653ece5441dc5a42cb19732b23c50c49deaa019b7ceb4456f35b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc78400cbd5a83f0b72e875810bef89ed649cdc9d49285a86b863cdc2e5b32d2632814864bc4afd91b9c5b973de0f73741832b85394b9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f57b539e1ee74f3d25fc2ed478ac5bee504f5a8c017660860e7972bf2a651368857b5fe0f52186e65682739c99a6bdb3d2ec7b0d58039;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145861a11cf5744796c277a35ec46aef907e3ebe575bf5c8ec6b864fd05449bf51ad20b9526e5de677af06941b1f01e7f63a9b2bc291e9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc39d08523a7a2195034371c01406088715c0631848ab4c893ecdf19f5bb0b0bfc21fc5036fb0fddb29ffd03826b0290997bf938b9bb369;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b172426fb55c6d9ba637312af0cba38c895c339d9693b0bcc0941307395472851b5598539494e97166411a933f7bcce15b85c0d8cad52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188de6aea1ae3c7c75e003701e7ee31e94db500efef7da9fbe078ab747a00d0adf8048357090e2769da50f05f48d28a1e2c2249e51a7c90;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3289f687aff07e18279714f1d08a100070bb52820edeb0e8e3cdd9e260bd3007722c069b3c25c4f032f77e5b2e8c271ba587c43436e52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he22de50deff45deb08846a7ffad2c63fd885cd0ab2ddbf1eae5cb0beecef01608ce9dfc173c799f191a3f329c83e5444e5588812138ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157034bea181d56c6defa9efda7cada851819e62a9554b85670d4252d02de5e09be46e7f8a46fa6ebd0709ad4c9c703998ec4d133a3a041;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82e538bef6f0ac0c70412c62be3dbf32efbaa979bc219c972342415bc0c5f9762cc117ac30744783cf99e0e6391a2f29d58fc38a3f899b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d6da34e698374778501ff8e4d0c75b3531393865ff2b63ce3860abe7e1e89cad557bf26c6d15efb343c81d645bc8295bb3af0b08c7616;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5797f453301baabc86841b01fc972cbbdcbe3d5a70d2598dc685af1d4fe575db8a2484f8c058204273a40c1d8afc15a36a0907aff3bbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2e16179df4a070135870fb5d2ead2e904173a1122a1ecdbe6df721c60f5645d6419b49955a29a2bdfadcb74ff33375bc002c259b82879;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b80a70c6ca4a6d97edd0615f37f389d373022c46c07ab856cc1944112709d20ded322045fb208e4c370b4389d097d799668e2eca47d67;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h841ec879596f94f7652606b762d12669af9741027bf4cdd01ae8bbf074fd2c22bcbacf1f7edf1b4babc25edbc9fd0dd53e3cb528c67e18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156f555dda896b47dc1670814a58ac3cbbf8329ff970370ba92297af51cfd5b4025baef84673ea062014a1c91549c2aa53a4f7180d636c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174d6506fab65734057d2caf41f8c2fea93829d6de308c4c85de7e951684fe6993f1b70ee7c2f7290869a2548ef45c2c5939566499e287c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80241a79cec81de0d7af76d98934a0c6362cae2c57c4a109be3370eaba014767fc5eb2fd85cff23d9861d765176861bdae0c1962d5c8c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7a6b868c9c80f253145ad2330a67c36fc1d234f46ca85a4b098345dfd24cfa6351dcef2435ea6154b4b33dace3c7203bb83e6f63b5155;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc595c2b0f3900c245d4a737cf1dad5644e62c801ab2ef09432d9ae6d55a70734f0711f415ea32c07b3b229a6af0d08d466a3454b2a65fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1172b293fa334c2f020af6340ebcb9d4d64e052a8fcaf0f5f7121c751a3564f75fe3993b8abe938ff139af0616f4db7035e4a7fe5afb6de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81c51a8f25aab131eaa1e90c549c4119894976665aba8d9d9466626f043eca94e5279e5b4256691d747f240fe60d128a6f0567656962ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1704477a0a0080d456d4ea5f51f2dbf399017f71d0cf933a65931ffe57cd7760bb9182754b7838de2f738b0408b51add1dbff04f2ab9c54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4430f1bba17261bb75afbe891aa404f1410c31c2e18b0eec6e42d9cae8c2f6251395c7af71896011bbe64a0f99c4fe98b7d95b2823d250;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c98d977d11faeaf849215d2f825f3462e99d9d5fbe733d695450498cc41f1ddaab82c3967ef46d0e25e391784622179ad3b43658811555;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd7b2a287eb1e3163c383322379966331ae30e1bf487918ee27c09173fc94c9c4ae6c9fd9238b77a9d1a3633b07dc86e592e46864f9d76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170650c3baf82ada828ed19240749afba218b5f7da29869d2e972c070d8a72af8b1b800ed820fb212c0d6a5ee803997ac938fd39eb9ea62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13da45d062f5ba9e576e1f239216edaa1f2f82964cc9a5896bcc5bba8af18850525b9b462740112fbf2f26f15631a5f062b1502bdd00427;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb968c6d1af2f3343f0799c5fc33b2195c7aa481e2e899844be48771046a8cee0803c1d479c3b20a63928803a6d5aa287dbac2168d5eab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca8403b56d8f37b10c9c22d98846abb82cb8325df71518bc77a287bb788c6ceb6c43a2f3817231870027d306dfec0c224f4f2ee9415a0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3584766e256e374d4629058a140dae2bfdfcc18a1f74b48a0fe506eff617f52770cbaf2b58ad0d2334e0275762ea0cdeb236128370e10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf299237477f28ae4d0cad3eebb5ab679d7105a2f4a33c791f56189be9138ef62ce6605de907266b2008e9a6c504054e441b599b881a32b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44071318e2d88c918b054d162bf7b13d717159011223f302cad9daf170fd3c72ef6977e32530f7242c1792c963ee360e3627e1575936fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d32f566f4f4533e163749e51a3ec2edf505b4f218d85bb469e0a2e1db4f0de8738ca908d03f26c37776124223ceb2a09fb6e71f222343;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ead35567a337fe67f43a9c9d63f5549e4d6e4889af4124172fbf4406d27c33a9547b5b8c771125ea42fad20ad68b2a034017008f3561c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e9ab59098480faf312ce72e7726f80571bdbda44937d4721c33cf8ab6606f6bf0ebc72dd28068c06338ffc4381fac5c337bc85ea7f56b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7b772437406e22b6aac403f0129de6a111073c1a7f11c48253ad3ce36b78653d52dceacbff26a50de9249c8fc5d055f201a5e07b74ee7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfcde2e30bb3a3aa6b97af168c71e1b5e0c0e460efce8c8a29f1ac2092f60b3aede48f57e199114ee3a7ef41775f124029433d2c01c7ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2acf4d846bef799ab8a32b4369bb19895a87fc80164b2841ff333b0cafc2bc9d43e5fb99bac19652332434fc63870076da366c7a0c562a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b04b9d10b9532f9304ae2391edb59850e80a31d32058cba7aea95bdec375fcc4a85208187039dbead7ef09abd484c0eb0b715f557d1ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cde13d39e038b9e2eaf75c9efa54601b04be48c5fd15d8ebbe3568b37b6e6fd073127015c19668a42be5726e3883338618ff6b5e4fa9eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7dfbdbe00adf9b121810227e91213519b3f1dab4d8414335a46798eaba907570a4d5ee7c4c84a547ac344d3db028ffd015f81d0ffc7d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140c9241fa9150560f55a1bbeff9117416212a09c307d2c6ddaf244372a17728ef7b1d7cab7172d0a73b200716b5b69db124139a023ee03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120ce6ad64a991c749a090645b2e78bac03c5c6c420f4c73a39d29cdff515eb3c6c5b1edef41d4c43a2f6c8337679319f3225e778658795;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161ea05340a612d818e3837db0c152aaec9ad5b5168efd6cc102e653f8059b4445b0df6d974f090fdd218cff6e08b2122de94651234d316;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6da727ab6132990c06d2e9093980e61d1aecaf30f2415802867560abf2daeb6c803c9e00adf33a2f13fcc0ee07652996e39109d0b41f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1042d14aa31f50fd94e5d873e376c3374e6e3e0f377c2edde2f29472ab26c11ec48ceff47e1282b44014303b0b76fa1add29558ab7703e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he07544e667d014986612c01f9862abbe58d6b50f590cddd5902e2eeba6fe560fc5c7059cc602bcbee651c9ac010fa381a6a46e0686008b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ebcf928d07544e26e09b30cb690e57cb5da64b5937665db3b92d8f515864dd0ee6771f275ed00c02ebdff7f5f086ddb5243a488e913637;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1020fcf630cf5680bdfd0d745f69b76aa428880601301c5dbd20de640635962e768a95eb97eb65cb0e8f5fc5fc215774040a6b748b68770;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e77511707cf1fd0c593927931471887985ce39b056bd10c940bf04eb3b52df4a774183730eee5247b1b22439f803646744f94d048b7a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24aee0adab8000ecb745cee32c371c57542742dba83c561e835a566bfb1bcc829dc7927d108177651ffc57644d8f750c2b0715b1942138;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123cf5808aa34a54eb9963d139c4ea9e1a564b10416b96f788e381fcac0190234e213f63ae7f6fac102c01d1e9a2017b405a8fab076a16c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa9115d667d92f8f054de4e5b6b5e4468fecedba006d317257dedb4d4faea0e03a1a253aa63486ad5196ff14fe5dd4a1ae87bc78466802;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a7ab88a2544314b69e21b236a85b4d3691037bc58428781087138eb8c86b6be1f8840ecba2db56c89959feba792281b60b7682000ee94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb05205fe4ecae5ba6196596c5698245eea2131490f831cd53a6d3eafa67b3668aae3d048da450c2f80e0788562d1541f474ce2b02f276b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b134d3661d6c3f470c4bc1f17692994e43966ca1d0b87f7c9c255150e37298ae8c0df7ed3e7d078a1abc427d5d481881ed183b888fb675;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba769c7087d8e7481e5e647033e5073d92f8f26b37c6200fe74d07c0afa99ed3980cb476c7f842459346979bed5413c3f79c39b4694224;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0e700860173e4f58277862cdf70db30923f11063215c18d43c137cd317e6113b47c8399d3f345c6a4e446642e2b55924351ed88d2d34c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe394b0015ca88fa52ea1c290fb85e1c140519ac53dd3325534890e5a0049f93a29451944a56c0215193861c288169a8e470bcefa378ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd07b89c24b5096d1d056abb4b46a042857f9abd1e69e937c441e0fdf3a4c7446a58be82218ebeeee609c48d34b4838b69eb51fdbdae806;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194292d9eaa35f96d43c9ed648d2c5133321e96ad274ec18bb39e2e4daa19b7d3c586c5011edbb0328f7aa66e480659358e96dc1745fa29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d688e51ab5cdf7e5ef99561a008a636dae53202eab09526c65820da52a0c6cb5ecbf823123800a95fe9d04c3a9526b33fa1011521e42bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed5b87557c9be14e8c8a9083f5619b79f93b285852ccdccc880de50024a6e00559dac531a80314180cd95ee3ab9b9b585ccb665f651b6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fd3d06a621c62073ea96e9da61934c28306b57698cb716d047b5e9aeea79fd9081f61308a56e8392f1b68d7a0f66018d28a938c833888;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96bbad244174e1f8b59007a1179fcce0c94f99161f5d447565037b98af84462c096939ffc4f1606b2db8d204786c787e92bef6cc113204;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c88692255503495edc0daaf3fc2431adcc1ee2c929cb48cd15837fb5cac1aa34d367ca799dfec1139d0a83e755a2ad846de9c4f0791f32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf99582b581a064fb22bf809db85cb7601ac5f4569fdb0ac5b46dccc37a75b099404bd7e97909af6beb313bdadbbe08e7e1488d4b822217;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d4421c0a6a5f0c2ceaaa3945a0025c6eb107c3a7d1d8dbb85ad69598f7b5b3cfc5b35a6a37366609cf62b2fee1660de477bda441ae3d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7487691f76af5b495fe095ab7786d81ad92bad57bf3845b5fe39992610d162eab4728263dd09b94a7b68f9eb0a40e52ec3aec7022c9b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd30586e832a0859e913f2567aaee77bf54f78648c8355fa4ed198cd6e3cb634d9c8fb9abc98798464aa3262023fa6ec142b76ba89950f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65dac686a6cee44daf9a7cca1368005254831702be2834ae9007c97503c66762c2a5f59e38cc1eb644f1819587349801f791c1f5dd20b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd39a581bfec082c0d2889ea375c7eb0f54ecf3738f15b23cdeb5ed730c51ef9cf8e057bcff82a62c5ec345562c5136ae2d50b5068f5cd7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbbe2eef6e9e4f0858f6e45498eb9b925717d52fafc9a429d426909e4fa79e2adf7497d45be1def68a36e577d85438c9a31c6ea412546f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h866733442bc8d7dbf4781cbb5629eb0985cdf10f13086d134946e1b5d704a0c927cee69abf329607357d7dacd526f10577df5c740719a5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a3a5307e2ffb657f0141401e5b71913d735e0e841bc1939cf960ea9e744bb34df3662efd048000663df109f08d3efe8d2e2157ada9b2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d4386b4dc877c26372a3e3958e74d077922c7b7f67dedcfa7076771b79c6128612755dc0aac9d12714053297f7e5af6fa37579d651ac9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a43903647847fae56a85102dd3036ff89d4345f015645ac70f1fcf35663d1c1c208fcd6cb583490d9057ebe6a3632d34ad0e11e94d54b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58f1f5b769941a78b80d7dcb0585bd20a31d59874ce4a0593b0e085cbe3ea2704167b3a22cf0b22e5b0531c37ffdac4417318228b52dd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadffcdd19e754e1aeba7571cdfff175d9b07f6dbce8c429f02a757d31cc4582e91f2fdde54977e62d7c34d23190ea7ee2f0dae8feac893;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0e2be3e70668d459717d2c3cfe16bea0ca77fe16bc2764f1226223c3e392838b4772a4febad45e8751633ad0274eb2b40eba74d58b56d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5f85f00e01e4825289c13c09b7efb340c87e6d6c621d153de61ceb81dcbda3b6b2370a3e5ffa948c7e4a23fd959234cd4d5e9742d0681;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b254137d9d8adbe66bf288369166b2526b5246125d1195f19344e49f0314247eb7ea85592eca084c70cf37ef300cae88633e4633f6d97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125c0c5edbda0a6de4920b4defc1cc7152ca34147f81659c0bbd4c027b9531a472f139c9c8c4bea685ea9d4d4372a788ca938dad4ee9993;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h836d227cfbdf22ba77f886575c8e1238751c87cc509303bfe9f04b152bed1a8a97443e39633cf65bb3fad8ceb1eb0695e882e45a443873;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44dc68a1417ef8b73b8bbd6d1bb4f56cc65a7799ee68e26d25d153621eee0ae1dc92da7c568d224ea7816cf76051e379f211367b3f8c97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142be6aef50602cb7b62f65ffa98e1be8dc39ba02613c826fb54b35b02c28360d80efeccc4f679c42217c432029f56f1a6434aaff4c7c8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4071d415adc8e64523a3e285e79b9ee4199861c398f961b7715fae0da3b93110d1b708d30a828145a37bad0aa43bfc154c1010cabdec8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dce865319d55a19a42bdd0155942f7d7a025111f59462db9542e33719c26b6b71a314e3961a27473536a0efd8806ce4c8535c7e4dbd020;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15035d6ad9892add39b5b94897d359ff200e027228c35e30040e4ccf876e5c7405e70010c5661a07729ee5388fce040fd50bcdd890441ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f90d33362b6e8171441de474464735bb5e6d2643a9c9e184126297553f6d4d795e05ea715e6dab92423f1db2f6cea37abcdcdafdcf7c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70d862c438d93f2e4aba4da0f59d84e14c04bfa8f1e979abafc6e593b961757adfe3805a2c53d1ff58e58124955fde6a3127e68217af2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c644a8b927856ae1ff792b3fc964ccb35eb5e310a83b9f9198a82e38184cfc5985bbb7bdab0f7dd95297f6aa171779ed5226d6f2ce2a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1407f93d9cb46a7e99a25cbc4b326d55319ddc1c5abfb06dfce1688504c124f5304030e0dc54068bfedffdd536cc42f6b59b03bcb64d64a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104bfcc7ebb218047ac690b00914af1da1eb4a542dc6d222e308dc429767593d63ca40d69ac176868b5c22624eb16fd06e41b217cfe68fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed389a9fc5d55c520c74a9dad7ec167a7410cc156aaa9afc541d52ad1214d7ecb2c4f94b1f3fd37a3c66c3e4d14a5c0e48bb2e4c7935a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a806708b03336e03e43986f4509cf2b7ec50263f4b9a08217bdd641393bada4c9d913c870743064a35d27671916927dc8935329a3a92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2f00be0977c125ca90c08b23cce91ee76d8b243c79fed6766a58bd46cc92d83b4b571d52d6389b392ed578456e0c8bd845a630108f636;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddb8433a8c44bab220a61a9e84216b63c2aac8b24c6d7934a403f35bca5e9b9aa64a4b5f1f78b713822c8dd66cb89f279dd4a2ccef3f2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1887a3ef3521562a2b455b1528e7eec8db0b7863fb4fe78a8288703061fa74814f7d60f9b511d6d80fd7083c3b87de4a82e55b74bd97de2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0a50c2ae3feb78bd7001bbf64e03fe317b020de02afe1b712190d70bdb3af4879e45c8cb67a0aebf137811ad06023e551807df706c995;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89bc6a33b9a2db8e3333e8ecec7b604c3755d6c648c2197098d5906f2e56160ae5bd9cec90f53eae123cba71878e12f6ab40e095736e16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1091bcc253ea1d10108550efaa9d06a60425093d34b7120d6ed0c862811efd082e1140ae424178abb755077aca3218d024f7c27217b4458;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16791db90c05450e6fa383005be0694e37525906899e602a14168c5177496bb48777d321dae93e19459936937ec8c12340fa116f0854137;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8eafbec9fb6031c58e7b86a6dac5f3adea4f662aac0a14b08e2f15f1244329825bd591031673c8dbd9e97f44a60509d95fc0847aa1476;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c23b3241f7d1612d66a0f5f889b0ebec33b7b68dbe35596b1544be941149b22e1739a69b423babe3b13cafffefa33c45f83fe78956ef4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d461d8a6f593ad433ebf0dbda8fbfdfc88261c8e6750d0c375534fb21a9dc1a798cbd865af70765f15eb637fe8c35d84d027b07a5a48f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc402e745dd5eb126291d654fa60158b7e4b8414c48126a862cc8d8175f52e46ef6cf631f9bc0f4c7c60a9ad4c8cc87c26679ad11a41b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac3f1ef48254cb1e9af46a21b3ed077f053c6c2c278905c08a4519b2e42de355d7d509a6a4b4abff865629833b13abaa1b203c79c757a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcbbb3ca9a1d3fb12d41d793ffcbd5e6ca6828a3c81912e78ce8ba18a4cf8678da5d92e5e53254e434f982f96850474798f050c2251712;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fc088eddce4d4924bc23d2ce74c1c538a3c90de1ff41c9b152b0c8b11c07ee0616eed4379f1b930b71495a8fb3e840a747988ec03ef29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124104140887325f382d7e577feef3755924c80f0ae51fedd0b63429297dc4a02961663475f98901eabc85850f1dce6779573678abe4964;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3707cea78ff925c112dd5a33ed29d612893cc5da2d9e0d7995ae9732f9c9f1322cd75b52f39354fff56670416c35c86b2ada103ae5c801;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171b4990feaf421af500a38cb36930cf1f9625b546f93618907ea18250e589141ccb4837db6cb75798265c6e55920bf6548af48fe3460e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h543dfea9b360efc7ab00b2db807b5f95092a4b391a41db7acb0497e3818e0e44e79118eb16fc0843a92baf1c3b6156f0e497c04d50a3df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16532b46c1f165ffffde06efadc15563c1c550edf3b820ec52ebf41b03bcbe811412f9abbbeb1eac77335c144b681ba8812ca880608b7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h650ca8352906f7c326c4e5419cf5e42c1797d0097d8dcd259ca18ab6878468688e297e29afdc42973be33f0eb89731b195d1666d7b2be0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4a3417753c8ae089ba7fcf825ff05348f31badcb29ddcc8a799ac996cda5a683476d47285f46bf5f63ee869c97e150e63057eac1e2ae6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146b10b59d9d4968344c6ff04889dc9f0d8199ed3be953e064ae04090b500df5abfd8f40c22a507909fb24f6bf02d87a401281c52a8a334;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3883514d2c4ffcea3589ffaa066e0bfb38fe92162db54ccf6d94e85289906fe407ceb96c183f2fb5f153dd01bdc9cf1c36e38624fbf24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcb6985a2df59650f1bd01bb630155dc2f34e4b1a19388237662bc034e7205288456386bd506e0794aa5e46d7a6abf003911c3ef189fb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf8a7b1f1b8feaeeb2a2d0d907511f2b8d5602bed01ea8426dc347a49f844b067e61bb048cf0c6b7352abc3b3714b8eeeb9ddbfe913996;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188f75b8a817cd4bc84592b0496c27bd20e0b6452a947ff7f3dd0a21be59ee840fd3fb069815afbe8c2612aef8abf9d91bd7c76b0490835;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab666bde5fac522beadf1885371fdcb2b431b8c10e79222196137c2938f1febd21852fb5f5324da54290242a08d195ce75ff581e96424d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcd401721ec27a1521cbba42348bbd9f1addf9207b96401c67c8c69a08ac7075ee26e2d0152913c42c15a474d13f211b1bb151121122ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c693e6017a63eb75a184edc9ea1d856ab8f64f40c34d34dd827a3a76cfa504edba5786b93b49b9b0e469cbcd6a5b2f5a9d526c4251d33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133e46a42cb3ecbba468305cd44c49d60919c20469c7fa9ffde3c729a78a36d63450be962ca1dd68e695a5d6d7367506622151120f4e09f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b0b69bb0477bb2b4d20ac4b9ed3b9348bf5d0757e6cbebc8850fa996a6edf9c184c9477edb52a6952f67b011f23a42cbd06fa9f8b0b60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2de3e7b8394a0885d4a2f32e8e5a36609bcd8cf231902a1eb6733dbe4e59a00171092cf1ec0ef2912a75ce2517df9f8ec6ff0449c63e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10703ef4086a318179f3796c86bf5d30630363a5dc9d85147924238580814d81e10895c29c0f157ed93e18d81ff70e07ea011990ecc8f02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151821b6fb32b3b19f1ae0bcb64f31ce050f620efe5a8b8a05bcb4020d07b1a5370f908bad9a8114f4c8ef99022358b1f8c9d9528c30bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4719a2d8b78f150c635045bac18ab83b6ff6af45cc020b0c44bebeb7f663f76baecb805333adab38385bc754a80f169f063f53aaa717eb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3ab4bb5f4e52b64984786ed14a9238d9ba16686cd248a8621335ec3d1a495fdc667c14b5bce35f88a2448d70a0fad31a067b63e25135c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d19e3a4b808bac61a60f4497824a63cf891fcde2448e8b0d230943220215bd13ada03b2eaa6ff3f21ca5b82a58d6816983e15518971a62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6945e16af800bf043f781215e5f5d3b30174cd79649c614b4c681532c91944de1ea7ea64831c94b83b32608700bb702600840c94fadcb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc451b1c5fbfa5ce14c7c95f4c926288362270f13409e830c07a6db427c81e8c2c87975d805818ca57ba04640d57d11c8419ea9be4c345c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1695f8f79434b6cb063918fe2e858f29055f4f44c0396242fe5debea31e790cf74644b5629853d584b24791cc1c55e43b31732656de8557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h281e10f504315658baa0d4b232489abf0ddeda709a6394b6def331a358b338ae9589da29e4dacdb63a47decb473853fec05213c3e4d7b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94e1d9631c36fa74bbb8853ef1f79b4dbfead241b7314deea8e656de4d931dc82f37d6f5f080def861468093127744de6c416e4f145f18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f389a4de6015044539b7cbf9036019874f0460019e45391f6cf87971aeea59a1ceb2071345deffefc6b4e29c534cf63b543ce41074fce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14cd64d7e515e148dbd54ff41c3285ccd329ba11484a78ba84b6b1b07a0ddbc0f247a6bd3e7bca5dad3952f64ee6aa3db71661877727912;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2899600e7677002758ae9b08685fe9e2b093345c15aafa0097c65b8aaf2688470721eff518458d594b8f40cba5c31f03aef6c7859dabf9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h851bb2f2ec2f79e9407b1762e3c0d48c0705f68ec2000cbe08303846dea2c7a26e414a49a15e4a47679ccbf208e94241722e4cfcf6ce82;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h470f4618b696934aa62a6ea4a0a36b95674840eb11e8961ba4241f22c5ea0258e01c34c25c22bc40b4dc27abb315ba6b7ce200e2c23b9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e0cea0f5186c4f2d748dd6f8a2ce7bb2b00bfbb6264773c3db63b180028cd02ec1692b1ed9a6d7d351eede2cf7e989fd3b57a9327950a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76fc4a1112d6e959be6bd0f127d8475fcf97249583a7eb88a8aaf4fd219765c16b814fb6c32564533d78568f11ff25b047dc25c7e1671e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe0033e87c1797c7a9f9316c1f80a352903a506770c2945baccf2f0dc4d5bfbcf10ae46f51433b4ead42921ceb43084c6425f4fd4ee725;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46d4aa9977f15d0ba76f701777567429b22fe89ba2b08b85585373287d5d625ecfe2e16ecd2fd0783d72fde893fa0dbbf92135d4143b4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3debc4fbec2ff7ad782854c409a7449bd8fb4409a12a6c9e28d8fd549f5b8025f95b0a56f50f902e9fd17c230c00c3a4ac8f0169950c32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7c9453f5348bfb0e9525d2599cea2e8c43659f82ef907ea64cdefb5fb705a01fba430c2f1e08c751a09c598d3063c4c74ba71fd38b88c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c2cc04f7ab4be657754c439729e26fb2dd3ffb36990dea2866968ec952d87160e7ebc2d689777654c354fb62c99bf3836c7601ca4f441;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he53d3da85e57db5c6a4bb369e3d5ad9aef7b0e03c8ddbb32fb970db9b7f80b9446e99adf65b1ca504841803cbe42365d777ed61a54863f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c230389c49582e04928ba37ce02c92ed67dca59202344a21da08a17c2fd6b2aba312f652f060b1878c9ac661aa0e801a3c75ff687fb713;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9e24003411b95435a3f6101bdfb434e982340c6e55d154c1146896db74480bcf942e61c69596b5a18cb289808cd887cc12fd94ebd2c2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1988992e40776c1accf52f617c22c9b9305856010b4d0795accaf811fa7eb6705e5ddf1fb7776f5cc24a06affe15d5ff55943f99eac57f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h330433aaff291c2879673208ded8b2f2e054a051dc3831103ad17efd8e4b8f83e546f7b8d56597f7a16fe491e4306b97e9daf05f67e43e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e8585d3dad3f2fa06f8b8de955f6776c297ce7b2e13c43934a219ed994505b259cf95fd09a1ad85db927c03b392fcc82a7f2445f0e41f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a7ce51764e56f70252ce41974e9c49bedbc88a5df00d926c3f126b3af5f7014682bb1dfe943453efde48a9288cebf0a1e54a059f9f02e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67fb20548f50e690eed211ae0afe8323c6a88e10dfb3f36a2c18dd4bc69f4ac2396f09b7a9dd4935633b3a119f778b39d109d370666418;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9de031945a3c401c4c7f7df0e549f410cd25e77c9f2ef587ec20f9763547fb78eed18d9e9e4aeb968e9cfcbbb327376d00aca58d1a7fd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6a6bf29d007dedbde43c89fdecc995ef848e3be1f8ffc98221dda5cbf4102c7c9b6d1c56071a453eb4339b81ce499cff693510c4ebd44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124c0347c06135ccbf63f8ce91ef2bb11bd9d40001a7883433c63f99e0ce2e6725729e01623b33c52087247e364126f2a5f82a694ead375;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2e35518ce40d217a19d60ecd233969590155818233d037d266cad37c66f72e8d75302ec91cba0589ee5b3eca626b1846a0f5622e96cc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16661c1dfe9cfd2e4e36158adb16a8b85db5bb2c83e92d30bae75886938ca41acb915850e20de812ff4cfb62e4ad8166a732a1f8c2a04fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1416d33205270cd64fdb84e90a709d65b03727134f1fd941c18862742f293a4f2bac6c4be52ffdc3c73abceace772777408ac7062b0202a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1119957a04b54cd1390ae788f53e167a4f12aa2ff8747e4473769a32c368fb79f6783f47c72646ba99674674fcea45dfcc8ace3a9ef3844;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca2e2bd3ff4ff720b519fadd4dc512e8579ced8466987dc34116cd73b259692b068997c7b116d657a00aa1667b7a2d24fefc3551ee337c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1691985e1fe972e8a18292bc93bca698aeb8d0daa59761eed72d75d03135668be52d9ba094306193d2b7fdc7cfc5762c50577c2c45f4695;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24e74a5eaba86d7dbd448c54f6ec5cab049b1e10b772e93df2813ac9c30266db98bced35a9fd1bbd9b3ab189a822a50951c8e7b643e732;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb96196ea6190e88ced0678e89add806f1f76ae373dbfcaf11c69097c578903db02398f2bbde2a6dab6fe37fa0293dbeaad8d958d17629;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7962283dfb602b1b979c1b8aaf156d1e0a070ff3917d3a7c2995979447cb4dc1c992c34a23dff33cc7f465172cadd60f3fb23d6429e88a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98adc68b2d372409fa57fbdc0ae32aa6aeef35e591028e3090b372daa0dbfa998f4f70deebb2f24cd209b19b0f09140dd027865d9172e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b06f097af44ef5137228ba1fe6d97662fb9b40564247919693ffec00b5233ac2bbfd8c13a0fb12a9c00b0da530b774053cc0ef83cbda71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c181417f4f80facca47d2f56c5d022f596dab222cbcf308c1aa642f35f69423e91e84944e2509fd86d72b782f9d9f33eb8a9d00772f56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c67147c1227bbf0e49c7d00f5749cf4734c5219a2590ee11499c26eaf32beb63405f7b913891cc6767b4edbad87f8aca5934a5a904cbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1041909c110fd8d0dd388e5e9fe4c680c9b604bb787afb40fd9e1f7fedf40f95c8e9518d5a0d7a0a0e257154be51b9753262da6d79f3276;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6dd395794609fbf4fa242de1f9b3f25a4269ab2a4486d4cf57a432f744d8e9b5422b447fbffd2dc95c5e68f0b534a17b918840c222e1bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1581cebdc38e11fc4285fd6513b320eaee2c06efc1e0a09155c805cb1056a4cd309e3ed6f8d3cf231e77fe7ecccd448f499ed5d1b101d70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h159bc9bea573f405643a09c8520eb9d9b4f10e3853dd6a4d856754507a0a346f1a816e7828528440c2d0f14be5fcf432006b0654d1c7e1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1fbadbabf5aa922da8108db2292632898c3c22e9d23f6f3001b7dc62922792f93567024730031b0842725c01f84edea9f0c3aaed48f11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde2a2926863e6048cf329b4ab6a845dd228825b9d83f725b9048bd16ea614bf25daa10f598e07f06733d1fd7f87b01c550b2c3472e4fd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c881d1d0f4935a3970f5c9576ff1aca2b26a5382b07391224b10125a8d8723ea4eaf40c5fd5729e0480b0aa1ee77d6b4e0abe0e633870d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d0cea37a77f0552287dd66dd6349a7804e65709eed98c8d96fdad3f1ffab4fd7f57bd7064398382f00b290a3edae9cb68306cdd6a79b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187726720b24c5dfbc042243bb1cff363bde8687554041b7391372fda5ce4f5fc828806b06894d59259ce70d1a7fcdb5576c165a21eaac9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dc992bd7e6fd8478339907ec6b4d228440cd33e63a1e101ca98c13de5e2389d2691193de4fab5abc40faa6678d39496a8a830da595342;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130c21d8b537a977123f80c6b08963ef9317207786ed459b32b326c637cf8302f5f5144335dd60ea5d074482f61a753b7bbfd5334f2d358;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15750ccef8bc653c8e22df8040a0dbeb54641623713d68bc129a2eb00af4216a1516ed30a114f305e021e1dced2a021c074d21acd56e7bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha533cf17aaa3d40f234bea25ef2cc3a1f1f8fe6d61762ecd74f6d6fc127f3f19d360132cedea8a097a66f9de53e913ac93acc2004fb683;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cb8e0ee1d10f2c24b06bf81331b03031c4316b47bc867ff72f8c75f538d1a43e411cc76541d62d6fa28d511befe793802643c1cd7b493;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd8c2682becad057e1f5c3e20b5ae5e861af3c6dd689bf17e8217241a8d81f8cec50f298bf54d774886b1ec725bd6631b4364875af9600;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146f50638690f8d5969ead55432d0e4ff0a379336458a1672f3b48696f2dfcf8df54f8ae120b31c6111b4287b3d47306d28e71bb80b9f9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7dc1b4f3e6ba17bb35ea088b87572c559af6bf01a71a8c1e810866023bc22139b85c4218e24be66acbb533be361ecfafa3ea4cafae4d94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9bed27eaca0ed627301d2dacec04c7de5f81c46f539d857d130dfe2cd6d79ed61c4649758f4c0d447a74bfba77cc44fbcc9b01c43bc61c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae5e3b65f332e8df37a4bcbba80a86c564fe4359d89ba0f5c969f9f699c9b0b03f575c4304f2ec52a8bb3a5330acddf850e69ec542cdc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36f015cb173d7858120d82e68d96e99461b4742a5baaf6b823c6fd3c6a6a682f7672f90986bec5b0e0fbdbd942b076bc7c4f199ccb6c35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h50eedf2d4c09809abc7f03a0d29b00fc2f8eddddb90cd196afce5a9202ac757ad8f49bb6675c39f65cc01aca7d06ce84f42b6b4f8ff48e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cff61ddd76473ad6b46b720141065660ec4f6a4148b2bef34a829c30f342a260d7c8c1c1e09e64de520ebafa620932e1d3a0311382aa9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1c2882f893a3d0193fea58eba8802f6d1f8ae9bd71176dfa470164368da6e7415573ec7cbb5f389998917011bbfcf99890576bde8d5a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a1a5e27213952c72f3f868bf7e3adef5a5c3f6afe7f8831c1913da8e2f23a742654d4b34434e4a49d57ff3316b1ad693584645df1cbe4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14999956db1112961116dd5920feceec91af5cc843f63fef9bbb27114e53e9f671d7faefeb0a9106c181d712600e569846805df0fc8804d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ebb83dca4ff4cd4809c236f3a856b14cd7f5d561b8e7c75e6b4b315b5372cde1ac7c7857bde109482e11ede6d4fa5713816ec19965bbd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ed3014c2b56b27f7e2c8edefc25f39c8a6a3684e3dba8da87f831b2652577c3e30680a1c1c9401707a851910c237d6052e330c62c18b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb1ce5288c1411e054d7b53e804e81456b6e0960bbe1aae47294a0c0c6e4db7f644d3c0252c1681ee1520e32d103f0c7e927915b85c1f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcc3af9b456785c0277c8be0c215670c84327db06d2bde9adf1052f15ac2078b651dfbfdd48b0de6806d70d9b03385093e6044d29e8a87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d79f8fceadad3d758a7b30c416ed213aa441bbdfe9bab2ded0353db3164f463bce2bd39940a33301fb77f08eb009cfa41a5915ca11d07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152854e84d94e8cb9e1bf8b16867e52f3d8ad4d57adc1b69f006ce663cbc65d6b02264e93ac895e4ee7252ed4ebf2cc87b5a67e5965e9f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80b45409dd0c7e50a48052bba277d59b48e10380bb1e9d04c3811e50a6f70032532efd7e8d0bf6b0dbd3e8770afb2723b0f0d3c69b877a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc86f478eab97b1003804142b108aa1c776554f37f0b07868da6656c365e76f944a02ca9630df6adfe2e4415a097119e2c0550df4122325;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdd75b1bf233ba7ae08ea41650ca33e4fb6efaa518fb4a187a3ebaa6520b8f3ec11cbcc23183cc789c57b1abc9fcf8aa1f15298cf4f300;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e6719659adcdf4d13f28994169223fd8f2ff82256007fc614cb66997bc6a126ddfa43fc829975752acc4ac2fce455edb4cd3d51a3fdf2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heeca7d0dd59ba032d5f25caa287ff1eaa8127e152ddf776e16d9cfa999d4d8b8695aebfdec3421e4571e27a103fa0e3167a5e61fd24e95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h258d40a337d4ac9b7d3a70f438d514cb7441b09103f599f01e21e11dddf96f94dbbc5f6961e413652e183aa197a73987d756ced33d5482;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c244dead3d0662b3d2eae59f4fdc8595c7fcd748543c5042201f4b2cecec572a813ea271471833d9ca9b7eb8131d3bfd40de1661b48ed3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hefb860a1cf69c058542e5e52fcd0a04390d6c8535b10dbacebb0bae9c0f29d8c59d864305050f9e1d76e975b50403cfb8053bcb983c9af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed9afd148de2e48cb29bb9de242027287da1177d946197c100ffa3f038346e31c4fad6175f026f7d956604df9cc3ed288fd0f78d377d73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h824b19261581d57b05f8969c28a7b063edabf8f7659e40aff1ce11ff320e930cdb6cbdc61190a8e76e030eeb7c0279eb3a75bca29f4abf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb15b9411885924897d8f3170a93818e9465b359791b5df6ad500e50eb61e8c46d2e679cfdffaf9c70f73942ef714809a4543dab8618a6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1505788606adc0df3e2ee7cde78f35480fab209f97d5ee5be79dc1da41a575df97f7441830c00fb239e9f4920e94541532bbc4d7e37229c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1269da583462f3eccb6b9cc14684195f686e63cc46420ea17361d7045088bbebf3d16ea954bc5ef36f16f5443bdc28caaa3262113cea60e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cd52c9cdce42dc63ff5cb8ded9136b9940e464ec7843226f733b646bdbd1b8ed6a7b4b451f4ac180eca737b15bae1acbc38e2c0bf786a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e40f088444cb429ab31b62a82a3140d65a5b30e9da7101cb2a87ab846cf7faa8753763464de94e9704ecb72405ffbae260128d9e1f732a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a8911823bd8e8401d2ad95e6c8b3dfc5d15a5670f938cacdc89d1fa3103a7bee44899eba3ee811d0b585eeae5b0c86da5a1c5aeea639f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bbc7b45bf780c6926fd874441338b8780b6eb0ab3f0df7a4b440bb75ae63faae7889fa31f31d62c2dc94a68d4114b543490d628dcbd5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58c4b8637d921c90127a9342a0fa9aa1694244027f415b14338a303231ef28a65488d580461d4c5e16e04ebfb55fffd1c03d2618cc24fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa3788605e757dd2de3a92a054384c64d30f8e22217be10f4cd36c426ac1fa8f273ae55daebf80bbfd3ae9dedc24b1978cec1b7adb7a47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c18bd4335d4a1572545f09ebc8640d7e613b773a83d3e54463f3c02da3ee2553da8673dab3669ad617459c6bef0a7842a21abd2410df57;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ce65a74a684984a17a25e3ebdd6e9cca8b53594ff9fed4322de01c8abf32aef7e080c2eee385e6609b02178e9a953b0802b95d640032e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a06a42dbff92260cac278be8da28bd3983f0216930f165364e44668e874857fab204e27a76951738cc68653b6f4d917ccdb043bd3aa6ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4fe284274c5417ae5a5df078252542269cd504c2cf6488a76b530227784f6114c25d112fbbeff479c2f4e1f5c5e63e0a2ede7afdabb4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1933f91c7901e47564ec5518d1c8793dd90246d86dd02ebd1bb5df55a7aadfd6f293cc3fceaa5dd0cea2658112ba39ec4321388828d3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hedacd9a80f77e4db5f475a0fc89a57cf012c40688fa71368841d12e8b0d72e2c116858e406542e270f3d5613f434e1c365d36d6dca1793;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e36b8c3609c31b7dc65748cfe5ac9af3c33105a135b76d27d7de9f43632b133f9abcb1eaf581d4c1eea7a42db7c393750ad2bd1636f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69ce06e0f25a5cf410668d489c849899aa3ce4b9a8f2fe377001da22004ca071fd1520085e71c9aeeeef7580dc568948a904904db3b2c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45d69bef6fec40a81ec32a0541ffe4ca50d50583c2b93ab0868cb176a9c5d1bcc5f718a7791dbf893f67aaa7ebc471d627804a067d0e12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcfddca1dc38274a0753f5a8154e1c1773dbbae81a53dd6deca7bf3785ac94977940aeed7d8dd343ebe57ffe3351761b5fa2638c4ef869;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f9ad22d05516c6645d6eddd674dee5a214eb7279ef705b049f9df3203275a2213d1dba3ace6d9c4ec75a34c7a5a19081241178c5a88a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce5e16580c6e8d576949ab4cb389248b6e4c2a10d6e7bf07eb6f025db4d8a1aacf1f1b0591aca6f916bfb89266f19bd23b372169610359;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc94acf6dff4068d9916dcfa1adef2ba569d28a14dc40f05e8d1b274b04cc225188e8a4a3f4bbb83c2857a7c9d429b8e05335ae1596786;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1500c7704ad4863d12caabcf203a3d76572ed16130428becf10dfbe6c59851859306f67ed8d61c7403597ec962a692c454ffe018da28f58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b71be41985108d515a43c49030dba6cb8dd99985f46dadbdbf0f12024cde0d878a576e812683f915e44aeddfb2f9fa571b36ba3f218e16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e8f7c745799907cfc51079b75f1f08853bad9dcb691b93b29522a0cfefbb6f058b51e31ce345da1ec2745581f6ad4048477177cabc2a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91cea6210926f01ad432a734089965ecdee92c5dc62af0b8e4ab52d3f7ac9499aaf1ee48822fa67d5643220d5319aede33b76541cc389;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a25b76bbe38ff88c9cbb087d5d6e40cc60abbc319cef1837665a8f18530bd01c7bb2a283e51798ef754170286493fcd313b22c1e049d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c513b3f4f1bfe3b9646f4d9b9d9406593cefd9b79bd4becda5516aef7d80e397d8b3bd87308328224fb0c6698065e7d8b6e4342ab44cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1173264276d53171a3a8be9f5addaba6ffb9315a182bd6fa0b9f53ba51d9c91e1780acd2fff21ce35c1f06e5ccd8d753fd10af48473bd8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a7c68b539406b8e2f44d10b6b62107358a49f2447c5f378f595b40457fd41acbdbc84db37c9539bca7f37fff60d357af76665476fae66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87e79952f22785447dd037da999621311c9f4fc27d78bd84247efa590d4eb0e85f32a34d0e92f9aa6a1c35633f47ff0f4335b52e4fe8ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c19a31b16e93b6418d2f07d7614f262b0ac81f2ee6c6d7c1afd369106364f72f49173274d916c8899781a323baa0c27cef3cb3fe3ebfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e9f00700bc37cd8a391045a5d950e4fe92644ce19d87033f6e3f9b093f9ab812043754995e060635054c9e605ae1dd5067d4125b12f9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79b1a04a10cacdd59077081ee59d2f6fe277d4027e469987432d2987e7cb2aedcd2403fc8d30bb74d846583ecc13e29b4047e3fd741680;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9893bb4720cf9e92a67a7a35275158e16790c70955f92c17d7711105124607dde16ff0854114e341ef374432dde1ce24939f0ef67bb6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h398d38ca9508bd4b0afe60b414e7e24ee1a434cf62631a3bcee384c810f1160893fdc7da42c5f6e0142ea52406277bf2692f9d0649b1bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14969f3cc881b5a251dea2973792914a4cbda8112ec09b668ce82a8bf69f4938ba34b3ff09cacfbf5925a6c67812e3ad67dfc3a2e28b36e;
        #1
        $finish();
    end
endmodule
