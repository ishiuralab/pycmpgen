module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [13:0] src15;
    reg [12:0] src16;
    reg [11:0] src17;
    reg [10:0] src18;
    reg [9:0] src19;
    reg [8:0] src20;
    reg [7:0] src21;
    reg [6:0] src22;
    reg [5:0] src23;
    reg [4:0] src24;
    reg [3:0] src25;
    reg [2:0] src26;
    reg [1:0] src27;
    reg [0:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3])<<25) + ((src26[0] + src26[1] + src26[2])<<26) + ((src27[0] + src27[1])<<27) + ((src28[0])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a937d5900bf43a9bcffa4b07b38f2ee7d385247b2fdcfb5ed728b64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172013d46ec94957ff566611503aef2b5a41fca0ce8c685b28f309b1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d20ecb444a6292c8abfeb22eb80e2508c96177db69d9f06e6d47c18e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a5aa52ed90bd62a080a0ad242b8ab964f24c847facec5f7dcdf93ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hefb047b7b3b93f0fc29986ef7aae44e594c202863e878a68e138a33f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1151e5c3ece08fcb2f9f0b06df36b2ce6f637df88cbecd10c0b8d71d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48130878ceb492ba9a065c2340a73707e6dadba9d540dd64aac07365;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac818638db002653b4ef39c1acb7678433539a2ff2ebf7badcc31ca5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f42a876c6da54e0a67360a077625e794304913e59f5639426c66e065;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11deb33944dffa966075568f215d0d94bb94f735929c69d07f990ba50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8238b1545fcff8c2432571335f0f842cba07c8cce2cb14d37c0c031;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0cb615918fb8ab31f0d5426468deda51026c0d4fa213e4c8860169a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f71187e81652ddafd9fe172fc95d93dcb19c8b41dc896b58bd0f635;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb1cdfffde07b8cfbc0d86dd49a678fce9c81c8869266d32a910f1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83dab6f0f527815cb67705ef9e1a9155a4066eed821149c3135098c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c559f433a95e8c77a517f7e484ac6e15fadf903417f16ef15e770ed2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc43aec7cd518663790f591e55be655087ba8d1d1fad3385d46719ded;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcefc0ddc04fcd784a88bd7ec3af57307e5e453458577d0d21a797ae5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a5d709df63d1cc10bfe56c093460569f844268a05940d62b7495bc7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b8683332314f11d4e75875431b1765b9903d1375a39e3cacc66e2e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23eb16103d3e9d732015dbeb6eb54b34f9a7562de67e236e783f4e2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7d437d87d6ec453c4da4c1c44f5093b22e662687057a3cf63f81c85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95737c50d2b5ec3ad3196d16213ab03d2b1636312d5a03a5feda0bd7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21d2b80ce8667c3babd79f17f6dc419f48c2d91ad6755187d992a867;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b24d29c9467578d9486dfd363cf193c91c9772bdc468741c2ce4713;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148a53e32dfa4468a11859cdf75af53b9938d37c6dd3ed80da7c79ada;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h527364f0d70f281529d61c8056eaa791d89746a80b2ff43e603fcf8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd06c35e632407d94f21e52a54f173061e3a9579b601459e5ff3ea705;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fec994e59b483cd8d0b2603a31626088b538da0734c8da55152e3e8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98cd1696d3fb7b631de01d9c2bcfee907e05b099792e0003a977c8e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ce62f0cb4a9a111ca17b4c20c350cec65634fc2c8fb5dff21fb0d50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cfec68bcb74539e51bffa6134b16505ad9d3d7e4d4742e4dc359d4d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbc620d10fc286f1b587bed7fc686a5b381a0e1eaef7db1e0fa1fcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h99e89f55ca9b545d4553a76db475b91064965aefd8e8248aad8a5e33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hce4f22d9408146242d1ff471dbfc64a3fa39b7d3306889112602caf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a62970e54d1201bb001acd5ab4c6b765cc3d048f64f2eb35b9b975d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a43dd4f383307f62235776e302bf7dd13b0914a1d00c8e991cdb1a3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a0b70702e2f57e6f2f76c83eae4f6e28313b3f8ed4ccdefa5f70b13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea3df3af021c3ae9ca32a9701047235c2f8afc3f30925da758bb186a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdab70523f6005712f059079ee4dfbe22f3c17554521ceaee7452cf00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h611262806f8e4509b24950cfcf3070165e268efb27336522a71cabc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62ff51c3c90ccda7d383d479b82e7ab40d1932c6e6e497e57774fea5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6409dbdf17a2fb37e439053241a19f9daed2ee766457dfb706c2a9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8813c9d44437fb0d42d93b531f27382bdb20f1c1d932a280566e7af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10efb5c3e8b224f628130506099203cc15356e9ff0877baf3257692b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70053060666f1d9421041678bb09ed6eb6b5e1b934466ac70e338a5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcabe7d31395016f34165926a91fe4b243ebf78d5acab403e85d74d05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h708f303099ebaba58e17f2cbbb40c8dce1bc6e28e0674e42e8d9a93c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h961206ea2061eef4a7dab29ee164d7ae28f4a31169a1f6c40e303952;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9100840b1a9cb9a56d6ff714f66439237a626e834754ae3cf52c8c93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1742f34886a633c61e2b14d9176b27beb019986a8a703e8340bc7d7f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a160a15d59d5ead4b86ccdb179a08800bd20f5d850a02ed02ca0960;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d64f9c4f03202780291921f6849e484d84ea906b094d4566630bb43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ca5fccbf298bb8706d9a1a3df789d54aec18d08e9c7875b9f6f5591;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45bc89c13e3d32bbc4c25e0a9996a0d89d091a280a000e325607d389;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91d6cfb6ffc26ed3f9c9a06b519c05b78e0382b87cf45fcd6665c814;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8628236a0edc66755660a0cd958c35a19396e4aaef5eb911ea6ca9ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddc2324b55dab22e7b6a4505e46edc0404f83db8dd06781a7c5a549c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cea56afc4d06a48e94197d4617540615d3c7332c77b3128500a0954e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1daacc698d912c37becd56504dc0036e5f1de8812e9f4f6c88782d47e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd6e232ca4bc90788656a7587d6373ba54c0721b3a1ce55ae1a89da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4708e7ca95c8ccf7ff4dec2d76f0ac363bbc4b3cf5f2c3fe257176d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e61d2abaaa627e048362854a5a7729f090d126488d135e0edd39c043;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f0f87c13cc1ca8ab16049e7f5667f72689e3993a690231e75986046;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1293acab2eaa23a6db75ba47b12256a09ed7915dd250c912e852f25f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h786ed138cb3ce8b9c8fdcdc3e1a3dff5881be59035ba32c79fbcc6f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd2f469bd928221fa042bc708ff2f2e6440020600867ad0711bbdb13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4790c2a124a0342c4eb6b146faed0533f921f904914496ac0c2d589b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ee47629604c0f121b3f148b005fe80b1f4568bee463e47951c91b99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142035a58adfb5b04ddce8b656b5642d951bd3c576b172bd569b9e57e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bfdf5ac1c6c14f4e210d230900e4ef41682f6100b46fe851021b08e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52071320e08f7b920eadc73af5181caa56c22ae302478fbf33d05a42;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h57dc56c00d3966df310a7cbbbc4cd9a7a2b46bbf8635ccb928e57c65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h118b779a302448d7fb9da89df0dda1af16548af0766ff586dc96a50cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb09ca9c396b9109161336f15791eb63fe3e6bb2931cde2f34d7697ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd1637f465ee197283e16d3772e4fc607898c2ed0dcd9faac34996d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb32ee29b9af2817b01ab0affabf39a347d99ec1812d70cbf7dcb5aa4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18326dab6805e5190b7dfab36358bf0084a5ee748c96710f760bded2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164d2536878c0671a2498f1930fd263d8c8c6e8e2407ff87cc6d15b37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1233b38999cca3ba3d36c46f21fb8d6dc438ff78d78400115bab768de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43eb2d6b3a30777b8a2f6dac9f086d73a8b297cce8f5ac7c9107a790;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb037b629bf4ae2c6a2ba00049368a20e11403ff90d7191ebb90786cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ba37a303630625c041508059f5794a71dddb00b090a9a4a1c81e990;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8463fdb5871ff62b00a05a2644d13cd4a8bf05ee1547932d2790d6d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37453206e9934c156e566c8105dfa71ebcc1b0b9c5bb055bd795e6ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf32df063d1dd3135c8405d3d5e2998a92175cbe5548e7d83b8128fac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111f6edb70b597578a8e8fba4c4239b583f3d6cdd737928de564de4f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f4c1399e2d3807e5575c31cbe9009264a22d278b795d2e8939842d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df0235a1653a63545928a408e56fde1dc8724ba508db5d0de58ef1aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h31332bf63a1439e0d8107175c432abe5f701161b894f4cbb2776e78e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16921bab1bcb282915871a78c329ae2e214329180446d3eaeb5b8fda2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd77c423a6e191df36124c2a5a438c01d44e39e3d850beb50759b6acf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24d3e29591d3872510862731aa88f252b7e15ffeae645232e15725fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a139455303cf898876d5900107ff38afc82a435522cfd759f69c8ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1de4a0e949e5ee65884b13a0deba27b92360d88f119d5eb288d79073c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40dd2ff525f2824651fa4cc24a3c723a9eaabee7ae032641e76f875a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1231c6d3d1d3fdf78a17bb8ccdfb8cf2251a98f23ca61ac1e74a80ece;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba60720de7760bcdc59a053e65094e71263eea2ad9245cfa2f986512;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4c571b1f7c6e445e7904c4288384e1bb4f2119ec06cca0dfb073dc5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7443e301140632b8bf956612e95e8328103ff23ba3bacdc23753460;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f303480535e33dba8fb5b377e7babc1a1166fd6b92867af9d183501;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21e01ed9ac712a6eade10974e78acfb484a4d2b9613e1269335d6826;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1487bd7b9580e4956b4d6b694ae335fde6c8ef62dcf44bbd00d77fdb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3de13497360685536eb205f0368e5d6db52f7cd92eeec71347707f35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h985c009f9b69b7600f920c51adde03234f051db47257864febad1e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11253d437e9be740431cf1b9162aa0fc5533226f64da6ab5e8b809f45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h722a5cccb7868f660540f6a63e05b87fc3dfe6fe2611d7f2ad2f04e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4246781249b5083721dfb6551712da44b68e788c953968e6cb739ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h67f35a49c105ccfd00f8d0c7e96e045fc3a32e06fe53173b013804f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53e8622eaee7fd07532bc00c47d748d030905076b137e26cb9635889;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc42a61591fe7da4885aaaf6885d00e02cabe6f56c1b9588f2003e639;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb5a1212231aa6a44135bd101e8aa82b398996dffbd7f7754d2b63726;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194fb2082dcc8d037a743f78032ac4819dbf048c504125dae2dc4fe19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58878b00762352bfdf11af53b1fbb911e575358359ce64e43684dd53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb27c93ddf1a4a6ab194f6ff2649bfc468f57b59fbece55d78c69e120;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d545f0e367b449dbff61d62ac19d5f2b7cbe0f86a37cdedaddbeaf13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3f13b7d2352f4d2ae8089de7b62c84c543321352ab84a1fcc349a8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51d0bc313384fa1586b4971a69a820d7518fe12ea51880af4d8b8c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h145fdfa0e08066ec81317197ddf7e7dc208b20f67855c6311684c8b79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7fd115437ee55521046db3246c3eb7fecbf7266f58b37e7308121c94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125753f35e54347e3c26645497e7a69a55d4d70ed17e1634e18cc5fd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h852cc2f5631079c3fd3a0fe4c6d46a507b814098ae6550d57c743b8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108828ce94388394049944578b93f59024d06fae38fe874435ccb6ad8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78aecac56c176e3bb165cb6bb0281f1137dcf0690b974e50ccf46a68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff52429a18ca4477099df481cc894d06ea63823ee355af4e9564b341;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he862060a54d9435c80fadc2b62cee2e05e85905db91fad591d2badb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf1b0f9ed0c049107dc0efe4a49d7ef3bbd52c16511dd4fa9e0b735d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6040607665452c66e53954058fc5b0a5a5e7246a693386f323c6536;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53a79a558651e4eaef186b1efd619752349f31898594e25b0ad27434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23ccb2db0b8756ba72a46bcfcae7207999fe4e4aa962a05b17dd01e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18aa8287814a5b977f84af3cda6fa613543d997c12bf683b899b93364;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbbffe95722b9f486d3630cf31a5f19c5513aefdbc18993f4e587760;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha61649f5f4919d77f25d7cdda28c678c30c546525ee335f65d615548;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190610f1908b8027bb5a84631b13e54e98ba1e48ac6aaa10a0a80126e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da298817843d5814e7bcfcf1ed543774e019e648d28ee331ca50c7c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f1d0d9a847e15404eb9cb48f17ac08023e42f8501c543ee7de6bfee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa08697379863a37b7aa111b771885d0ddfe4d6d77bcfb07fecfd047;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h46e9b9a8f958db51d6e15e9255d578190dc92b10867c4e7f1eda3967;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c99e2c31d9949843a83ef510ffe013072d2b2873ecd84f718fd6b9ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb6cd980131159fd6d74a64ecc96b49394e94db3228ef4b5381f4c2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd366665ed8fd415577df137bbc2d2046fa853233cdfbf4ac9fb9ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9b7ff7ece3dd4d20f671945b0f1bbdd76a4b9fc004cc2fd4c5bd8ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha813b224ced8258d6024b595eb7229cc39e20aafc94421836ccf3c70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c0fda65f67db3fe95058c8d7d4788d64e0faedb37df19133106a10f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb09da62702c22712f7ba6813231eaa71778941c24786e370ee0b00a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e086b1b5f4c6b6bf858be1ae00bd3f78f623a611e7692e5838267b0c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h760417f56de2416d2d7aed12fae30fa0183bf1033813bcf27305c89b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee3a081b368eae2899bc02cdd24d2baee388b60e97f01c0b8fe512f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb04cd2d4881423a5a1981a97d7a89c7e8d08c87b35097d133d5d48af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12cd4d98ef92ad74db80b89dc2eaae5aa2683c43c74b6e95c61f27961;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b0057a6b7fea757cb41a5065d967e97e2a2c8ae1a072281e4e174f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a482f1cd5e8becb44511e154c6c7d3c7992ef34a1f2d9e70aa76952;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0a508915bec670c0a97dfd88723ff8c38d34ef3954fb3f601e5d41b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17cd135a765da9c9fa20e969f4b86946ce8fb222cc1b3fed830d500f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15519096b9e7fc962e99c691aae1c05aaee03051edef20b153b691736;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddfc4e2f6607fe7a555325d133367a8697a6af50916a616222ad1e93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1211dbf685dac307cac1879d8184d94ed18c84a20b6aa5bd46d3f97c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136fbfa15e88c30534bac639525026e1b69eb76b76c11c20eb38112b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150257899675dd7adf3afb62c88486a0b3851249d8090ce61b9b0ddbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h112527db5348038e3611458a4af4d724227676ca113c5c3405a7606ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9e96d82b7a7fb8096c9c226a2ec08ab0b5815d5403be23baee7dc7cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fe7ca44b97528b09cb8f4aab660e0ac3c1f9ed17c2f051cc7fa3b99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a9580408cad12ca3192dccbbffe8f7bd817c8d4461c7e353b2c40af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2016735fa46f7b945437868527d4996c453d400f22409a450405d3dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5b7014aaa05efa8487fc7abce3acf61a535293b32cc79ef43c99367d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe7869a103275bff4cd78da785ca01d47189343219223f78265b839;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120f3da42baf2cf77951c0cd232f52a0fb18dc755707936f0869321f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195ea476961238e8a667d5833737b1af43c60c1cb4a6520ae9e33f567;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f9e039dc90b43075c3063813e891d37b89c842d3c656babc692dae1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c1df3131b868ab7e429fd73b5063302a08340bfe695ad5a8ebb49f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae964eb61ba9be1110f1ca7cb3666c69d5244725c50936d63d967ff4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18afff34fa945b3a79288dde1a57ea6e73bd5e1d874885cf63f2913c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd452869dc21876971fe809a6849a981d5666d6d7ef40bf18760578c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc792bf37d482280f3a01085ca1c955b35c0cdac8c6e884d38fd2f24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1367b9b491e5f67bd30094bdc24dee05d9f81aa1f754b2cba2220ba9d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184b5ec4f25071460f6dc5db492796032ad79865147876970cee90d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5877218b022e3c13495028400857c903f670488b9ae686572915d330;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1854af15e520baa099e5e0800af56881dbf1e4f9fbb1a0058ac4773a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ae5120aa76c9e13a922781b6785d8e9b896bbb36c43ec9308d2cd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef69afe807234594fa757a4f3e907a7c95effd97a0c7596a28bd1a41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df869ea7e1bdc176b5d0a4ace3b8e700a7206712178d62f595968635;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c2e575e4e949e671ccaf4ec05c6bede6fdd3fce89900bfcd0423c83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8c4f428bf1c649fe4933c25ee8cee011996e4ca50870ab5583a56fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee1fdada956bb517c7cb683820601b84f4edc94baf2755875582290;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d1e148b2a5987634e7f6285bb520d966b25d511c2bbf131c4c42fc68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdcf795677e307118aee5b6fda54321c9822fc5b542a16a108142c849;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df920f137388719d2ec9470a92a0087f7582416392733ca84ffe930b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f0b9b61b8ef98916704ca4283d2c6b6da53d543fb3f26f1825682aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7856b6ba1e7f6afd9ee97fd7758fc8c8cb20143fcb64106819a694e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21f77446edd4a291c805522be160edb431422f06fe043edbae4460ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0c55e5aca152377eae4cd031b61f21f50e9438eec66ec29c3c6d0fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4db916a9e96939d368d5c940134b50e6d7d3b4359da4e48fe35d4544;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf45c3431f112e44b3d70142721ec2f8fbf8bc792f3c46877562f4df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h946106deb0e98bddcc3406e90c48abd6c9b50514479c6e83cd7e3c12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12561e36bc7cca43a53bfb192953bc084b0e816b6d5979bd3e16b03a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcfe5b10521b94acff25d1b21f16905be4d110ef8e69bc19e648b6ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd162b76b4f604ca841b8f4814a6d36bb23b3e1f84758d88b3bffd04f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e8d61dafa15aab2806a001afdef0561931bbbf117fb8010f60f2dde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105e46ccf66fa4b4df293924226dedabcd9d1d83482291c357d2585d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2287a5ae2f34ceb97524a7843554bd5e450d509fffddb7e4aac8203;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h899bb2e6591ded12cedbc1bc7daa1e2968a96beec1dc15f72c513f8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha431207d79aa55942dd3a51374db1a1361075b12034fde0c74597815;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d3051169481158a557a616ce03811a4f6fe4b34acc57583e35c878c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5202610660752ac38ef485f108b2bbd94629abbf6fdead8dd70640d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f82d1d53bb1fc20d94df8ce945f17a6dbcea7940b24492d88212d24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb10a2e4e233e3338e0e1563ef87b6477094b0197e7d03e0230d2c03f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f1c8a2c51f5ee22511a6d9bc788ebfc3f11de0a7eef0d28647605b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hedb6e7fe5cd2849e2c84e0bb9a8186641aec88049312520e3e61dc0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4561fe373ff57d3e3434065af162d033ac60b60ea1de60d31ac42e27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131e9d238571f9d44111683f3edfa8c88f16b6d635005736d05cf6cf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a701bb849e888c6feac9e74a59c3c338b9ea3ab7e26c9579c33828ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1955db818822040b5ea40399ce5a822023fb385a13143eba5e26fb054;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he48e89a275b4cfdd6860f41734a2680d47a507a04957f25606474cf9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d1f666243fbc5cdf1d1966a1a162e0066bf68cefe6840de768f57c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a92794a3d5721fbef09fdcb977f365fc1a8695cb3e35c66705f761c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a2e59e10ef6fd38ec7b66c2ef7066916251f84f7383d84d55f75426;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc99f1c66d13c9b84b6ef288553e84c105076e33b625de985c94f3bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h149cad010a7231e73e291a204d39a2f0e9e863c49a3d480d67f61f795;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h112987da415065608affa0a93bd30add24a3f1203a4a6017ef1dafb4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fb7944f59916b0d55ad26052caab7579fd48c29ed297c4da0bf8325;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce754e7fafa7aaecc265c3836857dff9b1a9acadbe2040487a2c9832;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ddec5b4566a3535b9ec00eb2baa2469e6cfd91d529cb8594a3d92b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7afb7a971df1fa8a15c307111b5c477ec2728ea712767ca35c0e292d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a75f83461e7c904ac80272ab07c1de0d769e7b8efc0a977c73b7f410;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b0a32b623c924b25ccc73b6247bb7f2875f18fdb1fe093466610207;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f5a2e84b56627cc0300c9ccd7cd392411be1e03613d0925ac535ca7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9763463fbbea2ad31253bb3c2a618d3ea37882954e0372ddfc6926c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h124389d91da8aa015d5eb2938dea559b4968420e01ade3fc1424c3dc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h338b1bb4200ead9035eb3941cd52262a5c3da476cd8d8d23ef02686a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef740ef760ee552e8818bb63912916b5260721df5c7c0f58413c91aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h99730789b547c169ac1972fbec8722a2e638f0f81349d201d77dbde1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b2dfdd25db2ab3d5b2ef11783d35094c09cf81dc7d0337715fa36c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc009f1c9f54c3a5f161cd910c4de2d154b914de7cce8649235389918;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171ab6618c5cf461c84be59f0a8e7cce9aa5e397fe56767f4af85ac53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he2f7d94ceac1c45ab3a89c43a3feb25cb54fca34ff076b8a1e4e271b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17be7f402702e79be719a09fbadce5cd52579dcf63c3d7e9b6452040c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4b5d6773bd9b3cc850cc02e5d2b1d981a0cbaf1a575540aff48afd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43d0dcb1040183a34a44ef2fc2e3575b3ed43c99cf24d0cc7541d265;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a948c37558def362fceaa5d6539539515d9ec1831adbe4424ea04ea2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192e4548022fcdeef7ab25a58cebce4bc79abc18f0e854e107d90ce67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7e367a4ff18f6c3322d539c4cb426ec4ce7846a8dbd7c237f7121f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e383fc42c6d38a56b0a800250e2854b362d66109d2007ca26260c09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168861bb376f793cd132c32617f0060a6ae901df92770331bf195668b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c32d80b9a1ad236a552e2bbbc048a3feb416d056241eced53c7bcae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4bbe8e8caafaa007d5b9caebf80b56a6c2a9f6cde8ab1bdfaf373d5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h149d9c45d9cec3db3cf6cf7734ab12d03b0aa32399e0806f45e995f94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h57471f6f3295e2c724ae686f9aa4d71d81e877b0aca7e33ff6041200;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74a25ef8bd60800dff7a1beae911f7733bbb1c443410d0740d3b1193;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c014215f6e85930d0f4af7b615c1f728d3394d0e77a7cbd36221de2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2194a18cfb88a39c898a5fec3414531c633efcf3e3faee24655b8c29;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda2c3c3a1091feceb61d2f210ddbff3fecb5cf4edfa501f304a9530d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbd8908107d0a17ed0c18adc5569776ac41461e5b86f199c8c73b9d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc409c036b5523ebabe80e47fd6ae049af3587ab33fde0ee23743817c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d5f09a40d36c056470067d5bb24386a14685843a623a6b199a143e10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da1be924b56d95dee74a1ac486e6dd00d49a8aec2a2d8a3c0564feab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h107569920d0d488ffbc5905f5f416f5c0a95f8209d4ba0d0d12a2fdf8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c822e3ed264b37ccdcceed3bf5c7d5a434ec2a67e1d988db19519f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb209240bd44d531a2e8c13f056d0fe78d360d86fb85a4fcf849933c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fc57ff6f3e22c5684c87fb250231f2f7a194866bf08507ac5401343;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1181857d7b812b4a18b0dcf1911c7bbcfc1d7fec1cb5b17d503c9b10c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b33096740da75c1ee2f3835d11cf46e6cc1149e21bf7df26273b707;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b0b6c4c0fc5d47a0b39fa5c13909b038de89732de790c3a2d2e2c4d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5c5c8f5b036540646caf6309206ac84b9202337ddd45eb114b0989f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a42bf74064fcbd9baf8f1a0b41fb6850f580604db637bffec752d961;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h296d7e1e435321a74bd7d3f4e4ee740cac2eec604fb42b1abe67aa59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da144df5e4301d1653a1b125147ab2580ff09f05914565975dec405;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d19641a03aa432a5dacede1300234c96a36151c57d0e226bef8a1a5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e901ba9013c66568f289c36806adb189e69cd3c62b1fce7ef2e16c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10041399ea7885b7b896eb8f8e68aa4082d0a647462c8b95d213a6882;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16dbd1ad11683aeb723d17ff84d993874a49a0833d2dddd9a653f00f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d7fa0618402f94399ff3ce22999693cb226d310eeb8089b2a4d89f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea7e85e32605626ad63dc2d56bae3dfb47c379a0e98f2e1c582f9882;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d128c64e75ced7d733a33f82533cce3c9618ad04fde5c47d2253a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2e2f574f04c189b632474aa7256af79131e552a719cfcb017717639;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1337f815218ebb5daae9fe5a569ffdaab87bcd55f816ee726dd8377de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h197e0440c6b60a9b239763dab990e74876dc08702b03b2caca5d73ff3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51735059c079df5e26d8a89c9847822f49e96649fa52b6e45736cbd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e2c124d585ad405c66f1a6f576f2dae8a4817aeb0f969dc01455fd1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habd0d353c4031fd69c166068750fd70d0da261be044abf53cb32789b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7d1bcb2f53dc6796d46efe88f78c4772294ed08c055f67dbe6ffc51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f024a7d65917e8bf82646eb32045ef2b59ce34194381fa4b1cecd046;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5eb957921f1efe70cca97c5bf4a1f1396a90268cf4feb48ab536b312;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1904fa2a254a175833e621d6aa86e58e26b586c86c83cd876e930320c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172f0921500f43db24dc266ca0012a8324f4c270c6f8d097a683eb664;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f728509c572715f67182cb30490a0192ae95fa451fc6811666d240c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6d96179453247f72b407b1d0b6cafae7b5979dd41a24f6d6bd1ff47e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d74a4ee8202eaa22d102dc23030903b91b453a0dcdcb13949ffbf8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he40e357102eceacc6be2906b676e62cb1576ff9b65bd5176d4d1e1d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a6744cfc3b18122267a152ae2933a4690b0bf70a7327940c8d13d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce4f524b60382f6b70bd235faa3d20651d893658bd69d95f9d0d4ef0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190a325461d009e0ac1ffecd76c0556d9a1fd1cd0a88a5d379c5102b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e0fe2ec765232f02a8686f4fb5ffb85de4bef312d63407091197e44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8ddad3fdba909c088ab27fa2dd53d69234e1559194f14598dacc30d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5fdeea928674a3afc39fa5951377f5152632bbcc272176cca419f53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d5a4340d7d0f45d8d0adb4598be1d54669f25a49d847773ca85e5eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b62244327944d1e206c33671454f663e1a3d898def0fc61b31998e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f2eda12064270b55b8791f07206ff69b708562bdc4b16aa18aba3a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2b8ad3933e2cd1cd24fb3c62dfcafaa5260fab655e5da11e5074d19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h27f87f1105d9cc1b77d00f903413493838b658565386ea4f7ef666ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha67ef63b1021af694b2a7c12f5174ada1d7de2f3d50f2c093de42ee6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176056a78bd5eebf32bf378a2b38df320383c1fca5b868e973502b42f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c7151df5c0f1590bb0701c249b1001558c245be1ddda432e461eb8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5359e6183bf7774c3eb8e56e40a86ad8ec194ff766611302986591ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a2b22c60b2d4e8257d1692e03bfcad416f20f9652176f74766a506a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6ae06b59b1a2046a83af9274de4aa540d003252d87aa36a7b5bcd53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1532325a47dca5b1d507f6c8ce0a1e8175923be108b557195083fff8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6f80714d5650fd5e870a856713f895679e74ee7a9ea19f00d873461;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21dd6d7600523256f1ec49ff4cc02431a7235db00c4a090ec80ef525;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha2e1580a6b81970fa3ccbf5e746bd1be77550c1075a051163349b56c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d36cb9d47fbf0fed061d2c14dc8e3d2b14bf6e9310dda45902f8e01f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188e7772bddefc0393f81cd3a08e92cbad4a8c4fb19a87eb5d0a7ed4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a54c13d19035f828c09d8fb445615eff9a968346508042cbd264aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf97a85f2272de7b640e20638be8b624e4b590f9f2064f30d345c11fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8151c632d80175198955b05e2b1c8fc2a443aaa8c18df1e8595cc43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d9b627d631706b163926fdd9b2f902366d3362df9404a16f71f36f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1548010d23f841369998ad5b8c5f5b2108f81c7c4673e2b293b27dd17;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13058214cde5cf2883832bce5c7518f030fe1fb7bbbe14aef1b782757;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1069d4d6d3cc354055aa5777fbc70c7413f132b2f06afaafb3a339693;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b506ef4b7a2d39d9768e54c0ccab8beabb9fe8129a5c8a307bd67b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a80d16da998e61eff54a1782417b3bcba94ab8c130afaede6650123;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf8783479b965ca6dd4651eb47a1d4d0fdf3fb1472122ef32bf0152e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5190f472d0a3815143f22570b5f5d67b415dcfbbdc4571e9930f8b49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ac1fdabaa32031dc9df7464a07f8c0e429a513009a883607e077065;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141d68051f4a772ddce4c40e9ba9ef85e3298ffb8e242ec00b248ad42;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e372d45b4bebcc2826e6d3d41e80aa23732e34286644c6a39926810;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h180d2a2f33787fefefaa1d5a698fc855152fd9f04e88819929e85d2e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h87620a699be40ce33206dd3da651a39a4f239a113465bde9c50e351b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18aa54a990021a42ef923d4e8fa8ac9175aceb504d0138fe3175bde14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a5b2110aaa89fe684b293869a61b8d4b8f651ae7624caedc654f9a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2aff3033c4f551866ebbe7390ff14aea43acbaeb855b6406f2badb33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6ae04eb7b061480d98eafa9401e6c4ded05fab2af1590f6641a2907;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4e67b1d1bbd1091a2c4b41f571f1f75a3bf10233a9f4991ec26bdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1440c5013cf9f7e6ac9e1b286846bee14ee83bd41d4f271781e46cfe6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1bee7273a2e8f08c652cf1ceb9bf12561bb817b5c61cd24b80ac7c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf820df9edc7f8d132176e5218813d52c3be533fe99207128723fb593;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf593915b49f538cb77171cd973129a501cc1782c74a01795cc41bb36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h945d7ed8b93b74aebea81eb006cce3618e5ce1654e782fcec356b8d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f66e7b120a3d56ed4556c0695d225dfe87dd5ca7272f720bed718749;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e09202696e1058d8cbcde1db42d3a0959c4420b6cebc7ee0d99b6827;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108b4245ebd5cfdb9d423a1352203f5282c9bbc3b31e198d1de9e6b15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c9cd59083fbf4b57e60e00f7f3d8a2982fb91c08090266777dd3b6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119d0a57b9617d4ef0af4e612f1ee0b987c398d0da2ca68e032861a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habd677d375f865910a03b3ac4db11a9e54e85cd7f604958e64ec3cc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d921b3dee0d53e7268b833265c24beb1009764f9bdfec89f4a126fe1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h84faa054dfebcbae6fa437c45563f446ab150a58d93cd97e7023389;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9327e4d80f404c1688792e9f6825a7527f38317a71461fe501bc5f91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b3762d4630db4d485a8ef95329ae7edbac3d2d433000d70be0c0db2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189b641ddde5ff0de1534d7a9dd0a3c93f4d79df9b3f77534af149176;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca386e9b84f9d40ebeaabc4c1307194796c8a85b3c38c9c2fda5ebfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6f332561fa1fa33397c737bec2b36fd6df4cd9145d5d8ebf1b1e11e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h550f0d67e8a49938383fec14d2ac2d0ca867fdb6ea56ac21f6969f79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ae8b3b0d90b6e862f8827f2b2c4d6bea9d681e8046b778ba5f12f2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd424fd80c8e48951abc25d18969831c4073c0b490072d63f381a53c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d779a97b0b28e4c0fd6497321d3e42f9e985ff1bd9567dff0f009ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd40a5dd6a25514f3077eda652eac559e6ae42ddda026a18804c6e183;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a421e0b3880a0764a26b752a3132c14db1cdf066fbd17c6e2b76a81d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152173a72dd35c0a9436c3ffcd0e94d1c14e197b4e2162d11c3693698;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98a072f47e5722961dabefee82af49433165cd1682390e8faf384a1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h116c47b0cd711130b9dc020e6ef21fea6b6e9f7f20c45fc2cb7973c13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h99f78dfb3e61d7e34dd180639e11b44e220efd5a78b71fd17e2357e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b8f8df1e4b4fd7e4c6d68b732987a8426fae34f2864ea2a07fd1878;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81d34b0b378a19e24929e1e628b0e2de5c8cba2a5d8dbff50d131e8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7928424a6c412950a587c8751bf01d6bb45e27a1308081ac6f33330;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ab3beccc511a02641f08d1f05482947fb8b143b6ef05bd9d31b09e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d31919f1ff7d8cf854b5b1565b3b49ed2f5e13fe1c9a28ee535dbdbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e34a4ad35465fe8badb33bf97def3ee8af605c81ec76f1179f191bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd550639b02467796abc6c3fa2c5a4ee33096842dc17fa194e529a65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff6c27bf72bbf799467303bbd7ceb84708762f9cc3d68ff5298b2116;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b3e37c3fc7ecb7c0cfa631af6abb4350e95e2237845ec0a7f86f279;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h31e38ad1f446be6295cef875473a6a47d6fc59881b242af1c55d1164;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1982eb79f932789f129fdfb06e956ee2a12fa57796094a9357814aff3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b5561d4d5da291b95772dc7f7291acfb9461bee455375a674d96a87;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b916f99d4c51c1b272bf0795d49a858a317227cdf5cc233dd707558;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df6a725024119afb3d255d3f9112338896d5b3d397a23c61f123fad7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b5e05a0b01ed72d746e96e470273b66b9e409ed299bb836831979b45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2150fc55ed2ff860f2db40e5a92171be7978ac30c498d4fc73c232c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1faf73fb1d2af895eea2e5a6b99d786de3f5ac72a9668e860dfdd49b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h754881e029a2af6ab48873a8ee8345461fe672f52dae9e3521db0084;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d8550993de35c96e222c7f37c2efde36cae9e404a4bd2103019412;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17aa5610f0231031f3498e58da2f230db443c8c52ac7bfd88073f26b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1353548c6b30f20e01c3ca9b61e398653f2f8a0a790b127c14dceaef0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1026bfb13d0322448d9cd19e27bd6f045a782dbb5253c0fb32a949071;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b1ef9223f337529334a0b02c9194b76c65d0871e74a653e7ec15745;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9485433fb5415045fdd5d8ecde4fc25179a5830d4b2e3f88d4dfe168;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda82581200afe2d72f2772ad48650804ed17256cab79ca5be294a08b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb524d1ac63adedb4ee9f63549ec91081b9d057b347e19b070b0f4b4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e2f677ac902c7e615a03704846e01f67927a9847a08ef5eb5634e19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172ab35d85c9a8d77680a74a4d719dc7af71cac08291497aa919fa424;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14be5884e20a15e1b9e5dd2af2e964efd4a2bcfa4768d25e8b5d62525;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ec8db352f9697d2291a5b63cbd9c19c520790a220e820e299926d0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa1d5a0a9e7a0ac125e02900855f764653052363def35619a8b5ac73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17db68d9a8fb016aef1b1870ac6a7c83e2f668a5ae4bb5fbe5205f181;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a940a9b35285e63640cf1158f2dbab79aefc27156d1e8ba27348ff5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1383535a3e424efe3ad8fb27d3677bb7e20be37780f1772c3a3acb0e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32859f7563ef9a61dc9a3b3da7d4cfdda08d3ca8d9a447fb1b378510;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc72027dad357591f51cbd8dfa83aebdcd249c12b912d22e607a85639;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c9c20c752bcb74108e2d1f0e5c12362ae1cba8bb25b98f7363845da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52bb4f0b18e25ed4cc836a78ec54dfabcd282fb800b9e29b89030a35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137a0bfe1ac21e30d83a9744a21b4bd09a9df4d0c10b51ce561b948b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecb825465d3c8e6fbcd04c11851eb8f62e805fd590662b3fe8171bc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hceadfe900266a4a96d0580298618b4e89d1ad7a1a5c02d59f5894a43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cef14c19e83582ed7d919c903a3e85aacc2e26fff7da7794139204ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1beb47f1a74bd403e947241d8e23ab8fde39962945ffc09b685fa20f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16eb3c474b8a7ffa4551774918d4dd4188051a890f6252f674f896f60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb0f5ee1faf66552fa521984c61e3c6a91ba8a29f6a3ba0d54c486bd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d53fbc1af457f09189be6afb805adc34f8d16e39cab2fe0945d3057;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ea5d1717e453a9b1c38183f54e6e6856d8e4cc275670df8fdfd84c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5dbc2453ae42b591e37aa9e6370e581b2d52a1ec02e6860a9877aba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h662d85fc7cd849f830e1e9959ef810d838b841ac54a1297c27c846d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f8b73673ff204356df8fc4442148e9047379b2a0a0db2b28e516722;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0ae000205456ea78bfee30ae9898c90c652792e499b394a5e832f99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0201a50757883f4b5a44ab674b27d740ac6b1ab631636b15824199;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86f67e642e0021c5ecd125ef24f136886bc8b5dd355db7b6ab1d5245;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b9d0a619682b075b6f95a011e88accc46e4763c5be1098f9a16dd06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h158f8d09f3e1984c5483f729e0ccd08a416d98691d305a69ed6d963a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117fdad998b241089b2f79e229fc3192d29034fa3807a7ba1010bf851;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9901a62b206d188567414de1b0b1481ae544dc2ada6357a560be08b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdaa71e80bdbbf571d5ace397b9967ae502d85f7f555076a0fe54848a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10d079a78a142c07d86e197b9a9d322fadcbfdc0a9deb5d187b4ad73b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4cc3d3c13e16ebf60d8bb3ddead363c9ec1cd5ed5e09622e5ad56db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c9c29fb1afb47f2f75235f280d764c7cafffa1ab2db6e930751ae73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63d14ee22b8587cfa01b4d08c34770baa9313869aac360e57c0bc7c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h50a94e68664ce35234b77c279bad7b223a3bd86e841034a2144dd665;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17aba34b6a207f58884e6a9c4da5b7259b8f7bb724eb4a922a5db9e27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1478bd62fbd295c4d87cc127f17fc96f0de9f5a722780c1da0183667f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1040f43ed6775a3e5c1d8eb299dea4c6d062252d08fac5cec8e1f5e87;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5dd7bd27369743e803a2e297f138c338613c6f4d5d75150bdd19b0f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd53c52b285354e907313fc92b0e32975406805b492fb8637a5b66ece;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfcd159cc54353548fa1e040d0ef406ca2661434d771c35ad1888a2c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f934bc7d943deedb572c7b12ba372ede72847a149009e9ee71cabebf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc56a0087cb3e9797c181c0cc6ace691b39473eb0d9c8d5af9237c54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h655ea2f7b581462a83b1814a39cc7fb0881cb1ede076d37a1b5e421f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f93fc8fa7361796e52765eaea0bc3a9eec077afa4df358f0218634b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b280a36903b7f8c5a90bc050bf4633cd16d659f7a91f08a245f5238;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he66a3185c9c640df6054fdcbf5938f6059b49f41b549a7390d2dcc79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49f87b3e43bdd2018f3eb089bed85809ca85e0e5e29abf2f1caab698;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e57e3c48eed3e178c157a7c807d17ce4fc7f8e4623b71874244dbcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13266b484b2bea075860ed32d378d3a1f9b37bf3d971d69ea6b6d10e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1006cc97d15626e1a577fe345bf6ad2382438ffea64cf652a717479d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1adb2849c5d543fa3a717c33f3d8b2535b6c98d10245a63f8d657828b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152c7837263b367156f057cc14313b2d1b4200ff48bf1e8ff602970b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e9fef7a51ce57b8deb5f6fbc62375d205d434778597148c5ba253ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h197f0573fbccc3a3ef2daa6524bb50bbdf38e1565e6487268e70c7fb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hca32f0226d6bec156cf7e949ed70166d4c30b19aa5e8f83df2896fcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1446c5e87a953d70deecb5fd8c67b83f013ecc5a3b845c1329eca5afe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd1b6064bc8cc2aa5ef861a0aba4f571dfbdf6afbd93b78513aeac07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137804442627ba02fa26de55f762cae064d4c1a217892623d676b0bcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4c81802d2ae49f4830a6fd92c1386fad8599fac01006dd8d39ecd9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13890174025c670f6311f7c05a78282cb7771bbb6b418bf2e56acf656;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194f2fd67687113d8513ba134e33c96eca7c1bdc29464dbd6b4f094c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1e823b187f19e2386101728c8304b2cc82ed86d4607b408a4115f52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7cb2705e60a88d5cfed2cc274c7143aee6d16b66af759bd16e34953;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13896d6fe2bc35627fbf73718521caa3fa1b69568daa50f83bf5b68a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194c4d9fa25ceca7e23780b3b9154d79be172938692af2308c63c30df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h470d05dbebb7c62cda7becce48064a94676775352cbe66dd13711b3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150f733e572f7eb009d9c2cd60975dd56b992a4ea4d65d4b3ad1f59ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d693b9c463159193c9adcf4dc7eef7ca2afb520a5e732332cc9fa6d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb4ea281c99fb1c5126362dc6cb828096b1a5c3e2b47b8b3c1ba027fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92048abc35541874ab7923ce61b3110ce444ab311d85d55751df3d37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda49db1b1f1b7587b89d90314f05d95ca25d44f6b92a69ef82fa5872;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181ef34bb57b18a368f0c33d8f835d941df95a6747b9d56eab73c18f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c5afc9e8c8d2a5b70c793c9d76b255f17ac2a0ce2e07928b804bbaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1247a9172a9d6c245d282df423d29a728fac96d7e6f0a1c1f2052f075;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1c01dd40720981c1d734e2b3bfcfa11251e4ab082648429bb9f1e04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b23e3831e932ec97b65968edd5bc65a4d5fa921f22c236360e844d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he699d9dbf1ab3e35a229caadfa7a85d7ed39662bb9c9694b3335e905;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9157dbf5a9d9ef12099532212d48efa951197619e33bf68d11161569;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e0874d68229c3830bb85fd1abee76c7526639dd04f19b68886112fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cdf4fd124f39ecee05120513baf10b834a187911bdb38ab06ed065e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79dfc216a91c593904b9ba5863f155a9d76d8a4c26e4bbc3031a1666;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df4f862a7603952a4c9c6820107ba486f7edd1c0a6a20458a0f8ba5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a15dc0ed1c27528083c27ebf5c8a8de81591219fc02249b56b33f90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc2a03e467cbd5c0790d31706584574efe10c9bcb3a2c45755b24567;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h27157580fe58ae96b00c42b78fdbcb7653c669e1961355a308bf4f3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f5af0e9b9930d7e5135d5727b32dad7623ce2478ff877f2630f5c84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb191e98938d3e553f102d7a57c89fd43358d4f88382e4fb8c01e963c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h113060bdbf4e9e624f8e1049f8ea2c6d5f6d4e2749629e07d1920daae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148761f6887b7a834387f94e697dadfcf9438332e699b17b13f82d83f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c9bb8f981cf9d46fd916f27c7ae2626789c85c5bf6b5f1f0e5e4219;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e32a010a7f1f5004a9eef8a0978b51a4db9bce36387d71cb75612087;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hba412a57eaf37a3521e866e31e38873195cf877497a4c8b929ac8e16;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2a02d09994450629dd020c2708cb43d1ff336aff9f18d7767a42be6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c6b6c4938b24b142d0806db7ac9fdc2b30b0ca027dad539d3c83947;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9d529e3f8afa840ea23ee2a8341e13e8f0b07d018389abb30313853;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha04a8c303aeb26aae87cd7c04f307a90021d7d30d2a11b2203e6b5c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12763ba327d342136280d18f27add5ae14125b911abb923d3e870a0ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb38eab8ab74b582a83842c5e04a83b4e50ee30edb479557e1bafd63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17615921be0cc302716a62caa2494602edad3d51c48c18123b3c839ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcfb0b5faaa879e02b832489355b3c4422fcc7be4edb0f22affe8090c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba3b19e949ac889576ea7d06b18f3a5ad7fe8a6ae77d293f83346ba1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h124be626362f4cc066a2181747bf7567f8dc38e277f56186d0928ab04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3395c2ac7d53429faf3ce759eb7839bc17bee97e96effe425d30af0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108e56d0158367e7ee49f9509cf78410caa141fcbfdb0717f17d8efd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a770b89bfe13af1e239383a2fb3289368e49fdbc3dad6c944ba61753;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf70e5881368a8c5ba3cc854e5c2ad0e7a4427be8a8b01038a44b2fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac2e3e2b9245920f9094cf2eb94b367ddaf8e0caaf7d234fe15cf1a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b9edf1171d0602d737c56162012244cb877d850f67f07ce8ea4c76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e4092cad4d029efa9934dad593544199521f77c38c4152b2c4b95611;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha48cb414e72415405b843713965276c10cc8b2970d7ca5a67e70abfb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf87d10c13f10ed7d4eafeebd5a667957712077936080f315fb75f6c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d60eb91d66a5adf92e019b6ed229410c2cb41ece0bd89b682f5cc8e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6006e08e94c4a415d8039ec725be2a219f8c30c28fe18235831941b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h201e3faabce3800ebeae0d7634f9ed68c39172a0c96d9f09c634008c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h170ae4a080442a052af9a04c1361b6ae4d4ad3a805a1f74f0837079bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb0b9ca86c7e63d01e98357193d4963cf718056de98d03625217bc23c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12100fb1067412bc6e6c4ae1bb8cbe5d8cd0a46e73367f693b0dbfe7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ecc9b4ef8c398f55c4829f63e74dcd84ffe16a6fac0e855654c51e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19ea4a6d1586c59c8223d3a82baf03f401f4f012a7eed62eeccdb047a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h465bb1ffbeb96eddff5d0a36be093003488a5063a842c9fac638086d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12194e726e208a7480d30ec7131293642eb3adcbc2ecace84bf081b90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h592a442f2896a5f9ff349677e6cb6c96b37fcfb6737f5ca213e25931;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6df7697ac253b79cf63a47a7c32e743c857525554d5f5d615788e86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1e060685b6db88ecac5f215cad9087eee13fc77eecbacd9c4f3bf9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2df61daf2bbfd18500e7afc9807246f976ee418937e97e187ec2a90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49b75d79d08a576971f55c62b7ccdc74759bf3850a55fd506c65ab8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f47b59faa0d570c2ede38e05e9709b7b029aa7858a53240fef97c50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed014934db65efbe1f3600054feeb7c2aa48b796b9b252ba99af1712;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79b8662aa94d13a8b6d5765cc79511311884ce73d58d2f171b473647;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb61fe0d40caf9c7e187f66d97b6797289a399319c94a95780d4ebbc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ef38e42f6c2d09e599e756d2b5e66e3edd125f6b504269658982b4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h124402462cf1a2aef5ef2f125b4c475df0a43f3307937ecc5973c5a6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7ff95648dae5395065741e3146c4e8b8d20d46379ecf8079e49384b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1afa686ed52c934208df3565e83ad39ad7ee92e32e5333dd66412d147;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be714e5379fe58b53ac2862defa03d00d890145312a320efb781ede0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12794db4db2b8326ef667c83e9e92f1a62740c3ad01619f1eb0354ce5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha59e56a73c51863cf934ba9e9c9266d53858efee0a669417d9265560;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea89eb95f362974a9cab360dfc8dda09995f8bf83dcec5d9baa2e89b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f358c464d449cf67a53dbf84fac021458fa58c488e08bbb2821857c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16472c71441465fe81e5d59cb49d49718cdc8fd05ea7b0e71419c715f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb29b9e32ec82d3df5b276c32ae462eb9ea112533b9cd6947fdb157c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca41b3b78f1f5e26ff64c26d04e73329c86fb767eb25dfbe581cc384;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc973981b8dd99638b73b54b664274c59b500eb8b2120e91b3a1982c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fef14e655194f973cf2c295c5a075f27744066d1c46ef0e0227069cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc00e66afd3f796133af756d872d87ca5be07408964b35b49c57b538;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fccc0722a9079a12f2abfaae1e8c4c762043155049cfe128be5fe6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b3542ce6403866db78b42c66c7178d5f4d06d167dc2c1f0cee327d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb28819fc8bf34eda43ea1959f8a78a945ea575ca26ea224c193afe9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e6902381815ef031ec8333a91754c7e2057af8d8f72812aa5a2dbc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13442e9bec70f4ceeabeb8ea7eb80f16cead897168cf260ccfa154b30;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138d485f87958f1cf835c3fe01c90ca03d712fc5cb8545007400e5217;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h156af959f35689b41d7e09c07a40ee4af779ec41c570fb7f220f28bcf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da62a49918e4ca699f1cf88bce1473f9da37ed65e83b1c968e524085;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5bef52442da99e23ec0c18879614b78632bccbcc8456cc7252a23c74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12841b16ccd21e370b313a2d51a29de296d7bf1d85be6828426a058b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8abc8125ac2075e491c2e953356013e26ac21aad3ba2d2abe87e1dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b424802173efec32d062e53a2fa2eee855dcc84a0a12c63b923d216e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c20fe9fcd74e1d8307c0a401afe2ba811df967c7bc1be8421e9b6857;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c024a520f7fa6ee748c710044b6b0165ebc5ea989df5a8907b16b472;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d2cc202e8e26145c419630de0b3ba9bad2a5dfeb4bfa00c852b916c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c3a4e90e079de06717d7b5545da63b2253ba33310a43c03e94883ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12aba95d2478a69bea65c8682f18e2f6f036c5ee54bb969e3b8ff41a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f5a0c71bdbe23524438ad8f4b9863ba766f819e807dd6fa435aaf831;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h121d0fea35cab45b718c580a3df8cdc7a0862cd33a13c06a62155ba06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc5b1778ab2b81ccec3554129cb1cf1da32705cac47750bfbb92491b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc408fa9a4d644407bbc14367b9d0ccffcce8004800cd1bd85910f4f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3263f96641db8e5a97be3c032a5adfb5ae2de66d4cbf9fa69f315fcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha13df8a4532ab8839a16ff7860bf4b21f3d7fc0956969374e1a35f1f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11505a5e309809e923753a5143905a17d61ecd4966b811c1343a58d71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fbdb6ab97a230c656a2e4ecbc4f09592bd461ec1f744dc8e31f7dc47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1937b100d2b51e94cabcdeaf85f8f338857c1d1addb1812b16ef305d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h827f7ce69a5fc81b5ed5f9a6cf1256e6e327fd025c9ce20aff2722f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95b0efa31f0f652e4c3da62e5e084ddef47f65469f3caa98777c3edf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168af1eedb81ab4de4fd4112f52b6715c7fc9c394e2436af758feb5d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef2b86ecac2db49767565098dfb1befa4cafb3bc43d281a138e4315a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb951e349cc1ce8d1da74974e23997edc9f6ac62e15fd9cdfafa3bca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d461a4f03b13eac3bfe2b3f0a0f8c3877bb451045e9e5e04134dd0ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e36861444929ac5017e5cf04557d08388e4936df3b930c2384742c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43460f5e809fea83d03e74147a67a8d22c8075be01cbbba3702d27aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18547eea4339775dc7548c91fc956a7f0bc060c960551f279ecca52c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h60adda90613f4379a15239dddd20e341b6a85a7710b8736aa031b5f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61ce271bb9d47b7120523fef3513fe2197afebe1656c4dd478d6d1f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde1edf0d7fb9258ff7276d4217ebbdc4b7256a1533275a8a8f408839;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a2ff680b16e144d8df2722067a336563ac5e2d18003f4bfc7d05d1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a9559c6a2542631838d5c329701c9ea437f1b7f292372adda8b067c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3963ae5c2b2874bc742ece27a4822a7a70972672dc8f3ba2cd87419;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6686733c22333b73b3e8c43bf55525e3fb3116f24f48f71274f2d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7fdb6134c065bd2c146346a13ba832ab6e1ad1c1b84e6b336ede4832;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152e93a980ef30a07a0e82eaa5965e9cfc60e4e6acc439661e411d8b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a4f3e168947354918c2edc70592148468db080a656f7a5e3cb56f993;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8db1ad26c02a09f308960332fcf4cb7f15aa67826d99f4aa67f9937;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152d660698e596e100b2dd95032790d7bdcb85bcd04813f75c3fed7e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12df207027de66739195d22acac8aa5b97ca1360ae5a7cd7f7a4289cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7d836f26cb666fa6be260271a4aacd9880883ed882305c7fb934dc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfae51617f224cede553753f7e0eb1214ffaee1577d210b2e72c2b9b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6be9815d09ca528124dd7ec9fdaed82c18112b21d2791a2c2892d55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b8cdec432b031a6765c2479f8e0305af022c62e0f4dc5bc91da4d6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98ea3eb698ca4aecb1a71cca5def98d9553116570dffea7f48f75f22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1399df34127646addb9aa55ee980b4b6527903bd11a4b8221ca517afb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3668e580096f499edbb32fc6873002b75729324310c8761f4b8821d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19aa140c3228ea2ff09a05e4458d5a9fe88b62322420a5ea18ab2a0f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a345de7bf29869ed74fd4e6a8983df687f8d2fedd61f3d1b0343541;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2fb2b71c5bb157365391dcc6a01144188f4f51c8e858bf4c0b9d284;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1759c0faa6605acf005691323063b860be0c72f806a89a8ce44b666a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h682f11d94163a846c38e69f5f1973a57fa1e54179d7d30b3d5460a04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4225e40a8613a3bc120605b26fc06ef42facf995fbc613f5b5f0b05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6cd712169ce4fceee09dda35ecd23f5e6fc4d855315d04e12d4c2c7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h768c654e370bc68ad424a2f8d5b6fd9a22e8c73247aa63d0ba16bead;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5c4d753dd5d58ca8fd81e7484215c9615d3dfccec71b1d9c5203143;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a8ee28338497b23bacf154f5e1e5437bc703ed0f1bb945448b355b68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55a3b439a13467a6d46df7c21cd0b5ed749f87a7b740633b3cb278;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c77f6651af6a5df3eb94be4489d3ebfbfc4979c570ed09b18d7e3aa8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83ee271f21cf98aa70a03276a7c908aee7a3d77e05b8b6b33d66ee43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16662bd9d9b47f4b6f200cc0f9a8adfa2c00ea7f8a94280e8e510e693;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haca18ee41f67d067d4db81a03176546fb39c6ec49f53fd58bd3021fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he42aa707565e7c42b4ef3c445dd79fdf534e88f7382fc1e9c984a40d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9fe723d644b7df84d89139ba1cc90e95444a86e961c12f8ef12ba35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168dca3f3ef08fa53a4b453926edd9beda2d196562e2d1b2fea6e08b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49b1e7e20b8c421cf70fa161879d823440109d7b6c67b80301e3cd95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1498d8e832a159ffeaf8c2978a00e4a06d275f9d665ae878a66758d23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a25943203d87bca2ab5ad31829a973a5fed92623e4505cb4fa26403;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha354f51e5b1b4f9d42969086dc36df7e9c6e79c9f831d34fa8b5fe5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63b432b5a7e78ebc957691bbcded0af0ba90224a15ce0873922bb4f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28bf67521a6c56a16e9756797e8102209943d819aa81c3b4e62dd98f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h124da2ec8f8c65bac3df1a97068da5c824baef9b54dc14ca9eaea1272;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a12e5b3d2b9199a3679f30f3a7338c8450caa5af0244cce2748db468;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0ffdb1e294afee0da48ed381eb7fb8236701369d0b653a0e0a9895f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114313fd35056fa8ae9cee98e0d59bdd381e471c66079d9eeb181c44d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf71b649d3e189523ae6ae260c7e00afe204eac7ef2fa2f4dd8b51094;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1682ebb7d751e933a10bf2b9abc43879e0bb927cbfe878408237d0aa4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fad83544e6bcad919c15c511ec6d6f307ca0a129a942eb71a898ea0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19eaeea04689207dd3601dbfc2a6d0a2b4a0a34d80447f03e9c4f4f74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha2f7fb083c32a8e61cc10d47ae5591948e262429ffbc7bd1a32cecc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4c676d1a8474922da91438a7cc664c5ee7755ae6533e60343c287948;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c02280320efa24fe72ab04c5db477b36dccdcf776eb7706aae14836;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee54d6f6b57f37f7402a34db630a733c1521aa4c570e76e04c991dd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d099043a64b7b4806315770f6358e7b6b9a06e9645da92c805c1b45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf529a460623753bf55a1bc378536a82a1cd3290c09a58ea6f149658;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf82df12771a63592fdafc647bc1edffab340ed0546bcb369da1aa2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8fa7a841e20535ddd8b75314a41ab392c9828cefe464deeff08ebd72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a878ed83058ac65ee36cb34c6f5ea23f851c17e12df4055f79e10fb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e0e56d26fbce9d10e426afb03a4fcfec74a308e3d0e99c65d3bed1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e520cc3c598c187f1a84f939ab755913a40a8f8578ba0331778dec2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11695fc5fbaf56c0198e7eaa22b1eb76b85e0bb2b73bfe0d6e25f839f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8643fc0dee9efdd3084a7d80148fc5a1e6d2a5ec25baef78d8ba00bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd993a981f0ddb8761ffadbf980a31c1d766acb9c6e6163196287658d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d2904077789ae5d770a2d27c5b78328bb5d538f2c66f398b1d76c27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17131d04458c9a57ab73d5c5f27670b2da7085f4cc8e75b953f15cd56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6589014d48c86bc2cb9e2bc85137be703b824796e2a88f8b8e4d5820;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ccb70add7873f11d00a53304e34ffe6e3b9c77e17f1ffed463583ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3375bcb08421399552bbe38eac2db7141ccb0b44bc43d257cf197bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e161728059a7a7bb997292f6780dadeebad02f952e49c814e120d15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dffee9bec8d9839afbfc5b8ec67eed3749eac5d1e6ffeeeb6b72c0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a900937da373c5ba1c036eb4a9d3ad6478e190dc9bf5dad695f0cd22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189f26d8fd1122941a24ece94f09b44ede02ca03fffb182ac666d11ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb37ea67eb795786504f26991cb2ae8d83726726f3cee4fd726d7bc56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e9780ce01a8f149a2aedec3c82ddfe3c198330c359918763f8bfd43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h165b969c6b3e3825e8bbaf0dfb20ae03958705bca7fd47467c4456d5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12fa6561396ed1130202606be76560d9530dffc2c2caa10683aa32a6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2b9eb177767cd58b739771f7c17ce785fa5b5c063f3b28255a40a99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0479e542534150cf65c56420445362d586552a25a8da8dc32902095;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f9bbd3e6283135751186a985167abc02eb367cb131598a178e7484f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c9a07db8d53246fc469ef8365876e805e818f38cb24185eb2702177;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18417e26df345a1d981505e4e003fd36fc83a6d09d2eac6071733441b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffb082971ebf14b0187d45d05db24fe54efeb85c9c1b95b12b5dc8d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1113f229374936987be1582ceee45c28f109b1bcd0f2539d8f417315a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1335d116d3107b852263756c76929f14a4bf1920151f5d2ec122a63c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f3c2e3a7ca06a1ceec63bf43045c7fd749d92be2a474e21d63c8c6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1850f565aa7eec58c30ae26f185785c3caa89d19177f1770882b9a711;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f39964a0c4afce7438e3077fe472b18547f31b1861f14789bb6fe552;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h901a94c0193b93f5894cd89a132195b36be1e1518e01db9daaa65bfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0d203e22325f5e99992475832c427a1849287df76e3438b4bb5fc96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49bfacdbef707d473518977a5fa31951d1dd355fbf66da9aa776c896;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f6429ed6a65558f2f1249f02011aa281190e4d0b5d005fcc7ffab394;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa920fee7a9ced50ab0d794201b7df54eee05693de95c2805f2646d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf181b2c924c211d567c0d5f4b22de3b8d465421ef72a55524386235a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e7ad66123c5d1a85573db9fe12a2aaa4540756af836ced7b64383888;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e6225b5caa74d99294321f8b97754149ff46383dfa41e782e288c5f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h101d02503e1294891ff81fd4a1fecc3dcf8fb7a095d3397ef5b9d07f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h147937449f88c8097d810460c1ebda3a4bed4f9ce0bb3b181527d655a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8484f9664c4e032be8b5397868b929c493144eb38304f444e082ede;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee63e095c1d06eeebc7dedb6e1a7fd5ab7da76581dc4a8991c45de22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1079decff621b4ffa857bee549fff5494a96f6f357354e8ae46dc36d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h813e871a0f337bc9bad33ad531dfa99cc4a55a612dc57a4b0e374d89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91813fae1e7fcf6331486cc6993212067d9b509aaccb240603a69717;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc481b38a9ddd534fafbf9bc1530b6ba8cff91953c41d661fffa661a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b97cf0d79c8606867cb30ae42f0372972cedaeeda52825968f71db11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1caea3ab512526c853e5f7c71c9e90b3c0dc747c2d59e57ee34808763;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9e62b51cec00ef6882947cd3dc7620b2aa9bddf73852df3ad1ed22c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f117894bad4253ff26aaa75033e6af4c90ca03f486fe48989676dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc5daf40b01032880711146a58a5c5d24a5fb99b388168c9bb738960;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b47a7ed1396b0ca5bcec12b4574b2bcab6cf7594cc243d451f2e748c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43f561ce75491135edd49ac763155e9c0d5e5e73ca9e90d995d92229;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c1140b7091e3dbd7c7d527d011314841f1cea6e43a3eafbe0d6d288;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32434813d427104069fcc5599fa7745bab3290f8b1cc14c29c0c1088;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd8bbe6ee5fe1065b8e22d99b35037c4b86b87a95071131a470e2371;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1877102cf0fef0a28e445d93526260f6847f8a7efab2fec515e5e4f5b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha587310bcdbac89b361a3050d3caaf3a0da6189833c81ed0fbd299ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1603fb7e082fe9b34d893613cbf71cc88e5d939d34ea0c39650ef25de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f4e05e59cfafb0fbea062f6b347e756ab3f62c5cbc34587dd0b5163;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93666c25d391e270b6781cc8dbb49fb09ffbc7aba9123f41ba81c63a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbcd6156c349ce05787357012f2f72847268e88006adfe9359b1d2bf9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf7e060629bae8da9d39a04f54ad2a9192c2685166c59212371ac4262;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae5e11ad945e3975afa8a9b24787d2a1e28e0d244996700ce3a266fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2d217b886c0e95fb8531b5e968099c1573b445102d20ac7d9d6e72c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he3688d18d63768fe3a5b218d3acba76f6ea558b143ca3e39deb86cb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc30f2e1ec12cbcb33c84a7a43ecd8f2aff4f752ca0c982ae17a0b24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1701f6e404e9f31a5116bba7c48f4fc6240523f13a59f82b001b23bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8549eeacead0ca9bfb9cfa5a664e651b8392f57f8f9b7f23a57eb94d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f99b833dd8018bf1ef67ccd7b560b3d79842981cb2babda9ab80576;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11751c5b03f51a70df679e8bff29048e888fcb10efe1ca706b87a8c9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df8c8d339a62769da699cdee4c886df0b4b7d064ae682da3e3bd719b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185da9d59d86eec45bc11f1bd1bd6f83fb9ca75a6cd928d45ca9c23d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f71bd806fd5d566c247335abfea4be2135aae3fceaa28c0f972d0dff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45bf9128c8599afc950bf13e5004b050da6b8fa20ea324efbbb71804;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c5e79eae9addecf72cd669d0cc794ef8f0886a1e2fa1fd203f003b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h552106966dc52e8c89215d5ccc59dab6a1ebb6a610eeb1da680fcef0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd284fedfcdf4c401c4fb4183e3df0282f5ce123a446b1077b34c914;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e17658066dda13923935475a9a84978e5ea6dfee7d455049c3f9a5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb273a7b59a6999046191c7b68d7f43de25c10478dfab5ba420aff6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80b70e0740f033e828466d9a22682f6fb8220b45354b91c4d5bc367d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1681a2aa0269e9a02e81376df047b2df04189565f013b77d2d96161b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb61e497513f03413bd1978f88ed58dad35491c126d654c653fb316;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h44b6fbbf12816acfc53276d82a091507f2ffaa53d2d86a56f9b734ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c9e3a279f068d2d9177ade75eb200329dd5795b2b4dc8897feb1643;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb6195d3b66b1e3ce73834960665bb83de5ed06ef85f945d206b1c77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111b644f9cbdbe5c186af287f428fb1e28889e2e2ab7c32deca5b76c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ed0fd7a2dfe2b9c701739c0e2e0747b1bb52af2c1bc3c5333cfc40c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1462b6cfc46fcd102ea1c55f5dc5b7ac10b2a2ec4ff49e8a5b383d66d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h444ed533dcd032b51e96a520a5fb201ca9094760d1c0fc3bc8ce7732;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17b690f0a861beaaeece7ee66f09b3a7d52f672283e94b3836b3aebf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f7c5319db13de6b0261648670500606b457eee65df4fb565c91ff9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd68faa98329cfdb3a823dc248a021dcbc06e2d981f1374e4be0cecc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41f93f3a6bfda1db704a08f34b0dbb19f11ec9d758bcd3d838cff42e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd1e653ceea972d95f002c19216d6de937987a148e97b8b6face0f2c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h175813d9d6aca794a738ad0d8714048fc43ef96cada12321b96c04e9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d7a26cead7c4056fd95c078d61792ede12ab7973a6e77720b7b55139;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a33f465b4f137061fdc9b1bbfe331945a1fca2e2707e7e735adfe943;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he028df74f28fad92db9587ee61d245bcba0d6882065c6ff463b2a25b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c435adb0881c8c2059186fcfeeaecf3448cb2d65aedf9b90f0f0a01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176be1eda655dedada8bbe0690a7047e2cefd5c227f157de920e2078;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c990271eb277385b37d628fcb0ed3652b2be3103a733da9cc64e67aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4398d197d7b4ec68c63f94ec3231e8138188c6c68147a2b305bebe32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c0b4e2e7e40cfbbadae03ed9c6420bb58a013af39bded654eab8bc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5393007e4fff871df910adaa84c9de80907cb57493cf3b4a5750b07a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8035159838707eb80552d3570459ec4d9a64378e3063f5fd2323ae68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15eeeac7e153c5f84222f7ba6d3c24cd784e00e3e52bd61cb4c584f4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h938808ab54dd5e481409c3206c847bc05882a1ab795da6fff8bdd650;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc0b668df184d4c095b801c59b8449b21c77ac77a99056494d60c4e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf975b5cba7e2f4512e09b37a92981e5403b17dcd52d4b27fa7479dff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c68f7853899eee4ee3756aab8f2585c460cab584bf6dff7d2dec4639;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a22ea76fd9984338b4a5d3cc47582277976bc4062df73fb99f4e5b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he323bcb38b68258d4100a8500eb549ea8e557728f9636cf2082d7692;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h296797b7ce6e539c461b2dca5129969d7be0acb8d082a79afe2cb49d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb8d4fa272be04d274989b1a41b68213ab6d069d5421ad93bb3f2248;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16fb07f2707c5b4304926344c8468738a5269c78dd998cbd6a357cfd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91d90f0cea69d8faf323cb3651160672eca7f7d18ef8c81cb59c267a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ebaf3d085add7f56074435437b12800bae8467dde0c82280ed109c19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157793a05d72d71b2c4ee5c131cb95ba8000e29bed753e280c58e5dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125989c76883b5ad33756756d3f182062cd29d384ef6b4a0370c83357;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h318be01035e668a3d0f825b09e14dd94ce6aadc678ca8c8a388e8761;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76246f4a2b3ff5292f2f80afa9ec3cd85bcf832c93b0c43e04935068;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1190d12312f6636ba034d79f8226cd6e4a04152ce584e3c420556a768;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12518785cd8bc3c0166ce77a547c0224323c95c85070a186c7758c515;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc40a931db24cd4d1a2899336f76b4d44c34319da8c0ffc2e78a14dae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2aa55b0294e79029d0ea384e8b401eb997b6bad5bb43b692df9666c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c11788238255add6206115da7e290acec416215befb34241082c271d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h175b8fe18ec1bbe9c3cf497052e1b8a7753d573b105c5d84fecc6123;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3102b6dbe73172dbbe6092234b7924b8255f78dcf593fa4993c8f0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d6eb1c0912b59fffe656964d60c892b73985f968e58955f9f40dec2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6b6b2e5323beadd7ca453ae0494aad54ee97ed9770f5f5562c11abc1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90cf1defe841b1b7b8d637c1c6d4f2fa8e515a648adcb68f815c7413;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16cda3a24b9933385bb70b822a732b549731cff8afd94c4b858dff48d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a6ac6d53b273ed907d0928b6b0a8eb08abea280e3e1bf706e7b2c85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a042d98f2358b6d8ad7605ce4391a4061330189f5703290d8e099a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64a2a17b9929f9e978b38fe64b94514bf0599efdd7fc194f64ded27e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8235cd3dfefc52f6a664ae003a4dadc1452c24d47829d420502f4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d3fd512d44d32c351ab9a99cb126571df606d8ca254dd242bf22a685;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d748f574083851739c6d535bc889a4179da8d2569c1f00f432e55658;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha011087cd4f16dfb8163f17d96f303d62b7947959580786a8e442faa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62aa40de5f5028e6e0b99c724767464ae512f604195d06e011c6e515;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dcd33766083ce2f9be9191b11a0cec0e1dd880fc3b67e13bb75293c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8b34622306599b6e11febb3061ab2446b6c5436136cd5953e7d55ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129e8f7c209d983539d9390f57e47c415ff06995279b7f38cade41e88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b2350c652e79e7839064043a338aee4d22f0b10054289e27508dc02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17236fb6dc976af6ceb185f11ccac8650083ff9084a09b902c1ce91f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141bc094a2ee53418cac6304b069445a9138acdad3de3d832f20c2d8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41331f2f5ea7acbc0dde21f52ef5086b3e21a7bad3d58ed9fefe9f09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h121d160ba6a68927c7357eeba42297f86d74cea3a78805b45da77ff2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4bdce91d7068786fad37d65a8628d8e605efc8e9f35fd9b436c9ef6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9b8a1d9b702fea65070d27bcf988535de081559ef922d92610a28da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36dd54ab3bc277284a67deaa7870b522c45c82589c3a4d6a39df2e8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1872968464e08a752ccb5131962356c2507d01414f8fff5a56f3f5cc7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdd8cc12eba01150965f6a33f8fcf60fb833439840df6e484d2844e32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee6b3891412fc6108e9f5a03b3a4e5e6c1291333fad54aa9dac832e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19b6a5fd4ecb3be8687d98a47e556949b8c0121a01729cd83bb99ea83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f12917168745a359869185b322b72dc9e590eb0244e07a5fab25a11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha41e2c32041e6bb9f0f1209a1d98b884b8964d6e80230e75f2c9ba43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h715b695ca436f49f7638ffe2d115db9c802e9a07011f6c4bb00ad0a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd5ffb7efe51a394aae4314030920be2248c41ef814b846bf25087efb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1424279b9f846f41221d611da6604d5246308b958733ab0f1c25fa21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha472693aa99c77753d7f52086e321abe99d5b387c766c3633345764;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb9fa92b3b40364391604979984e1ecd0cbc9df53d395bd73b666ef9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a90311bbbcb6a254529b3dbb1f20f0d35d693c7921b0985ecbb9598;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f70e83bc21152037d93ed0f03622b6811108f95d2cc33f5f019a11b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc67e9b51bd89d7b1243c5ba891c3ba38d8704ab93dc07888d85c580;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h25c1dc384657ad73c2f587686c15b8fe05a134a3ca121dbd82e34bee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ee0daf249fdb8327039c5907b005205124b437d3d1967c728799237;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1980a51d9c57ced33d5f05d3d642b6008cfc445b276e4f1d22bf1708;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfcb2c92059d35f54f80503a37079a16f22ac1866fc538635ca28f854;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe1e7c0d8a836f4da85afcc3bc3a865ac2a84ddb4adcf625e4a0b64f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a884ed780f74bb09979d4005d897f209ce248043240d4d716981e457;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha23f8429ea6792ffbbb223a3685f085568c0ea46aca10e7e2a698d86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16dee30da1ac504e646f0eff5b191a0d5fcad616fd69aa6aa3da315e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ca92de5c63dd5d4f52c42513bf7df7ebaeb2e67b2ed87d7d9513a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f6037cd173e2197e5c5dffa75ee09a1e282cca24a08c948a9a4637b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f164d02942f2b0a2323c3612798e94b082eb7cf02bb5f04b529b477;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1edc958f9b9cae87a55696840903f2d401c2f6ae25b4ba4b438ab85d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8fa6263f5e317cf2e409b7d26d81683c01ec99f53926d644d74909d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h548db7c17a6740574fc538b99896ac803d0ae78c6183798d11116c5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd4e1288c180cbc87e87da08440a7a1c86ba9b2bc1749ec2481cb73f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aadfcf935e524390b22ddad43f431bf98126c60ccb1b18e702dafe79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef950cf93a1d8bfcc912c9bc70a135c19a8115896a28abac827e56db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h203ea129277debf49132a8020963082a9181a9642244f64560432845;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90fdfff891fc517d3dd4f9e5af0e6ef02e183801515f9d152fbe4ead;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19320b94341987cfa7187ccce64a38ebb527b50ce8f27d9dad54d0f3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdcae501b7a4e13bfbbcbd916fe24a72fa14a617f6027fa1d9a980ec2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1e3e2bfdcbf86f0a1c347e9d778f61086d75cc837bfab7fad5a0f89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbff8e22dae7aea0029c907f0f5534827ba387695894940f2713eeb35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed0dee436fadfb3ca94a82ea49c864cde7a0fceea97dad3e1346e568;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f0c616cf52e97cb7aaf1a4c35831071dc73d07193f400227fbfaa2e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11cf32d74b476efc0d73aca57be495dca4fd4adec1fd3b8f4e837d00f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3c79dd78acff7e2ac5fbdfd6d29d159bf98a8869dc4cace7aab571f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ae170ce468ea79ba9da850c3ed81953c48464fcdebb199664011df7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184ad6a12316b103f58f5ad52ac5b356494666991a8db2a4b0fb54725;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h287ab11a4ebe5f910ca3c17ae4b0fbd06893c3d5c310f0aec3b1d22f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac5490c5eb7eadb1e2c941a0c31f30ce8aa042041184ddb41fb6b8d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha2060abf81d183ba82e27e13e23617186ec5c47dfde6a6d22294db04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcaae97489fe0b2bf8fd9523e8d2771327de3757b91c46e5d0ed8ccd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9416e1522df81fa7594dbf5188b33214b421c3e00faad61555188c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfccca6bfa1cd674286b679cef969ed708feaed8e469abc961a3a19be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a1d7880def716ddce54245561b206d5564911c6564c3e74404e1b3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f73163f8724917dac9e920f9c2c330193185401bc91be4da69ca781b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9820a71603036eb4f3b63aaa97594dd0e529bff65ad74af346cf9065;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f09a17f84727827a22f17c6c51af6b8b73d0bc33adedde351c89d68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h334c00e70d43502516818b8f326c6fd62122f2e17a851b21bdc02634;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e17a42d7c2b6320066e96f7db5f7efa5b7a7b271cceba58fe50f7a40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee3127f258e8055608a1c5684e8cf1755470adf542e5ba532c35529b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ebc961d63e362cfe6b5f48a8634d958a01a59bb9666bc31e72936db7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a621c1df4871ba07eddc00651ab97f0f9886b1955b67fca3a76f2f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a62c8bd35b93ac5d4669d74300f59347e044df8a2a0eb0968a2ded0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff55f360eefbde6dcc89ebdc381c53c3b930ec4b9e1ef9c5ce73e430;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e662aadac3491698c97e1fa07d160c61d9b9b2c8200ee198874300a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15535eb5c25b1dfb170f5836af3086f44b3df15aec21c3f4f3b9d2b01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb6466532ade3af487f1800dcc5d27f062687f8c5bf6a277c574d07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191c9ebeedf5285687455eecbd9fbaa403ba3de8117591cd2e531849b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ef42e36416d9362e91d22da6821c1da4c9f7a311865a202682d7245;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0284de1c71ab70fae9635e8ce1507dfeec2d938b816dd035dddd0f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eaf696c636f527c806c942cc1e9003eb8d0aa17e325b3b76898feab5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he65abc895bf1a777b28631c621fa9f70a6a9c876b78d3bd62b14d9e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153d4418878a2c6ba0662d8f51c0ccfe3cac6232fc2c0273eb7c2c28a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h267f45c128604b0e450eecc223004a3f6aaf9535a739ca4f3e68eabd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30e88f05180a7a39f1f0061739f57fb5ebe259008dde119f7bbfea02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61335e881faacf6c4366ccfa7e57962528627e37f9b79c129e1bd9f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc875745c6c0822e809c727d8e1033ee04c7b3920cc7b529ce68ce181;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1058d5cc4165bf9686fe662e4514e73d72ebbe28bf777d3cbbcfb85f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117f42e46383d5714e6e88c3281f932d9803c9216c0d0f04d4eed03;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5d6aea0c015b0b8b40580ef8810e3003ccdbf43bd54df76983cd98c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ea0c50ca61c6f46cab872f050f1b328a798bcc647fe77722481c7a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c978589c7044113dd25e12e1200a51e6187d810cf46db771965f285;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heebb5c9c5feac27991d1588a096c93218a67df66e035dbc3314de596;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb58175ab6b745de4e1f8039b1564974f159557575fc901be756f0544;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7312ee9004bcc2ba7ffec1d6ac96c8ba306b2bcea5434dc75ddc085;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e62b6191c51d653b5d3d402bed95e4bc7998b37485b574f275781421;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e3283711241c0cb389cff2f57b42dec9b38adb5a0abb0c469cf48ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc85cf6617b75124d7d6e1cbacc28fbfe591d662265a2ce1fb54e8e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34f9de2bdcc22efbeb60d34e0febc2584976164aec2dc1ba44b5eef3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2e096e7ed36ca85161b0572e7dc732d67b85f4591a0fd94a80193bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha53bfac8c66626bc9e43f1d79715df2a2b706e7e2d84e906b955226;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f562f080fa9cb859d9677f4c6074350ae167d77d45be5772354e7317;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78bd279afb879defe734b774fba206233010f94bf6a0bc2b1cc4247e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1903711785e02e05183299a16442c7d6b4304220d084d71e39d5745ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6d3098a2aa021459c4fad3427276ccac5d5eff649559c043044ef19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41eb977040b4868d61874e6c138e376e19b29d6a369c6f8c0775101f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30d88e7604436d3154d7a8b2368e9e1baf5adfc0e740555847eead25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h406290bc9357a92e6d2aee1551779b6181cabb9673168402ed5931a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70b4f2e76813e2e0983a9ecfd7884dbfa61beac6219f51a4b4f96d84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ffdb61d9c77adb123133eaeef468edc7d8fd63230957ff90496f862;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18372710ae9bd415555d0a95634bde84e1ff8a41d35ad514e78527434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1729f6daf9c1ab22cf434a65045512240089c695b2416c3c86339b614;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c44a3395941488588068084bf776a3906f2a5799cc0507dd223bf0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haf52996818481403a6a491ed0a96c5ffa6032232f1709b59787008d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdac78b207b02504b739d71110915efb6dfa3cd19483578f0c0e330f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2915337147225161f24b766ee37922f9e224d0fbc025d6489afaaf1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78a6be26752fdbc8f0009196c9fb45981918d5e54bdc1a1d6a871c3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc038929b2bb50fd038a2f290effc8bc66fe69b7551ca697f7f2e7729;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b8356127831d25bd30130cec4b7a35a4b97e7d9b3910a4eb16ef57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111ff6ff861b7f1292877cfef595c44b28f837ade6184e81ca4a8d830;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7330e333c6dbb45def52d99cd3b3622547f9f74c25fed74ca74c9eaf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38635ea185704417e8793db01730eb5aa098a3fc865b1d1e85204fc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9458758e837f3341a6ee363a5093b784fde7e6e56d415c9f8e6e319;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c122b2fc9496221118d596572c701c8b4382a56f5b53629633e15d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde8b9a588dab94c1c9153e9ed32b3a9c6b72ae24cdca59ef3a3149ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc293d9b58a8cfe5905a4ac9b5b2db8a0987a7f6681195d640e9619e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h449dd822627d4ce3f6a3b806735410a648f0e2964fbc129e89f92a57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2dc309727571c08f31968894e6f9f1419163ea1913381f20f527e11e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b882e9a7ccb007206c32e0bda3ab13e50610cdb4b70931851a03f9ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e0e9989ba1a3fb651ee8afaba60ffce42d163866737e497f1f97740;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2688978da3d8936009443b029f8a6983a10715778c41056e4cdd666;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e912dfab155287731f9602ec131cdbd4fb31a13d8818ebdb4654a8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf47d02ecf3683cd3a2249b3f325ab68eea9875d2c0c3b6cd66069105;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f58cdb78990c9b99c02b1f349b25b591b550b05336aaacc1daf11d1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123e657b97c39a36963e4af30688f6588d2dd85654989c4387aa3b52d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190bfc142b5c49fa7b0bf47941bcde296dda8e3f99658184b046b3512;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aee8c68eb5d0301879badd33dca9f39f63852c0dbd37313a6ee7e85b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha364f5484bb4c3403d8f08f06a28aa4cd4532764060763376240794e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a6ed2429a4e7e14bae3f31017a6d5808cb4741039b0e9dbbd1acf2f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a658e23112e36884da107398d01b427a530051aedfe013b58790d00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2ca4f5c01a69a1dbc0a76610a9ebab413980a8ae1f01a17b68fa4a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6003d6818253ae0f447ad61899178ed4a4626e813bb85e0e1ed87a76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h160971e396d3259c7d3b37327454f09062e537723b3f3c232a6e25995;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17002a3fd979b73650ba867d8a1d98eca1a3d4ac5989c0020b7d26b44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa9c6bf6f549f3c64db3339b9ad605b80f3ef25cca26de9b2a672f6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d02d469580304fd406706913864637d0211cdfdd45990457fc4f4659;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1702ad87db434b66ec9f92393aa9c1282d751423c6866c1179f977f86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190a543601da7e1ed80abc5eaa79d4afcedfa2962aeb5b229bee2a045;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1367e7997b7cfee83dac421ad70e9fb504660ae51524cfce74f4fbded;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1514cf5179c68a6e977c3abee533466fcc7fd8a832b407402552383ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a25d6d6f6c7d6d68540568ed8a009d8622cfd379f873e32847dbb9e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3083000f2f3479ea662d11359afad93eddcbb753f09034dec07ae87;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb4074f5790097eaf9b8f4f73bfdbd2f4fde8a3d0c0f633298b6670d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ca8a1695f7af3588cedb34e254ca54998edd62bff3ff45c4d05e755;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a42fe64ce4e7edeb801b1857cf5c1027d6944a59e0bdbf90ed27b383;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b749f3f6673570a9cbe9f4490cfa054a092a6e30471d55fdaa2d15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha39cd37f17573a3aa24673267e637e2158f010b582224de1137b61ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc18ee816ce3110c0199984944983e8a1b53b4fc2cdb49ee4ca7b5e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c16e5d0ae94176293c41d132af5790e82305d7ff91760ba08f043b49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3952f5c62ccab13e4d18363fcac15f317ce44aedbed5fb3d02b4e87;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc5d88b7d189eb036f1ababe40d528fd51d6c71a5bd8baea269949b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa08919123e670db19fb8a19c3a4750ccffffca95a7d9fe00dfc3e62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc16f527b1f0efd1bf5f0f8b7baecdb7ecf62cdb1e314121fdcde947e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h69144bae7447376e06149e1fe974e83f243ae1016540c270a104a8ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d03612b6087b3fc884ff4493c511894d3295e13ba81c33f0d3cbd724;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4f8aa35820a405ab73fb4a1bb89f08f1e2e6e2e5fe33d613841a4e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ae93d6bce4ece7fca885fb75c6bebadbb8dedad5190eef26927577e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b667591dc101d993fc58b7e979e1b4097e0c7a30abce6f875b32d4de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf121e528e425602295d848185b0cd13fd9f6f16ccf6a137025fc4051;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h748722a38b471c448d4e317ad11e3c8774e0998a637dd479f49c37ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e63a4b8bfe8ecca1cf7cee783fb1d463e43d9fe7468e997b46fb5d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9d0803c11d5ad9563ee196cbccb8e0daa38634a095d5185f814b9ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1272d08bab07fa7903aea52cf890fd5f6c883fb0ca9cb7d4ba40b6686;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be68906d83a306e38b3704d5cfea141d5164baa2de0a2cec7d05e1c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h725b04a0b9dcd617bfc9c21bc12ad89aa02d16aa3d5d9f7912498929;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c2f2e51eb487f703f2118a770fd075b6ed4aed53757e94132b547c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120c1b208a9b8026d41ac99ae4d948d39b2754f89745511c16733cfa6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169cac4f71391cd197e633ce38885ea4903071fd3a6613ac92948c6a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f52c5c995653419177d4cf4f080836fa258ff4da496f573495dd36a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9cc64b78bc1982ef58ff8abb3604ba268a29e84439f8795e4869e3a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f578dfe95227ea4d804df1542124d3c1cb2f4174f2487b76118e0a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e48d477dc8faa83e14a462a10392c0a297227299f7ad27eb061eda81;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a707f0406cd1ff263af25ccb290645e84c4ea3a5b89de3fbf7b2d2cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a363795cad0f12757eaed463bd6da39c280376d842358d5d97390e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10881bd700c1a0b248684ec1ee01b0dd678f7eef296742d9162b39ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133ad8dbeb3f4a9b74c3fcc6a55ad7b798c4b42fbf77d3febb0c669c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f8603777e3a85eab6e0745cad9344889693e7417b1d60191ea78130;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d22cb29c72e43ca09f7c9b604f1baa04a648b27f18d25a69a078a2c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h145f7268e49a5acb4a339f8a5f42c7e2fad634177bc260c5a2d635527;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h543fe9e53b28dbd59ceb859a3fa501338011733a21792261b4db59f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14540d46c3a82a61aa12c514022f585245d6f99f89c8ed0ccc6931560;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1285945c114d1b37919a740759176c0aecad9314282f1d1a69ec096c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2bf7bc69fbec51f7b52e09d7ad83732b9067aa69fe17e4d1ff6acbc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82e98d5d98ecdf3b0019df6bbd0d4389ffef4cddc352376ae5708880;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b36db0142be46c2a31e1086255423945f497b5501044dbf1a1da3292;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1608c7a9ccedff360f67ce9c46d8601661d6bd130e0d214f58d330d7c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190c4c483fd7443a9b73ba7bf117d231adbe8bec217c487ff5e3c2d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d1a250c6d680f5edfb4500c6e32f6c376a3211928a2649dfb340d19b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1acb03701d7c17fa4ec768b173a5b45ff7e9c2bbbde61e46cf36937c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he555f6293130c12feb785a5a0504e9bdc9e74824d626a3e9c72742de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had85e6bcb9197720a10f3f8146f2657904ea46a99fcd143080823400;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h132df2ca49c40c25cc7113b8cf41dcbeff196eace15e0396b63a5d313;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d56494ef7cfe694344211b79b5819904bfaa17e07562fa54718e3b22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb5bd18941f1378970f2afce6a720208bdb4b2f80c4005a35e63205f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155db7232d40cce47cca5463c696292462699237f8d41d95af138a347;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdaef26493c8284e5814d1a5eb27229624bff57ac60e19fb3d06580e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a728b66bc97037c89f29407961667c0a759877d9293f75a180155f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b5a7705f170417d5d09d5f5884230ce44394a2f69918684cda80c41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1608c82ed5aa2fb42b3f8ce8da51a8a0a713d0c968cb4733249299676;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h890406ca5f10ecec0179a9597b65a75e77558f1c26b707f0ab3b5e2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd42c3b8a17af67fad2089caa8fea1343db595ac9d67d6d503e37e25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ad48c182d3c4e88c979a1d9b86a96750b652c06f14351a5a26dcd1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h165b2c569f868f872246f70383e98405c174deb8dcaf87cc318ebde93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142b7122584e7171ea8ff9f477c7e830a06bb37a945eb6f6c0549590a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbbd7e07e40ab363d1710c7098284d3c48125b22672f79ab44ccfd6c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49fb3570ca483108e398f77ff197e5ac263ee0ea7c97cc6fb2d0afb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c3d827e64ccf3a818441680a2509b5a287cf927cb496dfe99c3f6a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8343823c98be4dc230cdfd4ce80c23dab84ed7d48ffff3889cfc14e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181ea3397fdeea94cd536b36d060202c1a4a9cf8f55487f86a65e25b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h593e1bab90f9fde15758a62c5d2cd4c979e12608333c4f9517d94e20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d93cc586632fbfff99f75d4428ea1e9e84aa47698e60d2e3db52158;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3f172e6cd7cc57d010c43acbbd75e7f2d23c8db51d486e09cb1a59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b056e0c92ac095cb58efa725c2e4cc3e3dcfaf912eb931f41e185c9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h982d65a207aeb2fe3b5c3b3740693388717a7ed8c609aa8702e09ef8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129d1dba4a238c838df3840ee9e6de937db759a9396401c116aaf636a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef88ae63ebc6c4fe307a9ec2c92fcf1fd65e2845a468e151f9848d54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a3f7deb03c4d6acbb62c2567aa97b9106237af4d0b13c42d97b0a45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h403542bf66faee1a4cf3163c6fb355572b10830653fb96e557459e31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h980d7604741a355bc62688dafc8ced0d2a29553be5276ce832c32fdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14df17adb99da632ba86131057bab1f3f31380346b5eacbedb4937695;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h499c35b78efe394bc8c70ade24f94edcb87d6980ecb051fa0c9f548e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb9937bdac7e4b5b6ba67686d289575e0ae7d6588361002790d41092;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd63c0167e5008bbea7a9f52ce6d5290ffb22c1cab4a3f6139804594;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15fcbb6af1c7171e8ebb3d61ba2d38d9ab7197cef068cbd8820908ce0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e5d6c6b6a09fce4522d5f8a7e446ce23dc5b438c9aafa82899c198e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19181c8e30eba337a85912770e51029152f4786ceb31ec650f7596958;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e357d3ec7da351977197e7e228b1d99a7f47af8057c1346a8058631;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abf65528bf2e2164aa1e89e30a960a82a1a9cb7ff69e00528b103e4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11cbe207730004b16a4e8ba3fbb69984f457dcf1a88bf7dc0415d65bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9591ae9fc6723ae9b8f005b2f1eb4d8e4f892ea295ebf0b1e00a8b69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde4136d705f2ca55712bdf1865339f192ac708a87d41830d81f9425c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df0814ac28d5a62d4ef70c97598ae7a00c1a1ed880e96eda19f9ff49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e5136dbff2de9ab799ca6afabccf4f328f181065444db3c47c5c3c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb38ea3c283c10b472f5143a9155bd1b7be217042ecc86723463fef31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125f981574deab5017a0635b473dd9cb1aec7fb8a9fd62860c4419584;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5139251588f58c447bec0013c6ce84264489ce8597a4c063470a4d2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f028fd3cb9ebe4d5868c873b8e4c0aeae49f80741be382067254680;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d0283456072e5f5064b1640ab261afc185502c21dc0751947a68984;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1030347e8385d20bceb37dc095686e72d072fabf05619c51185e9a6f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f440a58d4ae93d58cee72fd57795fc2c63785ba7f33b4c61223ae0dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcebf3607ece53fe6e4baa192c29a420254d6c579a0c35b88a3ea943b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb4781d2d0bd7af11d28ff1f2cae9192b56d6ae6ae293015e80a9b8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9546f14c803dfee60ca39020b8dd4fcc85f1a251ef8c3de10366cd83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ff595a810b5a3e5ca4dac92b5a462c79b82137495afe0537465eb45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5147284119d53c0ba482064e837361708b240766c072ca73060baee4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f3dd739510e5850a690538c2f2f2bf298e669535d1e614ed5fd8936;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h715cd3cbf7a5283f35b37c83faec2922fd69796b4e11be100e20300b;
        #1
        $finish();
    end
endmodule
