module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [28:0] src30;
    reg [27:0] src31;
    reg [26:0] src32;
    reg [25:0] src33;
    reg [24:0] src34;
    reg [23:0] src35;
    reg [22:0] src36;
    reg [21:0] src37;
    reg [20:0] src38;
    reg [19:0] src39;
    reg [18:0] src40;
    reg [17:0] src41;
    reg [16:0] src42;
    reg [15:0] src43;
    reg [14:0] src44;
    reg [13:0] src45;
    reg [12:0] src46;
    reg [11:0] src47;
    reg [10:0] src48;
    reg [9:0] src49;
    reg [8:0] src50;
    reg [7:0] src51;
    reg [6:0] src52;
    reg [5:0] src53;
    reg [4:0] src54;
    reg [3:0] src55;
    reg [2:0] src56;
    reg [1:0] src57;
    reg [0:0] src58;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [59:0] srcsum;
    wire [59:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3])<<55) + ((src56[0] + src56[1] + src56[2])<<56) + ((src57[0] + src57[1])<<57) + ((src58[0])<<58);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ab46b8ead86e13b758519979e6cdf02415638e5adfed7fe8d7d5ac835f29f29a446001ac1e62267f3605777a1c15ccd9f83eb43ca45c3a930451c75aab6e015d9080695496f6d655c7e032278c7988d48503e67b4f08bbbe44e4400ff72221b8f770bc39b23339a9c5f283639c0bb369;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd66b587eb3342114477be2072217513d85f7d44a6533cf248b6e82c3890871f5b247cc81b0d28bf1a911edb40ed35dddb35f51a4ddd089f076dd5fcd9ff1a460e4839002701c042cdd5730ead4304d4a41ab117abcaab4335d432cd038325b8359747d7f0c464a01faebcc66127deef00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc07204f1a12154294cd0b89c58299c7137294d012d639e3a6a6f010b7009f576ac7433412a6e114b6b9a2c72d6a6762dc1a90db9765689c9054e53d9cbda7dc4a0e9ae4971422cfd94fd2d10dc0f2943fade91a3b37aace8f459a596a39d66b2f3f45925abbde70a45828488b0e4e92e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebf0488913875842fb3ba061f3068650d71e44d50c43205be8cee495b7d0a7b3a69593ef713aa3d1184836cfb45b13d1bf1fa1f86ffdcae1fbc9888a49b7b5e229dd5adfc3c11d43bbba61640a0bf7d49e3ea5e5153a0faef65aab74d52a9f5f077cdd7534f234d74b77005573be87227;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd280ab10972dd4046bf629e9562d07ae036352b3f916308e41206b8e0af23b76d2a1294f399e18a1adf856c4367f7c723db4ccfed7bd266cc0a6015c76d5bbff8e7de85d06b687804fa8c12fa1a4cf9cc82813af80c3a107cdbe8cc528f1430ce99f5edaa2d949fc704d10c1b083fa0a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4667ba4e021e3b676122b25d3fe11b2b79b8316c7e24c340f40ec0d063fdba3f249cf67eb408d005cc081df39140ffa4546d40a30aca3023bb6ec3aa1974f9211a8fe50a9abcadb91dc081914d1a23f3c1ab5ff5b392123ccabe1793323b5ac256daff4023b922fd737a6eaba273c910c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f290c8047ace1fe534727c4aecbd5b27d1d9587cc1fddd69fcbbdf35715c5458384974ff47813f23d19a5c203d9736645e9f49ad5fb02309ea95ad7614005b9f6c4f94ef4430df7b19792818a29896de381b367fe8e94d2b84720c9551bc15052bfbba5588d394277a1454fc94304b46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11bf88969187466d06616566c31abd618c1b44411a592ccfb2663e19fb2315542fb1397bb006a8457afc308efd63683b1c83bba95482499d269f80bb0c07eda3fdbc5433fce43c754e68ca4bc0ac24b902e2ad931780d0407dbe1476d28016bb9eff1209e2dca209a28dd0df9ed190e1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24bb38da7126893def973ba4468a6362bce579a55d06173bde394b815f14329a9a08f89084ab14b22746b15707b4e7ae3ef4b8534124220052e2a299119c0d98c3ca37fc10f35fb95d1146f9ed0005e1cf9a7afe05b1517002fe07ae9c01964cb06329c7835976b602353e8be8752bf44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71256b80318c9c47acde03cca3e605a5d148b0e435455c330ce54d1b3e32b5797346c7c323cc4ede60db813b4a401141fe4be7f4eac1e8ae19b02df280c5fede209015421d1e19084e5cc11bf55dea2a0d4421adf81fb33edd946cc4df819a5b9a75f0c7a669ee9988a01a3049a8c9d1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37c572a3d8486908460b547b101f9121cead21b4be86acda27ce445d0e34dfb9c5c26a9e6dbddd2cbe3dcd0250ca2bd1faed8e2a666914d4a95bf8265e89c7ce516b8c84424b7ea090f1d2917d6a3a167d5518af48e48c767d5e367144681a9e55d8dc23948c9b47ddd00bdaa2108100e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdd703f0713dcaa6a5e32e2a05645659c1434023690e44c131b57b2675a6b8b89479d29447f45c95bbde49de7740fdde80f17b2b7541487b61af4b2e7020de72211d778e0f49c46acd906d8a2bbd779dc5f5d1170df730a0fcb83ff3b6d900a8a8e65cc2a18b607c5baa7437eb5aa864;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd08c3aa2c4daf39b93994198ccec1767ab05615307c6de515cf732036dcf1a157416f324e88ffa8dd382ca05c5760b8bd5e811bbd382ad7c9c8fade7ea3319d39123627a3b3e4c86eb7c7accc492b7944599dde5bdb5a70f60d2b0a61efd1efa5f508ffecbf8f99029c15993b42f0b3ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed70c80f140be20041bb92d71584fee4b73fab750e7d85f52abe66deaf93189ceb7641f0888f75add31b6b87508b3fa8d4c159c6d8ccea5145c1d27ece229746797239ffed0d0cddd1850733931d381f4bbaf1978742b1122689b15158fa1e974fc0567006eae87932b7623ac896d7209;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d85145a0ca6d3fb14a2f97d1eb0a42c799e304c4441eb8615e20401ac440c18015737e307e1658db2a73dbeaba3ff0d4630e6f32a132562e92b9ea8343294aa6161057b22cf979cfb8a38a609d561e800ab9aec3eca42290f3cce910976e09cef42f8ec84a5d37acd95c0a2cf8690fd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bd0e72c44b6f5bfcbb32ff457d8fe6c8f55e0246a678b33e1dddec86bfa315786c298f5c1ce5396789147a5a61c643370fcbada52cdd0dc95a313e01033c2eaa24f5128c92d2a5859125f84124f5f3c4ca2d11a09ee6aa9af545c508857a6a84071ca06ac1dde44e49d5cc4d185aac51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd25802806c623d0a0f4fddf29fcc5a4015577728d1afa953503d11a98dab0ed4c9e998f6ce5cc27c126e595a7a3214c4f010802060c2eaf4a635cb35cad548be4236a289384f951c9b91948676aaf27f71e7fa958f0c877ddafc871a88cfa26ecacf727431cf4fc4225552e6f0886afb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1371669e20a8da07460dad1f683b793343aecea650d0b0f7fc09f1952da34c2c5fc0ce071b475b8168e459e7e054a134c53fefaf12d3543c9b3bfcd8bdd0d81506e2f17452e3b2e1bf3729e0b6ed20c611f357c2ff36e8667eba30e66c52eed19aa57d4735793d63815955f5322d71242;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28c773759a52e634c9be67f614d7ed682b23e669355251e8b99c1ea23423d2d7e0396653f9269c196e72f04232aaa48a00b69a4974f4d99fe39575e781fdd6d28199c0a5717d2c7b9c4ebed50693b1b99c282a5dc98f49874f258bd744878fd1389851c4a0dfb3a7a32d59cec1e74d9a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32a1fafde55652b5a6bca82f331bf49560f93f7d8afe4832f04af4a2616a198b2ca1e328ceb374d27c18797d84b1dc5c34bce96e8e12372f8788b3ec40895fceed13bd216ce13e632a67a2bac8e2d760dfb476f60bb81f52183de5ce8adf8ea204b69f9bd8a0916ba426b9464c7871079;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff15cdfce59c5d4c6084419e6eda9f29703da1c1460a5e797924b90012556fa6644ed93be05049674fa9e3a6127978df7e6771fac831bd02ca5bf56367677eb009c0d582832da1cf1374ba5c7fde6ea042c37e73af6398be5d3c8772da51ba59a13554fce6912d0cba4b95f42640d2f63;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc8062fb5f96f42bd6d1a1dde477b94eced34e949e831311351112c57523ff2203aa209b6b2ba667728766034f8248ef6118d40237fe2fa310c7b1b60f70d06259ac7c73e350a7d6740cddf4f5638ef5cfa39f56422997a5d6289c91a08fea0523c41a4fff6d100a71fb06aa386a7245a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3d9df6a6a96958e75d4b4792eefa28d82fbb529df3d872c24047ed4d55775923f7a6c09a88001dae894a8c1a031144c7984bdde3d1400fd4eba988aa2d7034550e103355caa3cd787deb901f8749af2876bdbaa08b27a70dc7bc8b6a085bb7893e10fbb53270b750e2df9617397d5d02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdecf622e0f2cdbbd0a3e445bab5177b34d1ca641bc368f005743569d082d6a68e2361acd839d522a592a58c1dee3256c4f83037f7e6f3e6138c744087d1f7da4594ffd15ea620c5b9d4a4b2bb9353edc315d959626f64e5a7151d288fd8ffe338e100b0b8034e6752bff515d5beb7578;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58048221ab6cc55e7bb0fcb478fc2e6704280ed4c95b75fd0eff352d5a527b83644e0fc3fb02832aca516837ab8ad8f0bb21c91ddbac2b7799284bf82fb7e78f65a46dd3141313d597d24b525bffa2883b066ad73e6b974ec4dae3c8f42ec403ee64b96e5f21686427639147af218a7a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8428a6203485ca1dd98bf7d4767e206d7aa8e239b6848509a9f66a981dc519c8921fb3acab02aecefdbe14565839cc882d844a3a586af8cc573a6dd4d99f6d944fe834447816222dbf4c617ac27ab890f3ef17243088452510357557a6ecfadd7080d4d78dfbdfcf954554d74dbe4cd27;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h536ff2020124a74e36a27291a3343b3e286b0e9b1399b48d2c0696caa6a0ecbd16dbf1a8c2048ff17c0fd8161f3d04ce1210bf4eefe22eea1482a1c690bc2b2df07124f29ca5d87261a308cbc8984d0980eaedf71cdae52d14d2598ce375193133109ec0ee4ce8a2fb90b4a2e1f7c59f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4819081b6c1ced7a09fb010e7005a4af5ee15aad61bfa90a5faa4fdec1da0003d0f75c62ad17a3469428768ef11073edb8facb66a3e4378f2bd29b8874cbcaa3fae5a976c0ac2aa38833a36f9b57d77ce43b048b30ccd17d921aa1c3761f96cca0695bd29d6b8bf7fd8e74f3f608c77f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe21af0807d019f5637daa9b227c75e5c32352f4e847424c8f06936d1c27ba6e50cd68cbcbf05ec550876cf5cd1684fba5e8f4fc3758047f3d3836c84d7e67264e70cd0b3f477eecb4d919e8af6188dfcc9e7a247d3a9f6684d60512b173f35cd44cd53668b07768d4cd1d72fbbc9806d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2ab7d029729b1d5bbca34090797b09709d4b5660ce3fb72aad420ef88a52e1a5711513a29c0f81d1f77330cf9eb1394d37d63cefef0783b9b5d0849e15f07b6c53d5aae2d28253f8bb46fb0e79bd86560927ad24036bb5012550976e75578805ddc8049446591b90e42af9c34fcc8184;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ec801b64d81d03fd92e4d6d1a31fdfabd35c4354f87eb32b5a4bbbf3ee71869138bd9976d7dffb8add1c225200603d6cc4809f8b133f9d7a1de58cb3b690e532cb380670b82af1b33528107abd70385caac74cbcbe695259cf6360b87631c9473503d4afecbca402940fc73c6abb2e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1317654a5b7fdd6b41130012a3ee0609c79732b05a04b7be6b94a455a99c380bd1ad2ef8f0e2726ea9ddc1a25e30b4ff63a4179822a48bcf44f1c809a6e05a8c0f6304bf712bfb1cc85b052ed1f5275106bd65f3b879bbde93deb00abd7d3a1dc007702277c12c42be4eb22fd7cbd2532;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4459197d449aa27838fbe9ce1a02f94bbe4972064d1394126e0b85aa708638092d44b364bcc770a85a97d96bb3d87fcfe7a929a7910d09a47e9d5f113cd2962dca350e1e7b3e42d4f401d805230a217bb4e4f5ac5498613576a4c6353359c6bac94a9b7840c44a4bb14c5772b1942d356;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb131a739d932c88ddbf5fece3b1e2bb09207556eee2989017dd6e5e3f230b3722a725cac3fc9ed93acf4758aa2ad71dd1353ab18b6a56178fee07fd0a821b7c1e86a63115ff018d46e8788e91c32ade0da0a2e0dba417bbfe65cba72001a1b76df05ba8eea05208c5dd99d0799d02047;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfeb2505ff9269dfeea765e7746825d3fe8c09639abac6ee549a50edfe1cf334dbbff7e75f546aa3a6580dc7b6c476ee65ff1919f5bcb483a0359a950cc3d87a7a676332aac82eb2046a3ce41bd90a7792d1566c222984a7857137dad80acafbcca6bf4b7dfe8e0e07cf68a37b4dbcefd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee5baff64ab19fcfa96a401380919eb0597fbb90bafe12146552c1e8712943c04c956b614735d895bcbe71b20ae1ae553847206942385f9eb7ca15ced543622d93fcfb5e0c1f3c245e97b801cfe3f8d66bdc5f56ed1f55a8cc2dedb1ecbd5e60a784a2e0d99d77bd4e0a73198d3742768;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e7c2a46db0616acf26b0f05eb49e03761ad20b40af3c99fcf3f33accc50e28b3dcfbbae07f2a66c752c4ca34e0f7e3c6706dc7f67fed5966aff503c83175d26fb50bca9dae113213e00078b64cef5a6d01bdd31431c6f1d28f67d37f42f9138f605acbc4ca59c39289794261c9adbb5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c40145e7d420e122fb5e24a1ddc753be98139924ed7b6bf9ec1f1e253bda31684e4a8fa335a093486e2aebd72030bee228ebc46cbd3ee81177311394c2105bdce2fb2831da171369a3ae70358585290c295c9d19351e9d08156047543940314daeffbfc6eafe37d7d8beeab2e804eab5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1da6f322a9d8f6798030cf5e1624f2c96edc7b2d89eb48aac31ac8afa07116641b1ce30487b0445567db241ade3bc6094e04d5f8f5ef2c2658b479b24c29619930a39524590d6e22972734b99cf7db2fef579c21776a3ddc524f1b48ada87a83bbf5b9a44517240a42567a07cce68eec3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56ca324f22329ea43ed53399dfdffc0ab2607dda761f1e03211eefcee3927922f764bcfd06a47ff9b6f7c1185b5efd6184c486862f0faefbed51c8d99b3fba28aa96edc9d52f15932b7e4e9b624c1c71f46b0e25779f6041c77a24197560505082ffe07e175725394611dbb26b079a5fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28a4f4b628cc01e946ed1c61699a717ffc2a10cab72cbffc3392f3287435cbbb76e8d4fe189c757b780998776526e847e541cf4631eaee763c56f832cb0d75afe3c4347dc7483ce3c9ab495e79d1519f3dc8c9daaf5d62ef99a611a7575230958de9e9a30151f4bb755e352064c31104f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf25ff21e126d0842336dc68f2d0c28ec9d1e1849cf8e372bfb72b5c8ae06c310e502458ec47dbe4335224a6acfa9cc80392e5f43497b66662046420ba6c40059b14650c30e60db7e76536d11800e2716a111832509909dd3eb0a1a00957a5564437111c62229317cc84cee9b1860683dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h517a3817dfafc616d425bfb35bf7fabc2343311587fc17769f0354ec15d70b87223d334a989094e28c87bdbcd34b0583c269744e9849f7480184fa16b803d9eeba45d2216546f64ac94d51202a006bd1364bbb94d9edf4e7be8742f0d89fc02de546a7cfe774a4bcea33f62ee5bc938b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b38ea916f56a97d733f32200cb1730e165988513e696e2fcc809c83ba50073121c243f571d3d65a4a5da95d2ca05eeb11af39797bdb6c1d4a362c1342c53ddc724d1b1f4e66a88327815364f4ce00972bbb6e473062b38d54ce9396dc157a85e762bddbf7347c864a1537ced69a1f857;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h929ba4e5e3fb23db58720b4021809727985ac09e1ad893025353dd5ede7ebf96ccb92453825e946c50076fb1e90dafc96fc27f89c657baef8082bf921dbd175f59ee3c8170113260f457d04665cdce5334d3d4ce9563ee2778ab2b37a9763dde18a5d4165301965997ef80ccac0abcbc1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe98097f518f501578a9f3735be89e0a5023d463a9967d3e80330cc436bdf8a4ee23c90b05a1709231551d3bb955d22cebbfded5b3a42a4984eafe9a0f9135c21566ddd5272c5a6e6eacda4e9c84a6e89d85f94268a7c1fd70374c4ae41ac6e358349215c602cf8abb8cecb25118a12cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5b5ce5048c4312488605a2b1a34f0bf8abc1c637bd243c92bbc29e7cb7de661efde9bbb793f28295b45f395ce320bd6f8c6cd326fb5f71bdeb411df95e679fadade99f6a02461b529b3f97189cbdfa6cb7ccd1cc6b0922ef27e46658f28f011a35f851a9f9223a65eb1f7db4d265ef96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha94949434f0ed5043378497fd5c1e0498da7fe58c17acf61513e26f0e646c2b1633c7ecf1bc507f9fb2579da419b70e760e54ca988421b749d954233f3b35da139b60df02cb2075f3232db23448d50e2224626c517b6e97bf437ed03af43a0fa2d57039215001eaf598783086b341855b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb41930fdb6771d8bb2b1c6e19ad3ae8f01d22f88ea70cc21596ac326d586a8afd6b43e4d702f08922a1d0a433ecb6afd35b70eb6293d02441e200cf52269c94a4c0cd3c8e74e9995c0e48a87290ca6dbb3aa1e9816046b54208b3cc10b7dc257d04a65595674d4281a59f876f86aa2e1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he015c25c05d98ca1c70f35386658edc378a648cac3a57361667327c2f9f1aa594fe21c8e3ffb00c1e2955277004fca5b2f057d80015bcad2296d17e02b6bc9a8576d7a267eaedabe9a36fe50a392349170826744a773bff5f7c53de4404204f64cff6747100c7a4ad8d8eab018fc4bd10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2065882d533f783d70aa419965c3bc9a53415df8ff3cd32f5fbb7f1a994fbfa69bb934877939dd0958f8b3300220ce56317ca4523c1fb77e75ab2a38260f51336fbaa1db1d4fd07d61fed937d3178d37050a3699c12c05f58c9eaa6a0d71a1743db96f331712c245ade86b3c133867b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h788211730fb70e0cb6a69170ab1e1e579adbf9d950314b6cedcf1156b9461d0b3db9fea1fbb1fe076df5fc1e99fbc294dc4f6dd3d2d8dcae55796dba0055d8ce91166bf7dc503c0f556f404f7dbc6406eda7b623bdfbfb82edd7c7f8a596b7f946b28fb1317ab4db226e4240c0f771160;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h109e8523c735cb29b8a2597500b40b4457a7c8f5efc36a892487e8368f3ee3754887b648f76844b383f3775b33811aa3c166edddf1a060aca7134deb2b2f0d39a79ac6ac889fa962e8db033a5edb3ffd6ece45eaabb89e3f868a90313127599a2bff195f35d3cfadd2983627564de172e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2b2135a2c22a4de7218b7254bb640671ed3b69d595ea7acc8f434a226444bf203d55c00224d71c38fb1a5b4e8c6283a5b2f64512be69f9551b3649ed3e1a873c2841216bc75b3a48a1aef6b0644c91bc40c337b63e723e7c10d6a53874e5133e0f2d7790ee23f68cefff9cbce5e02ede;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fc0ca0d2990e17d65277509595bb3fb428869f399a1a446a674b5b57ca74497408ddfaa61b463e42232cb485c6b01907163a1e983df662bc75d413e77ba01a6199d225e7b3bc743dd050c6dec11391c3a79a38819ec58fd80973509eab317921209ad4f84d3258040ce7fe500900adcc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83d3f0b2ebd584efea70aed8251a58b31ad6b90a05713370b1c363aaf8041b349b6d070bea4fd422882c567141fe25c59ddcee2172a7fcc5e4375e0c112d77d2d22f96de7871b657053a3131bf3f7cd222974a6799b1e7f446d12f8be49d9589e440e0a3af01223bd0f13d02b23e3e722;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd704420dc202a53d0fbbb870a06a3e98b5809590618487576cb4e7c4155c0d9fd3f421846274391791eeda0e71ec63a5f420320fd4a226082ba23aaac1e69cdc028c36352fd0c1799d7a000eeb93c216cd37c9293ae6c9f43871e879fa46cd08be12b3b6e44130c28ebee388a579601d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he62e55ed15998b306393450e755f8ae28ead64e5fe4039b9a3b7f3b287cb888626d0cff82d0c03926ff98ba2630661bf860dc8034b00d55089667bd983a5882ad942eaf5d3a7497a032e7952deb1240ae9b99ba436477ad8eef46ad8a1d9af84c430bad96c972778a876e785de9e20c8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0d651e79b5458d38324ced8b417faba8ebca75e220f40f7a5414aa05d40b044a7bafe0520bf752780049601b96c8ef5eb4f3379dfd30357606d81b4e5e068fb7e6aab09da09df4c1e86febedcaf3ba31fbbd9e7bde6d3a3cb4652eb757132a6bfe1ba703dfe79cfe4be1ca6f6ee88b0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b5837b3159e3be957b1486c4f75dc30919c69ddb9ff4c0cd4890427ed5bea7fd7d16deed595f6efbc0ad1930ea1ff36f6a5d275015a8d4f132ec762c9a25b429eeb767d51ca02ddc73fc387fcce6adbb486af15c9ec8d56a268fdb0dcf1dce99064717fed4ad201b15b46d928cae14b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cc1170038f8111f9926255648a91481d7226819231f02dbecb7145f1c9f4fae38440e327facb019e2ca8f7dae2308a57900b4937dbb42f11bf0d296b7b0e8342dee20a7c442d3603c52fbdb4119838870f264260488cb61f09a76d9febe0eeb0aa687c6074ef54552ff8c983832ab4ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96175315459ede500264861e0c052a53db1c0532bbbcd0236585e2e0496cc8e40d388c8ce248d9cfc7ea8ad6b79f265af7468a611943197b1b856625571db30789ea63422cd78bce84168a7c526df1c80440e45192648b59ace58e0a17d2610e80766435e1bcf1f2a352d057f8e34771;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d4b091618283e5991dc1557b0ab75b13d5975a81f5e1af237b1ac20fef0c7f81ef0aa38db3f5511c1b581fc66e7451e19cf5c8c946c876b327f291d041f58946631b2312b091e3e3e4e6c6bd34f30bf950684b5bc5b29bab1c9f02e9c8177adfa5c2cb217ba094d1f6501c38409e49e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h784ef4d53d9081476c62c9214c0b954b031f1105a14893a6f024b1458a8e068838d74e72a772a7f35338843ebcc843adc40f154d4f81fb729d976f46fd10094760679b0da219c921d5aab9d2f9940c668be7851f24ea5faef95fdb85ed8c2ddf5509d075bcd8a5b520796b43f4ff58a51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f23d2433fa3b048712ffb40ae9e2cb0da7660fee66370ba6642c98c009a07ebde76b9fd0b8b119657f0ff007dff17882a0488c976cb2fe6135cf198005a717a118c6f3d940d088c990780e2ed34b8a2d24df11a50be253e9a42dd4ccf4cb2cf850fdce0d0f763fa78d88240d83eee284;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2102af9aba1679b801975e1dc3334670941a2c79c0db1ed8841d6c05027abb661299ac940760f8ca4f29f28ea76f89ea491e0769fa86fe9717cfe6501cbbdf1547d91b872c1d840ded6dc4d602d92c93d7c6e74ee3ed9a463daf3376b8c52a2b9605adf8c4ca8a6fcca2642a04b93e92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc136e68b42be6cee193221aa74714321e9e78d571ffa8048bc1185d4d0188c8d6a7439b5df077e93bf2697c847b49ff2a27a4714099e8b269a0ece6c8bc053cf3db74f5f235ba136206c75b255eb3fd614213a6cbf4475d860089019af4326580cf7b7e748e71bc6ae53d36b22eaaed3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha567b0111f716078e22825691838f2ff7e02d357130a6bc4dd9b4dbe13156273cec8011a2d9cdced92a047cd48c828956f371e5ffd18f1263852887826e7acf8bd013676d3e73ca0c662048465779012eed7d1d38fb0b09ab15c33867b924eb3556cbf5e3488cc8b9ac2fe15b972c6603;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14b58bba1c69b023e5d3c9af398f19b04b555d620c3e0a35f34c260c6220873741228a61e1f91a7841fbac4b170f9af3e40d7fb961e76de51efec2265d5b50e88c93cb4e0eff9b0cc99f1b760ee99acd04e2ae5c7bc58e40615a3951bd4e5031922122f933dd0b0290fbe5a758f13cb51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2642ada752c724dc7cb9f595bc676d7981e97b9f407321963a3abea17e68665462d3559846ece1f528c136d21ecfd076f7ef5dbac7ba3c0e4996f99c88f5080e45704f68925173825d2097dd2943c849ed87776cdbe7ec1a202f0c4086017ed67de85b5ab9cc446d1072ca418d8cb627;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eee0a22ee7600f6c8c7bc42df13d034faed412eed720030330bdc0670fe63e26678daa709c358c2625379209003148ec6547b36049b2d679e0084b74ee4e573dbdf72e7d8e1d4ab5f46bfdef6c09556b4bef57d0c2fc215fc87a0d8081022b2e6109e491ae8200bb4e8503fdd38aa0f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7230e0ca75bf758b5788dfd28cd29a7712e18dc6ef69494ccf5bad9755c7fe663ff5ff45b3385fd50efb118c6ac8f272271273d76eaa41975eaaf943da644d10e6c5305273becec25430feb70b0e73078e241c8a5f9e387b033de630e2476c2acfc40e3b5c503a8b6b44c5fb8ca26a40c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51d7df7260cae2a141db253ed3423961a69751513903aa0feded2ef0575c8ed0d3be9ac63406d9d56832282404af4194ea469dd7a8f3631ba02280d059cbc97eac4107306f8f406db91f78246115bc1160359a6a0eea4a209f1f6314968fe6da43bac6650e6518fb716f3bbea8e109b83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f89a0449e0f25f945a04657a2821006e25b0a9cc8994937e84eb45725e8b2e33fd4197803873d9ec639cd9c206545452e928fe02fcb13e016c185860308d9bbf415bf116055944a45b61d3c08016c72c1e61095f7f07be84446d36308951dcb28b767cd06bd2d0a7534b7128b14230c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h110ef698fd958f5141961e46f9817649fcb003415b4eeb5aedde983e3b2748ea35d816233e51c9d44c4d70bdb9084c16e011a1c9e23b2cf2aa9276114f311b0168e015dcace936c17ff3e1b01aadd4d5a66fe3e7c776095859e7289d687bfedafcd551aa5d1f9e10f9e05afa184447607;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b8fe03920b42c1e7d0c9628e019cdb0a4b02c0e34b4951dd6456ddf4f5084fa3870093d5c5fd767a66d9f5b74c5c9e50486e9ab1b3bbba80cf189ae977dde8e831a49e911f049ba52154e4d175f770c7e6008872da0deb06ce03df9c051f184b9ef197dfa3f3f01d66aa498f3f86ab2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h598a6c0f4cb37a505dec90ea3527d8cf30e3c2003a67e70b391812b69f00418ea3270e417308727cd147155529d1612a57c40144b839ff2e16e23e0e712dc101000865047a9c957d76982c948ce48f0efff3872e68f98ca89d4223f4f6a89c17e3c9b2cd6b9fbc080d48994bc311c5ec0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h351feee329c30059d129d69bab781f9094720079d76071a2edaf9442a9c05cc614d5fea83fbb16bfd72da7c5f77ac54d5e6f5f08227ea8e777918033aacf6b08da10b70493f77135675e6df45e7494c547e45e7df86574ffa71e3bda8a9f4087feb0a63827bf2bfddb0c75e537ac836b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h772564989100e320c888465db6521a15d7bac12e2a6c944c7751d247c7dda0044b2372db2f7c6979b8d73f8cb666064012ffa3a05051204b0ad47ec379df73455323b87444cd7749cd20fdb9025852196912fcff5eeb44d0d1c18a19318eca3345fb8388f14307905bbe671d3e3402439;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h134e7015c879de8fd56750f2fff1c1213ebd4a20963ad894d877622c4702a13501b37b96a3dd6415f2b63977f77c3fefe839e787be29d70e0b331f294b6cd58a3a532f22aad85e7af0bacfdb5b8ddb36ca83f4bdafd2eb0c4f33167a910c258be8cd4a6096fed09ddb077cf433f346f6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8215a0f571c1ad58e34c52a326d46e9fcc446b3e47be6d2681f1edc586f0988db382347d7139136ea2fcb07c6f4f26d831c837ae607b90210377cac28a9d3294ea3a9f4c51e7b70d05e5058bc902cedc8cfb037b60bd14e52b6fd6c4ceca7e35bc178a8faeaf5b7f20c6997d14ba5423;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e839682618351390506eb5e1c49638777601cc07e8da2d1e344bc17ce12816f03a75354fee0e9b68005117670daa8f2f1b5c86c99e70fc1c1f3ad502f0034cb0be7d13f193bb0ec9f7af430d11e3447485d1155d9f9ecb2ac4f43e229d3adfaf3176721bd0fcc4330677df301b4bfc88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c53c263df0ba672a822fe2543daa9f712de43322ead408407d5032a90fcc60d9e95dc9d8cfb095a18af6a21c1e45cd7b274cdc4abe44536d34dd96c0957de5fa8209ea3fd34b4125586520792bdc0b2c41872fbdaf9d23a9fcca286ce0b486b1d35ba8b90db731c6be69ff7af2c9b231;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7336dfb7d38e009b58bf8ea278f729cfbf8ca8db5f7f9502976359e78cb7637005f4d592415f3f79214d92faff49b67b092971346e39db8772a831368091076fd747c9b2f36aa00da160f75133cf6e3bc80d690722b647ee8dd858e7899593d55502a9a16490b5df01c52aff098f6a69e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf1cf4f59a4c8978b898d2fba18b8059f0f7f5b16ebcc54f42f8eeac26e55c3c38c9fb82c948dfba78b361c4f99fb803e15aba96355bf286d523ccfd977193d36621bf59be35fc8cb4b8ef4c57c0323a1a971ae8931ea0cf490a42e1f1dcacb09a35de62e877cd43a89909c60220e560e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6820b317b6bb0549e694a1ec8624c6305c41d8f5077913b9a357394f1be93f3900180be0fb66f7fa496f02e18d9b2443409fdfef399da95a949861b255984a4916966a8779f5b7fe9c824749a38be1717801dc91d83548bc4e1c229780e9c0f4ea84211b7065561b07b4f701d86006c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a3aa666f891ff7abec5282c32e0af2b382619bb91ee4ca3bc5d8b5f6b90547159cb0c40ac561403302142ebc7ec21ed5756ef828a6c62adf6f93eb593978fa2f27e91d67b425efce122482bc08d654078d1a2a19aee2bfdd569686c72189f0915dd50d3c2dbc9d4b09cd490f34aa92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h612e0d227b9db6333300d114f0071f72d3d06dd9334a2f75ec8d03eb2a91cec7763300ab247bce04f53f6a14f4be3be6d8751be4ae899d8e8253fb726bcc62d947c156c48451f9c7b719b681d804713b9583df0289acbfee227f682995b938b75089702c9f5c3e9132c22ad91ef10b576;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4adb342ca6d1fe899d414be756ceb8afc88c9b3596942159ca5c18826db6363b21dcf2bfb94f208ed535531fa1f7b4b48e3281174153b481b3f289d893494db59f2aa4b3c95fa0f6ab30759913bcc8b8427d02dae0bef6ed658dca0617250a8d99c2a32bc4eac4fe861cf56bbefb3d28c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbedc15dde082713368e7a89ffd182bf7d862b4a8711467fa88fc88c1b6f06e46ae75d1407b9c547befd4e8263642fe7efec330ab56fb488f58808b1a9d0f5f3d8d7befa9b2a8358e26e44819a2c8c579aac5335e5a9674004f9241d00a79c1684da6c4dce2d7c5282f194a2c45d24950a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7705befdef945121fa22ea233104216ece1d3b1149c0f603b3bd518f9546ded5d4c1a01e771161f3afda1a256e902afa1b0fe87443b4d5d37cbf017dab8d061e30f2f570118bfa9250f1876416654400191e19bbf35a0a40276958dfbf87a4456e47e7766fbe1b8687351f0bc067b5b88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb076c23ad39aa114b02d8f175dada98c18c9be8b74b14c7697c5e8576e0bbeec07b6c678685ff9c58346f1cfa63d83118d94910a5a37b97e91f0e2e9cc68d40778588f02361a8d139e81e733b5e9fa749d5dd998964eac5a34f6e24eeae17c7213cdbb58d69f4ab9aff7c5d59da93a5d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d97c66036c1b49afc89873caa05e6bb1c2e7579a9ecaa7e779caf9e19a0dcfaaef6a6b9cd78157c69dbe77c13cb8fe3f4002f88bd66aa38cab748ffd2dcb8e58af2323718b626342dbea82afde12aadb472f1a7f4053e922baa8bc33f7e97a200389cb1d80e69abf066d9ffa3f8c4b10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc69af6908b617dd6cce8b895e74f4c3898d204d65c6843cf310e7e0be277d1795ec278eeabfaa1a0e30cb6dfe07de19bdb5707eb628c1a48f70b5dce5120e2327c3e92e69b355217f0a28803373807b7dacb4a194e153bf8d88e4a09331b51de6a6f3dafc77a480a8b81216748ecfd661;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97cdb23fbd193b0af6ccd18436600bbb571aa13a9323e939932326ef961a9ec1d7a6aeb5d60136a17cd58dfc615576112dc27c8515a0d7652395d7e2f5d36c6c3051b407c6b920fc304a6d4713cebfcd0c3e3e0a4f0f13fb1dbccd2ca54cbe2277dbb977154ee28a24b4309d9c24460da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37ff4e1dc9183bbf39ad3d645ca24accd1e00ef2b40a3ee9386b587b88c6864a7f86994967e7d5111d8f325ffb0ee06857327a29daec02d9efd0d747e21a8df072564075469c7d57fbbb1404c040a62b2d79a04fae669b7fa07588c3633c0334a682ad2e1ca079842306084e4ea21e29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1f025425bcb1e1ba564bc65aa379bab8deb1ea5879b0e4e634e8263716449cc3ae99bd7762fa4aef900de4821ec74ffff21ca96ba86d65f60995a4b477e4eb04be2ea00df2ff6bd8f58e1b2c6939af6de2aebe040928e6c89273e266e19360aa013f17132f9e760a8ba2568c4ac1994d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb023a6027287b3adfe72f8b0e7ea36cbcc76d3eab93c36be3bfef58e892e1054582267407831fa2c2b00570f6aa1be2f725bbf48efa29feb580b78a7a4af27d8da4d98ec521d36584a11a33ace4ed6a19faba42e8680dedcc9150452f5e1389a542aa2a8436696289ade1022fec898563;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee5988ea1b47822419ac930ffaad98086ac01e638a48e375945bfe1434e76f9ddeb67401369b7c8bdb03bc26334910f5adff94f8bc41192aa5734f6bb5f43e846b39ad902b2ce9ffff15633544e34ad762ba46c08de0fec691c5fb85832e41a92a481b8e2d8a5ec279f2679e7fd5350f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a87fd20e501f131cd29b1df54dc02d6a35264b46ce989f982868505efb55ed1a93aeb62d91ce46054a8feb922216861425449a348f8752c88df2a3babe8048bf88e75129e4aacc2ab0423ce42c1dbc96bd8a349e1f9e85b07f06972596f903542c0a6c6e11cb69c9cf516ecc4dbd9adc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb289e654cf7b3dd2e7ddf19d1bdf321e0f09f32c9c13cb2f879f7e10e8c5061c09da4e56feff80a1266e178d566e62fcf6ee852fccaf1ec8688e1db048bc1f77b0a9068eddb1fb01840c08fd395b2bfd9f78dab08ebad0b13e4bc65f8bba6be413941513c2dceb43d6f595f86166d63a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3b6ee35c0150ddba69651f26e7f0068ededbfe95b733103bbffe20b53d0b53bea8438b2cfba16768f4f1a1fe9ba8274e342446d47f230c822a7b2bd99b252d6e8c0085873e9dcb68e67a0f9eeaa0c1aa05eb63dd074ce4d9600749058592eb6e7a562352da57f106e9b063ed1e25fab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2ded4584f056bc299975aa91c0938acbdb0ad5c1dfa870af60db676cb0da80db97dfc52e906acf3674fe4ba4591f783b89e5e04e9521112787468446382ec128b82921729211ca645f75af66fb6c7c99a4725c4dff8672821d4fd76421a04e9956a22429113f15fc7a9eb6e3cfa1db2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d5b6df0bce2d48cdf89515c9098420c417163d4f344f7923aba41b18397798e4aa4c79dd55adc9b314363b54850bf4746129aaa90ccc064623d2cabe08eb03ead1b47c020b365fde36a690b9eef7b3958a7079e90baa6539f0e94cf342929ce9566a652dd8e2ec6483de38b2f270a0b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8296854abe384e3034801841111ad54a4770a4b790130e6158c920a84956bd662f0e083e96de83220a483c235641c841e2b9438762c1d42d77d0570467e592541a3db875fb34c13c83a95b6d0f7b6114e97174260ed53b6e2aecab09e2d03445506bc50e09bb2069bf6d4f2bc0985d9a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6faa846585093f1dfc7e658d73b478d697982b7194a0b452fd2ce210a81584dce4db556c62d2511116151de44be2eb9f3be7cb6dd45ee0b8d7afb1442f6cf1047f62965a4149099e7951893617e34bbcf2e21f85287fd355d791541acc9b4333c7d599e5dcf9a6c2a8e51c561f1d83c13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h711c54d6b4045d797fcbadf5fd0ca9ea9f006d1aeef3b8d259bc48f15cc53591b5d28d6d1ec969318edeae9663dd7901bd5dcc4df168b75ded94ddd7bf370d1f126856608333239c6d6e6a6e78a7454445f5e7954980b324f58b286dca2a1d674049a69b5b42c6316f0b4d761874b7b02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c164c6f0464fb35713528ad3d91f0cf2da142639b47ea6abe584c2ad18174d59789f460effd874d9fc4b013a70c020e88a8cce5688f0288b62f6dd615b1284e389d31606f57ad2861a0f6ae505c1cd1d4ea9aa1619ba24cf7cfe51d8dea963f351447ae01118e9cf7f2e981187eff17c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5259eb421ec1669a9264d5ca33da0cfb674f9ecf0ba6f634aa65d8127f4af77cd40bafae94a5fc8f42c104bf9bb028bc408078d708cf6b23a5f9608507aff82ef9e257bd69dac0ff51fa4566ecf59b5777f05dd7ad3c2106c41117ccf9161c9e436258613f0e21aee523268029fa875d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab962e4f6922504f70ad1d2a19802620d7341b672ff53bc641aae5e01f2712f6504c73a252f491b4efe2867e83a5c9ed0fbb3bed190ee1c697623f5fd95596ad90fd9e9181a50a6f39e0d19fab004987e9a25a7ff3a87f616e1e250056bd015c8cf18fe0ddb7d8fde123f0b888bfca8eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc82d63c44512ececf78a2f2cae98a091ef21ffe710e01befefd32ecd4a412e88c6b49dfba978ba89e492ac1b9814dd803154ac7f9fbdac0195ae6e52d4287d153d38f8b90ff1d46a0db92d22fbda242ca10402ef384c8ab90335f66b13677ac2e3b8ff46df3b302dfb5a1054a044a101;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1da81da7f4e473110bdb490ed6dd5eb94c3715e361fdae655d54da5745337c97b8a4905d7d2c39ec2363cf324ccdf67a80aac62a5d02e1dc931673cee2da580b5b4a7bee252f61ece1ecb78c0ac323e251136499f03b4ec68d2e752facca10bc1742600c4d6563d4428649e56fad8ba3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde17929b5e378b796463da0997823391cf5d715694ada00c444cd809978d1039af9a1173d00a056861b7567fd82f2a781ab3c3c04bb47a7cd29e9bd0f6180a0bb54f13b77ab19f0e7b347d16fa657997a0bfd062f2f977cf979548083fe01e4287161a39a8dc0a137e02127720a16c316;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11b21cc29992765c907d13bbb3f5123eea71c0e25f65f2ef909d1a7f8f3048cde85bf88a51e7862101934b9dfe4b572f223eb0f9122499db681a6ec612918ac41019cee936fff81d41f1a358f2fd76751b90bf478c0c3bb171267b3dad0cf11d7bd6075afcce2895ca974843bcb9bd9c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he12d6dcfd2069b208c0694383ddfcfd32fd2b1adc53e3989de4bb7172fa26a527a3217386379ca0dae884cb84fe15ea7d54423ea00add1089d4a56782cd044fb2c1fdbc9704df07301c271a5d7b25981ff94c81b42343b4bb244a8245c306b8a3bc19e849a61a68f499a42a6cca9d2e10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd59fb1538d0df520a8180a4981f25a12cbb2c230fdcef4927a26c0658fdf43b393637fc8eacc90f71e50418007d2f026bfb91397dc1d933cf725f672db9f0ce52bf9c4ee9316d18abcd6d6a5d2a90d9256d146311292c2f6e8b3136c9e3be6539a4fb020335c9881e7cf63d0655bf62a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h557cf5ee57ee3183a7b0a3af04dfac3e8b47a25ac6f49c1789e4c626929ab2fdf4de61f5964d62bbaa827f81094b1765412286b2da704c4aad7df4cb6394affec1c495766f3a6ab14933b6c89582695d25592a96d6fd7e3400f20f81cf8952450f655492422236748d4890e5a6fd25e12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85da18c29f195700be0fc71de0e47e80a070ce617eb9b77096abe6fa7239865bcf9a9d84dc3b847dd4de04aab471f8693bd96e2f0e7c165837df219df1f958ada3ac9713ec17df039fcd6b7cb95974ec6d7c97e40bd48496ef36fb3b3dbd1be6611e5437b29dc300deb25eeb47a216e82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3628de7aac2dc997ea6ffc51bfe13abf20717fc80ce7e03bbf173e3e2b0d041bd908e11443a533e6d352691fd0af2b326ec4569ef03d48cda563be52fab12885cc2c41e6700f2b2dfb55336dc13e226beab0e0195e94ee54cfd549fac582cd2141275706adc2b7c87eee5e29d4479da31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedf89a694a6130619fe03c2c186910ee7380a33ceb6364773001e272ee96a6d11531d02bd78cc713be4a25621cba0133d91ea5997f2f027f8b583b0d8dba8f3a8fca0b0e6e67ab4d7bd691b418583396f58a51715b9d7c3f6ce72a9cdb047d47f7a3d1a18c362edb8f3b17fbaa25fc50d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bca237bfe7b184273ed12196396719f3768d82d6af20f72e77f79ac01693644e6dfca95b7fabfa9f9a4c2031bdfe95d845e554955ae5e93054ac690cd690f9af1968fb467aab75db38caf4e4548fffeee3e32fc68a25f5fddaa45f5f2432b7574d2c2e4b6a2b6c545e3d571024384e66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13a1ee13cc6c90c1e9d798cfe4829ad55ad1a2a9d49bbf0798a1c768a3d63d399349fd7b830d6e1993972ee46caa026d46dfd406065f3f94882b1f4181da97ec985bdbec52106391ea007345c853f3dec7cb5af6bd9183faedc8a3fb7622caf0b5b7236e4e17b3fbc1ce872c5b826000;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a7f390a8229bae78ec5b577afa8ffa146bc0913cf8edd17a923e3349e0c9401b33682071d5f9ca3cde66d41a6b68ecaa106db5f90c7aeeb739693d134870ba91904c4aee7adcca6ac705847e0d6816201fb83c3f886968968bc09a386a3febd545dd10404a4d3769fae8741efd9ec995;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd996c1a85c6a2160dd185c26d5a1f2fea20ce57f075106290c8176d16a654b5efafc379122d5f5d07c9c12475f6efd5d3c46946ba83a0d3de656a8eb376b1b36128cb37b0c396647fbb6e3b4bfbdb4c9d843a4f06f94d1e8529e08b1a07e491f8b0242cc8fdb4dc6342164218534c627e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8103a330e550f7e96121d220ddc103f88b2f55ea080ddafeab0be9561758d496195daf93e174e901f467a09ee6a25ff2f84ae0041baeefe6879c20217e3ca9bb704279f498a5c4fc2369f728722515db9380dab355758562c3792667ffb2024f34576a2f946406d563ea338e1bb3da31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91fdad1984f26c8d6f4d2d60cc5d0b78140542b073d99be11126091696e4274bf831a9ced237a5b500ce0b24cc8ed0c9bdf840e92655fa71571919eaa41efe5cfe9f5af80f53161f158210f398ffb139c1825a60a25efa949601e5d54470338cab436aec576768f856ed6e634c8e01243;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe2dab6fbca49e3c65cf41dd8feaa485e65cd7ba0a7ed7513ee0c39ca705d11d7867a626b5965dccf1f8490e8c2c04fd7e1ad383fa69862fdfafdb3302449085946af98c46d104172bd76f57f378b4619aa7ee96a4b6a186bcb8ee6cd1416cfa5f703c02da17e433f284e8abe2fcfa141;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65496baed586eb9425d0339be3a4a5bfa4dc03ee943258491838b12bc398ca7da982a2c62fa99a3c6050cf32dfc1a0b42ab9ed0942d85dd90699e37e59546537463f8d830e748d4a6191db96bb4dc327e090f9fe20c069a9c9ed874f47b5c7e7c7ca2e53c5e904d321208eba9d0c8002a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d72678e80b9c067cc4c6bc644472e15318dd98a5d77294dde2575105594c88d8fb6717424ff1a09062e0d35b7c961398c8a05258d8aab941ffc177697f5762593d2b8a510f0bc34d2b9eae21a0c8d464214daefb45082adb72dd21f85710e426b038e892eda8dd3c24316c8f99819b83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf10f55cf50d3c6bf81003dd4ce3d8ef431c763f7e9b8724b09c23bd18f68417c20a247a8b490ddc880c81bf9e7557901d4690f811be5c9a1bda7be87238be0a23984ad9b2eb31767f53ae27a6b7455e55a470c39cdeb3ce940a934862080ad12c2cd7985f61edb2541c34759a598c416b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf87ee5de1feadebf1cd70b09453da2754ec44a864a38275307df70db2d777ff0cad5d65947310ca50c31d8852320023a6790a58c9c6bbfed95d3cfa0f02a567fc2b2b394927357d5e4b9f2377c520732c0bb27c36b1f8422dbe35999c3cd727a463a0702543d4da901ff3dbcb649e2dd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h685128e1557170ae0e06a456fa520d841f2af9bbf05adacd08ebe92c521ede1c133be5e402f6df94bbcb5f8093eb7f7df3e074b97c80e3203ea1f9d084caabaaab56469d513b3b324ec56ef12f1ba1c15689d2312741b6342fc50c8a3cad59eabe95770371a724028b75b1395b0894102;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h703d434530b1d84539917fafdb7b4ef160cfcf5ccc3a9e780028a4c6430ff2cc1bf1f8da68930a8d962047971a4b6cf71daca4d2710158859f8ccfb41f570e6140a59cfe9470b99dd3fc49aad79401de476086b0aabea9e64b84cd98c948161c1fb42d723369ef0e96b83456ea0f48451;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf44b1a9c9ac1a2218534e262a2df81d9708b31d9a86c994bc3bd04527309642f4e79d9d20160bf201b7d5f28ced539058dee0d7b1233cbf406608d4c9f857c1ca8cde5137f48ed5b5d11f0bf42384359dcabff70da1f5966405069c0ae5b17f1713a9741c70e6f823036cb3167741a49;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he89dd8465cd213203552e091bb10ae4af4c2b433386109718a11eb052d4e3f46a036705a15321cb31b1c72bb55cd5a3d253426647a05f732a6af3dc2cf4242fe75e5f017c9f237247bc76394cd4635e53b191ebdd63aeadd2d2b333ae61db46b4ea09f7438eb1add994eeabb39c71b19f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84e0c92aaafe7b49a40eae633397a90cde4e8922c519acfda4f59e780388386639ab548351f9d93a90e3cec859f7953b3244cfa6b8bb8c85ce3fc098f04873d72bb55ca9f8d395247d91c1da50b4856d1edc07bc29db04a4111949600452736d36b01f1d97df675154389eeef1a84e7e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77b0ffb8772af3fbeb5b307964b8256a3843b4179bdcbd29d1cb5313a74a33b0bc7ddcf2d3c86f414a6b8645ebf5c0d1f36c9eb6da4558089bca0ae7e2543386f8c073f818bbccb52f8211ee4fe58337926663c65e552a5fde3c40d7f5a4939974aaeffeee7c6a3633aefd299915b3236;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72b77e495a8413abe39d37bc53bce87f978162c854b6708a3ba8276b4d15f16e07e6c3f56438fabe839979eb27f90e77e17e8dadf439ca0d8226d566d7f13d7bc928fa21d58ffb074dfe2ddff2ad564be73bc88fa4f48a59c22c2636044dda2b9eafa4e081ef8e663575e7bb925acbf28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fc8c1e7475948ccf0609d977cb393ace600d426f708029a1c9f85e83c4a6ae02b4e8e90850107c3ff4f0081656275347e399e68282a511cdda483ccd33bb837dfcab4e0a40e6d6e2803029f3e69bac3ac9102b584beb7b2dfc5fff58c7f6e14f8aee9a8e81f09422bf7926e2995a4c22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e91d58159f4b79254f04ee4ea47a7031875c98ab52b64c9926810c68a2b3fe4dd7ecc9c817e06c68d27660525515597f1856002ffeab92d8c163e3f80a827ec4a143d278e57120c63422f65006bb42907997bbaed1aacab43d6331b3b8b64ab02d1f45df1068c87eb88f1ba7ef469a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eecd0b7c18ac8108fbe93abc42ac5d67b93e5080bd3d0afd6fea513d4c6381c893585c4b2a0a502202762d3c64e4e4defe63cc8b5b18c5fa5a0b21d2c0ed84376ed80a293383276e251f1eb2f2bd745a52716e54314e03ff9c190e4624a9424ba12727561884c6a0d48b243c7d09a49d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h485280b785c3f9791b1e22602d98422b825ad2feb02be2a79b62b7be3fe327a8d2ed88bf8551297b466120a6cf4feaa801e98ab6ed6f219630fe4a4ae74b606eb2b8ed7bd4f998d85627581583d923696716262a856cd0d2dfd8719464788a1bf14a81d407c666eef2f6f5997d557b6cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21e9b58eb1fed98d91664d1bc8f7b67c993baed2eee112e086836d29edbf963e2dd0239e56f76438f510ebccfc37d2cf1ae5b3718df1fcc229c4cd814207ab3b0f22f3137643a0be4eeff35b7a16a4dca35044063f0d0ccc4de14d4557db39bd2a4fdc8ff9f066b78983b322e3e8bc221;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda0c764e9668c6c380ff82c8f0f76de1dca3355ef51f0ba7255c8917927da68d781df2146a61494a8af4546156d65306566852a51c9f9ad7724af483dafd20e74bbca267d585c9ef5d3080b5e89bb2267e1c590106f22eeccf144c9ff394aa87dee085d87288c0052d44bb6646cdd3112;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b3c817a36ce1272590716c3d5cf424ee94612d5ec8260887988eb8d36ea91d312fc0f1dc552f6865dc06a7343ce5f48f76e4d7ca1d8d2888f20993e1802f23e288a7a3a8a5b04f1f3c1e7e23476be2cc96ed715c8b5859619e5c33114759b825e2ec4a49e3837d4e52eed1b721cb648c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69223d3ff127ea3c7cda2a9b55b7aee4691dc1936667a1cf86891350c68c301550fccab983e9ee3901d5a22e4bc805ff1696338608f09efbdb31fce30338c87080d6fa3436b0bb1d42e747b10b9128e790f1128854b64c855fe6da30c33fb1d0a57d54e3011a79b7fbb144d71eff04739;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h415121f7031f039a2c03a8f50e95f6d5fcb720ab4adeeef971c28d459c274119352ef978e3449aee24f41978005062a0b42f3ffe20ce9d27bfee0791d5f75970cd69309ef977b77e0fd6a83e6d7d45b9d949872c684aacb6c1ff1fc4a7a947f3384300bf5b2d745646b13c50467d8e90a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha160104cd0810b9c41bf00aed15526c6500399c9e598aa95b217946b2b946cf6c4dd202fd358e50b58bec49632de35ec3c350d428b72d7b523d502548f61bc94a65af2f038652ae8df8f716e756c05eee4acb98c95dc7366c9244f320a5f564d775af99dc7064bf42a14b6801abcfdf4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6866344e347b8bfd0d427a7a9f01ea58912975b91a43ab05d940fdfc4318e8265878bdaf3ba8326c5fc7adee3d0b20476c1e47dc0276cd8ee6335ed31b961b5c7889971b6f6704b45fd2220d8cd84ca7fd216821a41e1a4722269a61692bcc912e430b7bc51a8e0ef7b10128653b3b83e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b3a0aa5ca7c2edd98bb43e505780ac4192df85be06c4cdad98c80aa60468c0a30916a96208ca0fc15da90405fa7d01d46649db7cdabe86593eca469d626d13ac182edc131e417b56325537e978efb9d75d381cb27f9acd37d45e8e996c1ff221fcb19f9beb75569c8163c1cdb02df060;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7f62063cd51a66e920607b0bc6ab94bdb085787a4ac8e526e35cfe7096f43b1a924025d60b7e1b2bf765b59db0bcde698a2327507eac116ee361fca296678b00e4103ea32fcbe3382f306fc84e91b7c8ddf60cc952857efd4912bce7dffbdaffef68ef583c1fa94b55a673a29c89e001;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h398229e2ac93a04e453031a3c8c2fda64ef6b85af61e711bb4a82ce1829b90f5ceccbe44f464dda6946dc6a2bad69261acad6b0952550ffb39cb866d915fdef3621e0de3818124fbac3e83b82148aa1e58acd89fdbb0b20e5f348122b7bedd3e79db33b4cc697f6fc59422cff186132d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2659e1eb5b1a5abebc3ec318e1a65411d7a1647b0e5b65b8b1ef7185c564ca3532f6ffb236ce1c6debd3de5a085adba262f200d6a0449778475f9ad74aaa85b273fd0dbe60521c394b5e0d4757bf3fd512ceb59689143c74399b8f75d168f9e24200645dfbcd244d0eb07a6c90053266;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6733873d12dbd69612bfd732c11172c691fea0fafdb351ebc4aa9cd817739a10da95ae607258a39f9f1b32a7c26b80352a9757351f4f00b2452c26d0bfca7a41342111a2cc6a26ebaed359e65697b33f0539bc103db42c4999ee1fbd244c38b9b30d4be1bc1fc7261a96d56ce52170876;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h622a568a4a3e57472bb45960159a7484c69e831035e9ff16a72420e881d326777580dc0384cb10a02fc4532f1d51e5ca865d9b5a07faee40922faf42394316a8da9c4eb223b638adc10cbe3221d39b58f79103e63f020d2b3b0e4ad9725ce0b012e40a92cb2a979c67dbbea8cc78b1725;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15c8ac9729345132853351be1580287c5cca827bb02b06c450d5569c36d4853c3c64887d275d133f8595226cbb90cd19c7ca348fd82aa48f7261f15f5c4a3678a8928571d4430578679d4977b813ef0d5ecc9ab24a84298775bbdc4e26c8da47c35f491b8eae2744aa478c4d5e05bec3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c5c582207e280167ec91810b646af766d92a1aaf27907e96235c730659cd70fe30bf6959df0c4e9ff50ae1ae763827ed6bd7c75495bba2290ea3a3ef0f8d3428654c79e619216ecf4d290f3ddcc5d0c32d1fa9265d0299a152488d5ebb756c30a76149f9a78f919f278a588b59d85260;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19c52bf72e5d6ebb76e3c630af2f86f9becc3696833891cd76fa8c8a0db25a13a75562fb11a234d077436e86d582995f0a381a4410808f25d2019fd1416b9c2933d916c233f73d4e594d14bb34bc3c6a46e1dcd093539a8763a2ac0b9dc3b48607b59984f1dec1c26e5a1725dfacb9cfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd630a55b79fdd648844f6c34d62e8759f73791e340ea1c4e101e1cab95307493c2b8e23893b19df57a2f292e7de328ada1b6f6257501fa276570e396c6eb0ac300b560984a63bbc8369e02814013c30e6bbc1379257280e56933f0159235daefb561f64667697d2d9936016c12e31c2ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h452968d691854f783637f896d2a9c2c2b55eb8103ec05ea561a569606b10fdb5bcf38ebc25699c1358fe4e8dc9414e818954b766502fda8763edfc1b2de0de0e7f83f21753f5ef1304d71de02a3f58af3d8f9090c17f02535bfefa0cd6e51d5701768de7474600dec3f8a48dec905e71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28c198c4215720496135fd25e5e7bfddf74521a014d4ff26b6ed0cbe5e27b7087a26e92f4c1d138519e90348b56d814023c683a6d4b43b471ad2034f4c5c0feca04c960961705dc33c129f6bbf2b5fbdce4b41d848f2882e2d205ea196c6ef7049a429e7ffbf3ad14e0bd833a1b744d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c88c2ad3acf7ee935e463e9f9c2630a67e4b314da647514e29d6ee448863e3c849237537567fc6043d2cb41b57ae0d64c30b24e4aea4fff2549e2a8d560b99e7fcad385d28aea611b355f2f72fe96ed1013720b9b0898c01278d06595f7846715a8c62dd0748e05b817b5c8378e0bfae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5726fc36cb69c0b4f256b2c948e581d562a6ce5000b432bd357da7635f6d12764b93a8cf18a03c2a919ce9c9a48fa9405b96e1d5f62ad99b1a183bbe25188bee9cdea6ce1451df1b1f7ca0159a82088e53271c1b405cae67987117e43e4fdc62b7a75a95ff1388e80b6ab3f47b9ebbff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbe5792e6a67f88a28243a3f19228ec9ecdf1675942eefa473474a818989be9a3dcff11f92f8ceedf7d6de2a1f0775ea8141b5e20c611b9049daaec1f95a824220a73f59e3705bf1a784269b864d9855deaedee29f09ad1746d8c77bb07980fd92eb7613dc0db0c6aa5db08c6bd5ad237;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b501560926ba7918f21f6db2b36956c4ce5d3c48e9d700fffc2cb26eb81503f8bcd93a52717f780f04b0771dbbcfda53332abf4e0a7747ccbf0babce018a33407cf3fb37485f729ca3cc5999db995dc6566bbf09786c9e0dc00fa4132fd5d9976461d68f76f4704eec4f4548b2bcf2f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c82bb9261faed922e010e2944484d93aee43a6068d6bf9b42315763ec67488f42b404f2b35c6d867a31a10be3d38e5d22174b7f0550fc0f4182f11ad746be513843d3dc9b520e532e51095ca5d7cb81bb289e71e61e34a55d8e4cb448f29bb7579a8e8f91a164c54085858b95fc4d8a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdad856dd44cf4062e2a5c6f4fcd5116b70e30a95c703782846db9b08f7b11fdd1f8c8f8ad7aca0e206dbd09c2851e8e379dde1b9bb590eeadb6e6aea90d444ccfdf9a436602dea672fb7595ed70406bd25a5b61d15b6eea68e95c11342d826a26a760f24ee2788fb29c73a211cdf9a255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb81f31e81b9ce6b419594589b50ac147d041355b247f2b1d3812d2ea3a9eedae341cf74d368f73ef4e9e80734e359abfa55d2f485eab166e1d2177466859d4b349747a252f82597a548a24fc24702592aca37610783fda6d7e0be7e1c4fd0cb9ddc1b346c95e4e8e54475e3a17ce1ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a4302e6dd831d574b858326c578e0ebb9ff6b1c66e5d2b79ebab4cf6704f7c799b2cc7d19ce0cc72dcd3ca3577ea080dc6ea4b604059309913034d2c96b882c95e2ae07005fb4693357e26719b32f56fa660ca23e3223988eb2fb24704cfc756da732ed86f1fe0e43bbc7a5f0e3e1880;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3615d09c9d16e3ace9a5d134e4ad5f99fbf0e5b9c0dba23b1872f3f3fb88f0eabb2ce9608151a1b4f5e81596e93387d44fde76dec7eb727256775290314479af068082ae6bc16301c0bb5aea332edd5a0c89418f5cfe83556c418f0e1f8e81ed157a3274b2f728c064d3795436fd8c788;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfd226732da123aa8c084b3fc9fecdcd5075cdc28417fed8fdf463c0df3f41496908839880878e3c9399e3397af7729a6da4f190bd571d77941cbfd06628909bc09ae78c11219b9bff886f7daa3b76cddb0a64959155977706a7de8f57cb4beabaab34b524df5a4114de95a3be317162;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h358f6a75ec6382dc78016e08806231852008eeea1bbe11132dd6ded9a87499f4194404ce608e11578f3845659038767a499770c8452e239902d8fe7ea89051766133714b4ae2c66faef36c867e9235de6b0364b760081bef920e6179ecc3f92fa6bb9a3ae11e4ff4c7ef5523968fbe6c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hede5fd8ab91de587e8b774f83b685dc4026b245ba170d01967606ff716f844b08fb241e7d135ff43e10d3468a0fe2697414a639fdbd669860dc451e50687e8c06ac21d361117aa02c0787cdf4a85733bb8d9e2013e26761dd96bacddc288b38c59530e9076d52182ea0ad85604a081155;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h637ac8fa16a73bec6f55264cc26f4949839bbc5d67a4e724541241ad4dfecccbf03aa6ed0686183b6b208a04e66cf1ff5b8ce05fc9615027e3686fbca3e63b0dddabe5aa023e5c0c20512a8b3f14f653828d022937c0a022ace9ef22d54f751369646eeb4aa550aa4a728f0882c2d86f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6df26b991fe2ffab873e866758ee3230cb31f096db4303dd48427d32fb03f6cf75702674e639a5ed54f8a6a9221654c1d4f6118b2dc338815b47b01e55f2a09db093bbfa534ccaccec733e0da734abd665d45d38a74d7c712aa1a6fe40d61e30705b7e7cadd04b08660c3013ab579d421;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cf2274f7c61a20412be5fc3fb7529c45b39c11886931fb9d5e52773171819564fd83540e537f8f7d64485a9fc47724c3794ddc110934f0e59b2ac4750fbc1a0bba2e2fad6aac3258a6912a9d9523554f1918ee9b34933ef7f1b059e020969351cdba8435021875771749e88c54b8d5ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h915d862a77cac1090461da0ed37ffdb98926a831a0001f1263df7d1104d32343d31e56b95de026b320cca7390d3f985e4a06f3830963d5ef43fc12274ce2bf16cb7b06e2b5189bd30bfd608cd5eacccd900d268bb5859c37a4aef084eb3a409f21d3588e0ac46d0bfdb1368de9651b41c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5bfa7164894ac0a50ebb21f9acc17c9fb2d21ccc5166d160b3cb23a2868929b43080b4ac910f60ca2c58c6ccf0ad09d20bbfe1d10286d27a5531f5c9b1ab0cc55dbff9467e6f5db9ed17c4911c1a55ffbdc330dfe158f3491c5b575651706e3e76cb4644f6d12c1aa244a2f893a3771c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86add21115a3c21177f1f10cd555d68d36b08175ee8b1d477749946c88548ed7e076e4140c337924e4d1a093ff19c272d29d25ce025acbf941e6dce6433b7e17a53596f41184782bf7763f0084f2c901cdab235050367590697964c953537bdb2aeba7760f9e756b2ee25d6abc27ba72d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff111c09dfb4d35af48ef05e9ec0956e4862ab232eeb2a6cddc180011eb226d112f07eca0e52f02c45259bcdd37029cabcbb1b13b30f17ac7c3e088f0320c7f5f6bdacb8927eec82b532ca11d898158c0133f551b17750338d1ec4d03c5adfed256db43348fb4beaa7c546d7ea67e46d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4718dd06a79b8f005b492fbacc2b96336929c7ddd9a939346cd55248134670538d16328977b36e1dea409198a49c6a17875e390f75aecc98fb48e4e41282ad2dbf5a18ab0f441f3ef8a87fc3c17141c0bee6864e6854b36c3e138699f7c22ae93fdc3adb7a2dde0adebe4a38ad4731f91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he805efd6ad6259f4612c9c124d79cd18a33d1b87fa8d1c579d855797187147667a91641df8e8e3b729fa92ef2cabf5cf73ed82f54be55bbbab9b9067bd240e6eea3b4c9ad1a5bf8d27bb8a5a4de2e52a325a83d9923ea8e46fb1acea621e3e106fb70eea0f41598d34483373045ae9bb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed6645fc6d05a4af4e07e76027365d4dd9357a0dbcb81d343b846fc61e506620aeb34d3b694204a22103a8426a8749bb33203c455b0b4a161e527b094eec21bb2c35c6bcf15c176e5af3e44bbb0936d74feef2f3649fb99e9a5801f5b60c2455c79fb6563cd52b73efca877a0c0249c0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9df86fd932ff2189cdcb9cdcbac70a13b9e97510736006b265249ebf6eca38aa257d99755d86984a702711c3e7bfdadf796f0c4c2224fff6f219ed6d82cc87c764f5fed2369d31a65fcdc4d5cef202d8f89a760e5d9af4073859d5371732f0b0cb9b249e8e04fab6380952a3586b75a87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41e7cbd44f5587ac12fcfea5b42c4201affe3ccb4885e0282a2aea3b2c27b12a16166d4fbd02b3f528621ebbc0a78aa8f437de0172b6910de32f00d5066ca297d5bd926cf198d1cb5864850e0a3bac7d940c83ed2884fb63fd5b44b4d4da8425dfc44e19d9fe6982c8b00337941c21cff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he67f03084fcf781af477b7d4b821fc319f73f222a8c75b89a93a237667fc36db3c6110f392835918abea076f4d3a2088de42bac85f420bc063706b457b8b88be486888a4cdd8776859f393e8de55252080c241722f0bc8fd300521be5733451ac9c7c3ef7b7ed28be907b530303b9a922;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e7a363291816889b8843577c475243f1b3dd74abe2bdc97c73d9d179348dca312f6c22721741994553995b97da963352f6c4f995d1277cb07af638018742c0afbf1ed005059497500a5d2e4bb7a6049a2237c6686c28891c18c2d2cde7d62c38060ef760358272d6671edd2434f23e81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb12e50372816265ee6abfbb2a29500bf8c3338c719415737bd02d8ae63bf1ae79c529ce00bf637fd3c1e047ee102ba6b8bb476c61d39e9d454c822d5bcf934003790e569b0b02e1a3d064bcc5fbaf944b846aabbc853855736bd2ef119b3506601693112816d8519c73d453728c918e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc829407d3a08197b26e2303f8a0908be853b0faa570cd0db20db4281cd790b9e9f517815ede04883fb58cfebc9afc1e10f62dea30e47e4d9d0d9bf2fe866e594e3ddf3932c61b417b3f77c72a95551779debbb67236163e83e1179822e89381a04f55fe3b98451820e448e47a5353ca21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e95e10db00ddd88ce158d86bc78771370a45a9b310fa30dfee9dd089eac740e15197b0218d4370fb06b7b756fd2e961d17a587a9d644ac999a1e1a3af543c404f48fa6b4633c973ca63dda0bda6d00c24c8a4b0b7f0941d12192a8a2c99f0a4c9ad79713e9d8ef6290ac08c096c2db0c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc8a5cbc245d173d29bdb81c7831edc6aa17587d8f4b0db64260e5ab692730f564e566c6e31b435e3c82f1bf06125f99568fbe14092f7a4549b40713d273826cfd9d395d6030c5193cd2f99d55e3808c625a80d36bf7714646eee4d657fadb1767836299cdb88250ccf81f65f9b743162;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5213946f4cc582b83f3a3036ba698782bf548e50a641a76fbe214700ce61f99ed7f7820929e3f5a629ea0d34929c826aa440a7e2d728734bb4ac17c87dff0885a4d4e61413b1781d552df76cbc231f0f583a06ef862238f276fa516844a4b7e74af51775da1cb5a6e270321216a1096b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3710894350cfec03fd1e6b88aa23bd18aa467a7c9a1683bf3ae46939dfc3ac7b81c49cb1735489897312f825b0d20b9450f936003079c3155600cdd5a877663f9518a844c15d880596e52c37bbf561fc8c91cb3e61cb8e1cee7cb7155fbc27ac3ac668e143f06f3be342cda64c955393b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7548c5c58cc45b44a5f77f33b4bd292cd93f49ecf66567887ba2d3c4f4bd3f9efe30e0e8d065c65dfa7a22f5ddacfc97e68b509f938d0cfe94207e7e2d21af0be3235021d1abe7593f01c0279e69b792629d9a2a9f2f2ce5d35440418e2e29d19047eafb8e552893fd5fbe29d7fb2187;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d82f263d0d9f9344febf46601d90862c250b64dedc3ddaa8a9e2d71ce7acc77ac1c75658f5d1f5b97c78ca0ee1d9c652436e469a890d5711b738e5ee6cf1e9700949f8b31375b735b265d5c1e863456046af384eb6d8df6476187a03b3a9d16bf252aabdd1e2095803d559916c602b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6ede08f91b653e821e176f3304c095e27a5872004e4da37d2ddb587811861ea4d9de90033ee2fef472ba250ece8cacd40eea7bba757343efc335275cc0ca0ae43916ab8362acccb6fd6e719c9b2c54a00f4c5d8c7f00869b32bb5907cee5130b6e96b2573afbdb233d9dca4c8c716c38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66ce4e1a498db8d51205b5a2758510a002929a6faafcd4eecbcf6a101603774727961403ddb803061071362000d2408033e153104b24abad7fa8939665a14ea7a8289db61dd25ecee48b6c7d24118a0e17b59c240de27762d1fc1bcb45037c9141a36544ea48f7cb7abbe10a957c65d40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23e7ef2c0e02efe1037040b769bb103791f9f8ae8bbc5694a2e0ed682b36ac6d65d497683be1081f3e55329fa4dd17af503cc74fc008256f982d9bd346fefc63cef90aea896459b5b6c03f6031e7ea71bb23956f907c556974e83660a3b1219e37b3a22537cc7916b98f44f8aaf10c2c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ae60b4aa127a70d4bdefa2bad2bd142abf6a6003effd46161aa4231a64c874589a8e82b2407dc8b56ba5396c585f2c6930afa7fad5dfda518fde7ea7872fce2821f512f1174706e7a585ee9fc47169eb7db59905578a64f88f985bfd47d1345227f4af998094f18e51fa23a56cd060cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8d1176b53f9e8ed9fd87ab717c9dccf27eba89c16f696126eac03fef6e791fac291312ce153952714f4633f841dda3811347c56330883354a973581681d37e7a07733f1a1a4e0928bf398ea36973891c5a705f7a203bb0e84ed0c794f2babc6087d3e39cf7bb4dbd8666ef18732bc80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he209006294675b3c0bfac539132eb3f363fc5c044fe599aab62d49f4b74eb62df4987840f346b0a30db6b633f448b7ce1de72337d2f894152d0db587938ffb9a51bd93c15adc20cf88830495baef78a241a261b82c4ab0d8ec6eec1e098d88dad8c2e4468b1d95ce2ea512584e684e9e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4987ed59467a629fb3d804d6908de6739c4492edebd2fd27cd5d90a01498c92efe478e16d00c966a41474688b092e1e7fedf94f6e288baf04d6dbd67d5e1dd61ec27394906b135658037dfce8e135c6c70315f048c262987eac229a2c309ab9b9323a6903011b2a2f46a8b9b8507c452;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58104b2f8d6570e37604cea9a4293610ae5b915b7147635ab79f1355b72d898184a32f646042bffb0cf4669aa0755a77a00661139b329497a5a5820452a07dfd528189e823f1264a16b33bbe60e3a39be6ec70a12318c08ca19fc776df93c8ecd24c5afc50977813cb6e19fbefb3a675;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b4cda2b465a3a77101b5547bcaae79a00caaa195bc5a130434be313acf1377dbe74effa4d3a5516bbf80b6f35dcdcb254c32f73934f8bacaa51fc1d40a493f90000da1924a31e803ae17cf5ff374668eab5b253d8bad26afbad21804f79d8d5cd6e097091428943a945782ef9047c02f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca360eb42112b880579efdcb7dc02cf546b9868ac13e6f5bf17f5c9c35c31b8288f0775d353eebd30252e4fde01da63c4054bc1e272a5c3a07c670fe9d4e7052a419cc80822eb325f8ef4d05cfc9d4455a10d85b1a9dd3c5fb2866b3520b836f60431dc7500b66c23d2ebe69a9c22dce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1eb3c00e306edde7ea98f2e9b932cc085f0875339e5a1d14c6e75364163999b91c0f27a367c27f2683e93dcc4333f40d716f780606a0bf1e85fedd6935b791d83f55fa9f47efd50bc1c15e5503d78a86259d0fd805ef4c2643518c0ca76e0420817ad4421d4dbc8e3eff1718da11aef79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb094dc3c152bf0f5f12db13f3ad479a694720fd82ed466b98f838f48654337445fa463bbc72bf3424aac57f8f79a1432a64fe8c50f406c86313ee2cb93b6b279134db41c02f66381ab69726740fe366726560d673d2f69e7c095b90403509aa7c5718872820c932c3bf91f3f28763d512;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h681893c97e960d2d1bba88a24f60809c59b43aa966e44fa8ab4ae99a6eb4d28757e3bcb3b172e079a4bd1f1e33dd1348d63910f553db3dee3e287963bd596f1a0ebdcadd25d90d1f5e41a178a2b27415ad7ccdae87e3cbb3fcc037883782fe0b8e53c7767536366a5c44aaaef8cdc7ee6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1da9251644c9d50463a7d1a3999c50830308bff0db39c4ba366603595ae46ea3a4361fc764dab7c54ff3edb16fbbbb8c9381f9a6eea80f0e2eb9b4fc453f93cc8682bbba450f761c8083dba31f8038b5fca0e2e7e370e99eb4c334f0ee3f7880f2bdf9acb132fe7ccd699fe838346418;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf89041883dff7750b33185d1113fdf96c49b96e444e905edf6d412b6f47badeb849fe26e6c57e1161589b877590f29752c1ce5f9aa21b68a4ca965195e937a62a271ceec690f50d6e5a05c87bcc4cb84462e598f76bcdb56b63f200ad33c33cf5b229c83d43afcb9fcbda67f8409f0217;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29df9eba8c68861183f76582c881457d88776bc2fab1ab5a80a0d285cc8ebf7edf5968cbd9de909be85fe2b8a24587e66efa14769596453ae68d38ffab8dc2371ad5bf5ca9c18ac409dfe1b9f33d16adb8870131512fa9edde9fb017bf812edb0e70ff4042a80408301262110bcb7f966;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8100f2af15aca01ff04c12d46b723fcdf69751e0d31a6ad6e380bfcfa0e41ed4dc06539c6bc34a83ef65621b5be01f31b48e92a7281b579741dea105d503a3dcc641dc51a1321f6558e5d5a8fd27330195717501f8f74fd45aaf2d9bfe916c56b8ea1c3afcaf59c30e8f5e5fc550bd4e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7cb06e58d188f457dbfcdbcdad1fe1ccf120c3d7796e9aceca96a54b0a97b12f7a5fcec30c9a7ad9d325a4c72af93c64795cc50f67589feff9198286eab9c18cad5c697cd2f35e73a76a9cd8967c3c09ca5dcb91b7bf7d5f54aaaae180449751816e19f482f38f9089ff99970c40c79c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h952e6758870df17feb8db4482daaf8f7203152e9914bfaafc0dd7218e0671f1a73b9c60bc225d1e705c6a81df634a463f5e878567343e6653a334fe68fd71c8da9b47cc7f012073b1f76188d2e2a97c64dc9549221c60b96bf61ca79970788eae1ee530d3e465d332a4c165c0d0b05cd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10cc9bfb4b56897dfe4c0a2d87baa6ad147a32629caa8bd0979789aef1b9c448f68aeb89418e00b6d517cbb991577239c30faa1211769b8afc024832e1db44bcd1086b60c2093553117a15e5bbb7d7737512a13002a6a67df85e6689aadb354e39ea79ffa0fe49caabc07c19eb5b9a32b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aea5345495890a5a70b43bb40677b865c7a6cba11c181a017502b781dc4ff6438ca3ca6336b047225859ed0a6261508d01ebc1d0e0ff233fdce7e683a68e91e7393247e8cf0034abc3b32d7b5ab5e749fc957db5e71ce13fb4b389fa916fa1840963f3494488fe3a05d9f89cb81a798a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbc3ed474417a8031d23ffccc9558f8b2a7406735411e54f352ce1487e1adcfd66481138d2b24b3926ba56fc519bce83b3312f41628f0e56ba11d689ae2089d169ae2b0dfba4808ed7d3a8df411d3355b4843380533d18e440ca9251c1cd87a2d4870f3e159252012a4dc5b64c8481c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h675d8ddc8611682910384eb1f7fcf8dac5b81ead95400099b7bf7801056346d41ad790428e4c5965489c8ae087098c966e91a4edef80b205b32f30bf4dcd7458d1314554d9d2ffa915fd779a314e58ba3c30bbd2cc016e7513f2854c4dad9b4654f4e49b8635dc2cf8a870a740d6d1c65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8607f6d76a34d35ef86421cede4a8c72558831708a16957aed7959e31767acdbfca4c8e0d232491aadc57997abb8a8780a6827b1082ae6a6501be7a995906f046cc5875a7622a85ecf8212865b212a8d5305aa0e86a36a3c61c43fba7793b1c579a5a0364953172cb66634203cd93ebcc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21260e29fd93a2bc70a8f05e44766d5ac692c3ecf064669bb1f5c5b989d5b678759b4bc6f287c40a09f6aeac2186c4aad0d7701f8c506508cda3b2b753173a491a33d5039fc12cf45e2911dc412449957dcff124662ae0bfc0415fe01cce1dcf0414ae7287c02abc46291131e9a36b173;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedb8dd4583c5e242ae1b3255d08408bf3a0d8818487050144ace9f291c2ca997e0a48dbbeed670648b0d4163f10b63c59efcf440c660f9ac3ccdbef2e1bfa4a5d8fca77ab85c27b256110d3a59b664d79ddb3ecfd65694905615531e8d92f5a78c4cf1c1036d9e78bc7e38d599615bddd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h611a95f6551ae70ca1aa30a48fce7cc91a4a5966048613511fdfaf88224ad8ee7f7fe1b3681bb9d211e59d87ff5bac25f296300a530f2ffa47dee369c8075713fb7db8093778173ec068e90cd11ea884e877e1b6d10ce22f697ef3aad45db26c64010498e7ff1cd51da83a26a33c7b6e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb068325febbdc507a2fee004f0dd95270214b6d5c17336491af3498e57b6f46370f20b4101f8b46fc1ea83743105cb163ce9de29737d3557793d44a8f2031c581cc153cc4057742b69d5f63ef5d0b4de3857935bf2181160ea233fdebae2fb4170b57df2e5b0b170d81442bd79707ecc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf082dd99a08c18be960725f635b984a58bfd10c2be0ac8a975ecb5a3ab4077a3a357dfb8837c96b10aa5bde747fb9a564176a14371a8f332ec5ab80252ec2ec228bd33240ed92d97c9b8884bb0b42d48b9bfa546be31adb6129c4c304880b5bfd9bb41d882c85dd72d72a70f41e081e80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1d95ce319a85fc04dea2186b2ff15dccce8c70fc463f0eafc041c5db6623a0db2d8056efbecc9b9f6dfe1855735e6ba04799d26028c001a9e2921e3bec429264f95adef19be340529eb7a3827533fdd1407579296a14144d0df68940299ccee4e3ce164a6f4a157cbe2d0bb7b95d061d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd033b8402514276d8cd95e69c8a6efe7a164ba5b3964712234ca9ea4e8d7f90bbb4d5dd27d9adc538e091a06ea03e761f8d58d101340285185f0499376aea181bda9ac6dd45a272aa98164ff6b11d508983f9c77224f50e3a5b7274e98367e49fe20d4ab20ab4c68811dce7b83c2ae61c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40f67ded910f68278cfcbc225776616a0673a5713122dbb4b4936e2676da0cd61383c4b567ccf9d7b856cbe5c192d2477232cc481a903c675dc6919302792d2e67da4b50ace3a4363052324118806722959343a6aecff8003dd7dc72f15f76d408e3e7d5b92ea49efa07fa4aaaeedbcab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf06a18e215a81afe5ec3a9a7acffe7c63ce1c45883afea312dc20be29a664bea40dc5e88f1130bdfcc898cb7cb74100fde5e1cbaee7543de7c9d2b3a6481fe01ab0f55ad745b476ea19e4003d1c1da1e9fb3de4f1d5c09a5b3ce20c8389b9c850a0eb46eac23e1fd0a739eed84d491624;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f0826a5edfba60f33d5298ff903e4bb38f9cb985e1ed6ff7e66782ab020778991818d26e3059e416f8c924087585116e99c97a130b66aa299fd4c3b0dbc3e689735c7a18d074f482b67ec07fa214ca566e756847ade4504b62dbee06555b1da4ddede79f95ccbbb7a518b928578533b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1567dffb8975cbd743fa9cfa7dac901bae939259520f7ca67535e821a4537b2c2f98c173f8e87e8f79a10d5cfc0960814efe3a0d3e6ea0b8533a7eed70dc9a8eb51e1a29831e8d986cd4a681a5ce270e140eedeb3c88f8e676d3a1da8c3c3b67cdb5cb8a6143efdbd71066df887677f39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ffa9222aec1c6ddcd93f3a21481abf7af84dc4bd1ad30ec673044e10c78d2a802a2d483b806e2786c2970100bef927fcb4d20267d0ce17537e96aa8ab7ec1b798ab76b28ce21595de94ccb3a2b5fbb7875d6e2eaa2241bcb2a67ec2f7b8cc98591540aa756f0e89075fa928154ced77b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78e25bb78409b1917b0be6e3b18484392593688dbf8a99de18f2bbe50faa9e4cda9db57347ffdf01b65e73be01b190817c9324e98d50426ede2af9b5b31616e4494b4e2d580771648b2d7f0accfd20850e78f83adcad315e5c6c4ce1e8a5debfa8232e0a5d67e25812109273c7f231f49;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86ec5fcef1e78cb4c5ecf5eeba1c56a574a9808f4eb317a5492fb7f5c27d1579fb97901f3a82d7c23e4a385f5c9192a9f1e7542b7ac1766ee7649dc0c8b59b322ff97df58a0ea79c62654b8db49a9e8feb1e0a810d743f494ca64820c81df3733cbc24d02ba686089db9bc39f1891a7b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf07e34add119fd7387dc29ee928084ddd5f3d1408456a7a5fecd68a0cbeb5883c70803a3cfb11eb0bb6eb81130e9a5c73f06da73d8f1332516a31a214d532b28afd80dde412cb964ea24083afbc32a0a508863650d10b3cca23a078ac93318279b45f1827cd22246477be0e541b08142f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4f0395a4832aba1bcb3ddfb0107da3875b1a6da5bbfe00421dbfb38c18da6a6247f2b1961b336902e8e3ab94b7d70f8028808d4f953a7274c6b0104b131f0c8dbfc2ef1fb03d113785e1f8e060b7bf3c2243439a1de35f869c37d372d8a34da59c4f16500bb50be94007b65f141cbaaf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8132bcd136610510bad20c6c709530fca74b2d5fa346d3d5697da2febed014e16ae0050c6da3fd08de69e66b6dbd286be5ec4340200a25d494d3c1e9c1ca131475aee254666b4c2e39a4533f19237c6512ac2cee2a5aef061f366720bb341f05261fb2f001bba04fb61d6823f5c9b78a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e154458e6780633cdbdeb5952e8c68d0ec4ac8389951e443793d14de884c7e0cc39dca779bd1f6f2c9e9af6387219de48c921f276acc2e0d623ceb6cec2ad9a244dbdcecc0098eb456ca66e05d8b3642795a36b4836818836c4b2c56387af544ba95efcb845be0bf09a5cf81596fc5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76c7e25272c0a1ed9054bb9e89819f9008b66dcada0d87618be653a35f2b2b538c2d51f6e5ce363b0d7668d54ff5a5db53e2c306af5bf088f31ab069bcf60a705700cd6ae214aab372b3e1f353ef44491580b9f6d4a817802d20add49f0d60b8c55d5e9df6083136fb3d6326a3901f155;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76eda7b9aeacb9d9471623dc42c475615931fff7a173e438fcf21c87140e596a53754082e32ded6207a72e649aa6dd0acf1eb42327c4d1091359dd081f1e99eed855095f0e715b352492e4247844e092ecde94119b9aed16c875636dd0933818cdf2deef24aed2499ea67926cc8cb6d83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed3c40747434efecb57fb9ab233fc026a8a6682eef720b78686a4c63b2b075e0f050e21051cd515e894e2855b768e3c37603a46cccb780e0e7c1a04769f0edde55de62ab2c59bd19763d169223937cbf969eb31db2ff791cf934cfe9b20b01eede10d97fce387da9b701c1da36821b9eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf767569e7a25d060aa20199a5182087586c3cf72fe801209af8fe3547be6861a00a1edf0b3f659a95f8c64642592053e3c8b2f35366530e63772aa3c3c2089aae1a69e52865285df4d76876979f7367596a564f13ce801c1e8ac8cef9d53fae979b61711b653777e1724b145c3df731a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7edc7ef20724f0107f93c8af173af4fbb6e64bddd1d07bd5d983e7644092c34d51479fe67cfd458e624fa2138435f1b4d52ad2f1ccd282b1b9f5e03700f95497b46c90956b6c8cef6166652672840b0ca867d04349a73e835097f246186cd0a51a0810838f5b06351f7d6759cfd0cc74f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7f3a0c22ec0f66cd5c947058eb5ef45b7cc226d6e6812a8c30d9b3dc0e890b3fd501f771e403211a6125963db44681ee7ca8f058a1ecbe24849c34f9d8a842974b552529f19b125679a76eaaa4eb4c5f872f577c85599e92e6dc654c8da515214861510d0c4769c775c5a547f2a3852c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbf159af01f4437425c6fb1dc610d6169a6dfbaaafddd7f70390236b6149da751fe8545c73f51143daeff31d8eacc47e10d9c2b629e1cf0cb2a4d740d49d2e040a7dbae0d805c90df6902b5ddc51950905dc547f11bd6dca03b3acea098e8ec38413a6cf3d79db19a540577d2ccd9fa36;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb6783b84e2b316824b1450a9e2816d63a4fdf8eab191f846193ab552e94d0ee35e8503a8e7b429a72f64fb0de3a90ee3493576bb61bacf705e78b920c2fcdd8384c62722f1c2defc4d631d617c484fcefbada33062e7b53e08e95314996fa6c97d88b52f6da17d20a07b84f764c08a24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc316be757ad3a7cb62ae142710f220f3c39b681e3eea23b6e39ccd9091f8a2a3e73b6fe2cbadba7a74505cd70e2b653a4b0cca7152fe8bb29727cf4a1f149fb061d55f7cf548850700da7c44481919e21f08d10d81dfffce980f21b37bdc4e37a5a6bd01523a22ca352040ec75ffd2f84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53cd63ff983b72ef71787de6de8c5dbc3ee78d4558dd926cb099ca0c1635b619003c30e45d23cdd89255929a11978abc1a364d81811e16b20428646c611f01c8087c145de7cf6646fe68f9200103fda90c9d8321df9cfdaf74325215f0bfd0defccc64506ec7943cb4c5e982654c9ea8d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h998b469b45c360b033a7fdf998a4122ef1493144958324f2e3bf0bf9efc5b87922eb1ec4be049cfa62365c802bdab5144e5215204eb5ea329de50d96ec146392a872d02b4397803cf59fcba79694106f41fedd3581cd8631b4a9283a62f0e6773b0c0d7a2fdfd32f964bbca8ae89968b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8549c3b9b0642c602ad62c994c4994e0ac58c3b6a52355e4e995eff196087c924f7ef083087cc904d6cee232d005d5eef1fa8bc48965b6614d546c5f1d443b52fa9945011a7b44b406dd02f17c2dd3549a7bce33347f760a8789ea7f5c7cea55af03a32b98a8b51a43ac7bf396fdc4a22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba944939af4129010a17caf40949bc7cb30618b6e93ef46aaa0714d71902b1c395b18d0a971fc74467ccee579a40a0448e0046c1fbb1f446a01e6ed676df39ff30bb047e9586be44ab863fb0ccabef1ea0f986f34524fd080143fa92d0c2d0c914098099d6724ece31e8a0aa63116428a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26e85cd722193945d4b7e9d05a444106ac62969594ccd06a9db51671c5b276680e3bbfc7f8f5756cfdae67b1a97662fe1e2919e9b79af86f9cb10765cb870e361765da015d5c00a80ffd27f703ea5ee2aca387fe2689aaef21fbe4bc26f034dc8eb78f1bb1380eac5e7d620ffc71f3cf9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc85de3cd79c9eddc0d46194aad079ed26876e92867655446fcf3b9975a17fed4eabcff9eebbd8508ad4cd19a2f04c35b39fcc582fb7506e6c660eb8e2b3c83f859501fabccb8dec96aa592c5a257716668a8a6ec55e2a4c36ec5f147883cd3326fd4b0a46c486157efc6713846b417ea2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53e810827020917c9e5d802c2e72be61562c03590a6eb71b8e6bdc4952fd5509b2fdd9485f338a68de69cef2479466c1f986879ae4f0b75b2600660723caa6dcfb40f3cef2412b73b71cb4318a13b7406ef75ccab7d6d701d490653acee8f19a242a293364139058ef1d61cc62f4e3c86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2951834df1e78aea329b9cc28c1d7f6a0954c46f04ac393c9c6cbfa4e550310102c9acc050f07c6bc5ab80eec58d2d559ac592f06fdcf70fd117d1b68444f73b19868f624480e8f50c45483fa631b01e7f08857ba9b64fb4dadd750e89f047de4fa550b045df0643fc3081720eb23328;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86349210464dd3a79915cdbff8c23eaeba59f984a260cdd60c20720170428577ee897633455e907a9008aa0b770d912f8002209e712d94426d40f89088280652c1931e9d233ec4c9e2ae9f808083bfb9868ee95dcb5e5a92d9d27fb7212cd65c113df89572932ee164e4ef2341fa2425;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37674d185d1f280efb368461d2b7055ed14d6a847b9a823e8e15c4af0ebb2167d541db588cc60e5c420e8b797d457b599c80152b8aa995d3b50f284b6945355d0fb536cdc3fbe52f1f4100059cf4af39a11277e4bd7c16fb9924e9641afba336b135c227f7e14b2e0b1c6c323ab8623f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83d8312d857ebeb72cb93daef20d9275f8d85fe835ad12f2de88b7c36043ce43691f7cdd38649c4d7babda2581782873cfe80f5adb4fd75d382201e3eacb49f3d0517bacb8b016a9eba4869be85d4f5c8850dc265ff710fcbed3949caa04d068312b18d50984eb0df6e5d1ef881db54d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11051e8db8f960f4fad87b2d62bd26a3679833c5a5b181f9729e34f1a0befaa3fb28395caac86deec8f3bc91602b3ef9d5f1e9ffd5dfee224eafe42e368ab977ff2ca759e8747f22cdfe97f761b4621690a3f245e503da2c2157c84cbbe4e0b376345013bf595d6c86587ac4c977460c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1677c9c9ad89d67813202265797e2678a3a362c896eaa7cd1a450c073f83ce369cc21c76968434fa684df2eeef2f253af3886cf9e42f6c97bdd9250fb774c7693048856caa556a52270e40ae086ebacaa4cf427867abe8b22fd1a70cb9b8812c11fab86dd79b7c9be6be5112d41b50966;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9fb77943255f4026d4edc1b934486dd7bff803412a2c1f2f703f58e02261e77b04bc2ce4f5d6c5c22651b71b3fedac53851c6469350061d6abfcd3691889c9a4f6ab33f30d40b7ea6f03a8b38440e497dd17f7b7cb9efe6a5c44b8f99aede0b016c7efa93622072e838f1d6235d748a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd541d442064c48c183e8a17635236d7413addce3c01df0f0c4bf37ce1ccd976f3d831ec28ca4a78491e3270dfae59984e0878e52ef824d326cb18211ecbf4c17ff47c36fbd5625fcdb17cb80cc61eb96c693c5bd7309b069b18dec3854e5d25ebf6f02e714155e6bfae30a2a82b13f16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ace10609f55731514033b0ce54f56a739c990e2cfdd66243412327abefacd96667e47d2c38ea05c2153367ab2de56e7ba6fb7cd9d6ec5504bca6e163f73f3e3399cb8fa25c45f0e14d2222b807502d397f37f1e533b990f0209d34897e9e86c04b8452e4f36965c4b4e62bd8dd4d5751;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h284f32dd73298a1c7eb8e05e534173008f874a746db5f5c242c7f33fc8a27c892a1c65145be99141882cfe14a6d433086248bb74fe630c05d6eceaf57880193914caa815f35de5edc73dfe5d3a79f4c2a38c0aea122f969b794b327984191c2c430087182280713a07ced2db64ed5518;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7b14e8bc74133045ee5f94069507027304cf3e6958bfd85759e8b70b4eb42dbcfcb6324bfc4ec36b67b5a6ecfa2f0f18363a193e13eb61e6dff2fb137acadfc46c26921881c3339048570ba126d3ce19ba10f53d4ff0881683e7de67f09f525b7887bb4ef48da2bbf7ec6cbe72014b48;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c92280b2086ca9bf43b0465b08314d9a68b7530065494cf844da032ef4a882e01e0e056bab53c93193c94296075d5604f10ecdebbea9791982a6716d8ebaa325bc8d6107f4728e6ee6f046f7300af096f4941bcd34d168c1a76b01bc57dbf4b3dd344383b96aa4a3350b863fd7514a24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a89d94d176a7f1f214cf1b5459842544e1d8624334eb71ac16b3e519f924e450b00f127d0da63eaaf2668c1784d95a2eb0eecd5deb36f26e636410c6901936144cdff17307d2c90cd8ed63c0398569db9217204c3b696c581fd543a4db2ce521454ab64ea23ebd1e99b155da839157d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90b0551ff0d666f5ee447de503645b5269b3282909a0baf27e0a09241924041277aa41c511259009e3ef0e0f876a6d5072a51521aebce85d3ca51490d0bca5f2ff7c7066f4b19d2b34d024ce1757247c2ff8c26198cfe0c24876ef9ae81f071d687de65b88396f5ae653b2383ec8481f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c12abc8d265382382c018a15aa51f846a27d91dbeb3cae1fe470f57259115a62fa6f75bebadf2d71ae3e0cb8a2351d6478c8a5f7ec3c071cca1a879f1c727b979c5d9a67d0d458460d3d9290070a0acedbb3294956349b518d168817619dc840e3f1f6d4886c274a794b66893675ba2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd77fe600d0b2f73575dab2885a19d13e9e287112b7bb84f2d5b9bc047a2b6e6427f8d498b771de4328217a8723048ea9309145928ab1e5fdcfc771bf9df9c7cd01eb5a1846383ae7882380d053355e96920a12924c6be689921838c5a953c673503699026df7e312873ffdee95bc661e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h630f1cf2868d91721c8df86d30d563f3b947df08a1bce8f17f3e4a7c98a7cb0489ff586462cfc630db193440a13976e532ba7438d3b989ef1eb14ea91470bb537b2293ad3eccf9dbc87a43ce7752fd1c2c2f781fd85a3eb612a79da0f6a0d4888dce82f28e27079b8539cfe23018388a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2f80884bf8bc00fe9fb8b710e220db6fa5278e9528695f99e320f0e32617bcddf6554b0f2f835e6a3bf670cb16263d5c408bb060480ef3d930014288749141631eda8270bba2065e84faeaba2303df7beb72bec0fbe3abd8d54984f018846c548a1a65f2e30c8804db564bd5af6e83a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b564ddd6b0e78dcb419e63c8ed014c0aea8d626d669df55ccfdb646fcbd71a38b82859cfba265925f187f03ee8b28e21528ae020504b8881730db37919ba743e9155a60b52712cf48b8cb60e593ae70e34d3304a468544cc7650c218b6b1e4c40b3bf0cf72a193fe4a86c771c13a1b85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac1b08427de15d1914a744178b584c66b34e79c00e2818405309cdfd0d9fe10bbb0581cf446f2b98e74d1eb6c5ea22f449532673c96931a792536710d876229f97a5ab35c6ac350fe913d24f6d82450841aefcdd69c49ed37db4ce7e30bc40669e31a28c9c1734d835c2ee286c36d04eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc484a0b373cef0d6667d59c05949edc198f1eb5a39094ef0800d9f5ffd9879897c5f36efa4e9e9cc78c42dd42ce193c1f46895566f039ebac5636b03bea6b310a08e7c21464a24cf0d1fe49a8e026f22875b6effd790b691029cc95d8c289dfe9f33fcacb617b8252d82b36deae4f1da4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcb9ab43efbb5dc953410177fd77b1cfb841fe696217e7133096bce7d896d28d001e735393c599d0096ef259723687fcf75c43ad3d9d2686a4441b1033240bd178971077d4bbcc820d7db73297609abb5831be1f19fcccd371353cd1316abc2bd5078bb88a2d952c5d55bef2d0e24996c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0d5dbfe7a83d4634d25937a920886397a69b692a26eea27ee202674f95546c092f77f12467c1c0dcb0f11e6919e008ddbbedbec85e3176f837d9ca88fbfc1ae3832580b686a8832ee581d27d0569a21586e7f0df640a75da09f34f6e615ce06e135fcaeb74393ce5063d390dbe420b87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15aee3c26b72ffb836f2706a13f8d59fca5d6fabb19db8f8d69bcdf205314b00975875258b1fbe2be0aeb12651c93947c3e642f2010090a1068a9fecef29c0d397469d8a8d995df1e07619d53e6f7af0862152a70f7c4d42ef93daecdfecc3f89fc91d9001def20933362df26d0038f7a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16e2914025a21f72ab0a801f86b7124d849d2127ab8e56fec347ff4ddbaed517a9ca8f82cdc663c1ff8c9d1a1b8892b0a722c352627df8cfa1b0facc0bb2523ae4f09f4edb35f23259098594fa28aa24e38b71cf08db43638743f336818dda1a802550814d57e1d2ef6cd498fe069459e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f5f7f6da3ae5ed4391eb186743aefe5450e509ad8fade13743cc8e507f267a12e60616f7caeeedca9c7e7600e7fe146eaf3d997939d2846dc38f8d21bb9d34aabafee3ac1502c264a5542f6c5802f498ec7a68553e8da2fa6b60e552ce0fa66140958d49cbf5e6cfc59b0be39010e321;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2bd3128ab8ab600ed05fd92bd442f5b3d93ee0b51c156b848244c076d85850504cdf3b7276ba0268aa4e7ed38dfe52df139368a713bb0ff593b0f085aa6b3350087c4f26927aa491034826f332389bcdec4735c7d39bbd816e3a7c5924270a4fe849b3ab71311c2292ef11075f9847c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47ba1dcce413912a037726205866c1e5d5eab3140731e035dbefc8e504a25a7d353e35c25956a6075c5b3ecae94c79fd0d28eed7c6e5ef282c19ab61cb5efe928d44df566453cbc1dd7ee3b4733808a6ecb762da3cfa864917b2d078a0f05d3f4535c07f41102ff02d6f05093edaf6f91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1077dbbf8465b8152fdb48f3372018a20a164205b45f056f246d0cf5a3e3100ea7c1086b6365aa3f8b542fc83fbf2a6e0f6a96e53e6f32fb913e2441e8fbf3ef926f95b3a333561559822a9bfdd19df8edb142c4e4465ccfaf499ded8d7f9d10dfb23f851fdf93239e23d8596a4c231d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf94e42eb828c21d86f19e4173c3ef9e063f65fe8e05fbdf992b7bfd1fbb961f1eb4f41ca82257ec6ad203dcd956352410ad3ac3e2f3521d9075326e0cd9353572bb110fd3befdb5cb4dd361b7042e53de52ce0bdbdad3fabc6910665d369a1208a36b08ccbdd95bbdd0a2ef7cba80d3ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbda3036a3033436c45b5aba3ad21134647b284a24d36e301bbb3d34f33331e4fbafee2ff1d814bf7b285aa5269f67214976ca7a818b4896c77ac1299045ec6b0b2f5d7dbc4624f9e104811ca20433cd5d871f4addfcd9782adbc27b4a2eee81a217e14724fb6508e1d849a0678b283495;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82e4610e017caa2303d13aae6bbd6430380c50017cd626676f163fa7d9e06259423eecf4d8e187219383b988de6521575166703fc022d9e1593dfa2d3162e2b22515aece9d7e9e41b51abdfabb5167d0c3423f7f83c4a73609ac7fb1610abec7b1852f5c2674a4f9a2e4d3f8e1697ede6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2da135450475ddd05cd24239e72c4cdc0e564e00cd149a31607c0ce1b509bc33a158837ef2d9ed602581b4fc2c9f3e3d98453d080860cfdeb4af2192eaf273deb28415a7a5c4fafa42d54e3b6de5c401301a3b2e10bdb1b94f8df4ee0db93cc2fb4713a569607dd9095f27113fadee8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5f2f11dc948b8c194e3f688c5f59d1a5e244b9b157e669a003c2aad78e0a25cd68ddb424a19c3fcf52669459b98bc96f7add94d758661898f8d473da612568ffbc2c225fafd3f9eedc9a608e8727ec5e61731d38d1d848ea21f0a4e22d8e2f2d0de5f891aa057c276bda2c4d0e250059;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d0d8b726053758200efe7f81e8f52226c5b14778335497a1c837ccaa476316960eb3a456a28d6fbd3a9419746972efa95fff5ca1a35030f99fa81ed839157f029b9d471ebb454adda8962ab9186054f20bf60cb70130a1dbfaa500e89413158fefee2fb1f51174bd810696a764654c61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbae0e24e5e3b8bad8cc08096b0ffa5a7f910c40edce71f0adf0959659a09e7afad38e2b6f512d3de13cc50420ebe60c7adeafa91f0fd2d8ff225aedce55392f924733124bed66c85cc98a4f3e92dc87ee828695f8f332e992bc64b8b6e388aa06b62e48ce57b3fc94f8b3d3461b6f46f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39e86f58a661786463e65f7cc1387056af18106d9e557b4536903ed3aa45d2670fdb2dd17e356da920232d81f00fb97d14059a1eb4537f7b30377c9a92eb2dd39ebc3057bfbb47cb1748d6194d19c6ef336d4bf0c08617dc693c85fc065058fa6976b40171d622ac2dc69dd43dbfefb57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h557a1c229a59157c62091c6159a5df21c58fb6400a25af8934636aae2d8ecde45f4c42e0d758480d7db3e172793ada9a294cb439de24b462241e0eca1c140657cf700a156f52086167576198b1a21d5aa305d6b0a21d1bdc28f65dac5d7b54f804082c87bbe19214de26c860e5b87e439;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85e87e52a6580d6bf162027bde94d8de0061d4b54f901f1dcebbc0b480c8c7b066d8d9d7559283074573efd5d9fbe8359bce29512c9432f39534c439a911dfbe37f83ca71b251106193dbe9322cf7ee4a0a74998379f6683e1d561bee4e2d19621bbe13ab193e7224b26e9b7225f2a3c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc242c038edd676cdce404b647183f6a70e1d2c8a61228d6c84da4bdefbc16c60a9816ee7c0632bfbb36e6f3137aa12959e5f1a8df3da60eeba343efce3db634b4068fbce61a668a65dcfcdb2399314440faf572e41c99a29e1f38a1c60c67a109b986b828fe3074936d55a99057504277;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb84214600a79f9ed796a2979e799232ecbfcca2298089eeab9c4fe782c07b35c9e7682fc3b347a701487a741b1717e4824af00a1572a49f26572de2b3fe639ae184bc420e4bb97f913369057a9cdf94de4b337a45f892a66855205d9e0961bad9f57bee89873d2e9bcf5a094de6d42e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd54e4e26f0b28833af3a545d54419f64318ef704db2003acf66685e95e40d7767741945bb32b60de41f5a6ddcd23be1defe7d8a342639ff448ada109069932a644789ebb3a95ef80658ed4bef474da61ba0c395e86a6bf96fbac2e2c187cbec6b7ee80e797fcf332b82809a4eebc7ada5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ff7de15ddcf918cdb782108055305ee9219c15c6dd80d10757dc9650b115d9e05d9593ff18e5cd9db6c587ae37f7ba7253fa3b515e270df44d66e9399b5c6c340c80e66acafa7e402b197783ec35ec4d3d2ec53ef72f1c994dca7e473ed1e884547ce32884d3813548e803e1138fe681;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h818611e29099695bdde9dbad7e9a8bb6323309801c4dedfb58e31e025196667041b4b42e2c7cb955391e81021d66ba242f8d1c183cf2c4dfcc175dc141e1f2181ace0857cc933d190a2aebd14ce2f8d729303dae291287f02ab2bf9a250f0081c07094a73d8f1e2bd6697e44fb4fd0713;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf814cd7c36496159cb2634d3f3ebd2a2e7b16c63ec72bc3e625ad0af71027a1e8959138bae9607041490fedcff567a05a9d268044084372e2b08d10ff89c99da86c707d77086424f773b9b210ce63aa2762e482ced85162c8b17bf4fbdbe31b89132c131cf6c9d9938cf300966e808efb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13ce68d1bd94f4ca5be7651681a8f7f532117dd6d892866a03caddd4f7e310cb26761b912240089a0ff24e23c1477e4dbedfc63719ef7d7b07b77810c62a4cc69a4bf72788e7e5328af93eb56409d6a088a4bae7a6fba2dd96a327c69f12aba860be50540fa503098409678a23cbc2660;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h422ca68d15ab62aba65508d49b64eb312fb5ead6d64a6b1e9a85e0b1f7fdeec90f508d061f592236254e7a3e33d20db75f38b0b935f24b3f2ee906e25d4c8eaace3f8fdca9630732f52d68f8fbf698af1f0b895d1a60682a94d94dc9ee768533be9982a8ce6fd7007690789bf8c52f554;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95483180813f54848228f9c6c62d8d830200d1822e83721e7ad2d82d838c1dd4d35c16d53c7ac91d5789dcb27d027a62614af5e19c55461384b8d40be0e6bac76a227c5d60a0288f1caa53a8d77069e0d5b0a1491423dda51b5211676bd6b1a5351e3988207ec16d708f58c73109bbb93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ae0dd9888f3d9944bd940d8a93323ace3835f62f45f2930f98d1d07972b09983ee0ae42d0b75a52179bb5a4667a57d067482c3671ef75f9311d33e7b15722119215ea3513b9bcf74b459ce0d8b5faca7a65b677a0935c3b808ae7122a973c7fe094df4940d8ec26b3b228f84435858b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8decde0969d2706a60d3d5d9cb4c4d0fabe9594416247cc685b2d130409bc65eba9c9482069b41d2cd67e41802d50128e747253750eca02f06df1dcc63f978baf9fad728e7088d7fed1cedf4833d73b121abfae8535e14dc75cefb470cc291d26c0b85244d9f8cb1e42eecbde32d4bf13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ac366003c870fd76f65200e2125551ef00eb18af1c0b9d6fd69b810a6753bfbb6e36fa9a8d51229fdf5a85f2902907f6458af299f0c5f59136d81d36946e8263759de508f80f6cf4269dd992329f5b67240069b73edc36a227fc8fbde96a01d6bdbccc1d6d16063e63a4466318807374;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31f563c15d712ee2674e1c8664b9ecc10a0f72108adb37283055dc47980ab7b36fd62ae6bcb46687f68791505d81fb76f63a3f93018d3927855ed82b5f61c78973d683f8572e7b1afb101c90a67324aed0b6442e87b94fda7682f32f70cdacadd5cf0ae522bb08d302b07b277e90bad0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b9a2d5137cbdf115856284fc7348fe29e0237f7c4de7d3e71fdfa67c84ebfb86d2acf8cdf5ef670e6f7d297584519a7ccbe5da8e5d9581b220aedd47eaaf515991abad2be2ae8d57928fedbca91135cc5c12586d754882a58dd1ab9bf6a3f7cd925829279d28b3ca383cb9def638b234;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h299fee3b08f47edf9de27d31a1093a560e465d74a17ef697e9d175ed0136e9e21c73142943356dde0011c826585f4d4f2f83bd0eeb1fea79cb801244ec8091cfe45ca4be576d17d9dcbd61eff4d855f0cbf8713b129345194bfe5afbfcb148b58ad00c43ea9de054cd05e948a288282ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a512149063a9ef0d4d1f84d6a96d962c95d4594430240e0ef2746ec377e62ae7b5a5b62155dd7ca44d710444f2b6258efd38cc911457726ff08d91322aa1cd0a385faa39fdf9a23ecaeb6c7bd498b53b7fc30cfe5a44c59381a3f192ed4736a8d67e2ef4ee33f9c50cc25024f01c8894;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he930599688ea9dab6647f0ff168fcef439bf93e4da00676749b3fc2cb507173725ddb7eae9bed2b87ffc6d12a0605d905a2699c398e1115e878dcf7822fc8d20d375f0d6dfaf33d0134f7869a24d08cb331c910550a9a7db62ae948d70007f0f8fd17d86e2959065074f6b5221ea0f8c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6476587c01de51cd010a46b9396654af1f65537a2a0538703e43ac9d1f57e0b93383efacabd64814372f25f86ac7ee8371284bf770067f44d972b58ae93d33427056d5f663ef4c23f78ad58e7992714730a30b78a211c091f0d7c24f987b63fc8ef13bce0c260ee6f894aba18349ac255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd595c4909ba09520989905c37be33c99616173f56a85fcc732a8563a23b9c0fdff7370e24a74eac1fd2f77aaaba8546797eceb2953572648882fe7671879a86c028eee79c261fad570744a32409d67dfd9c4923f10cc7d40befb5e5d606731e3179ea7767300b55a4eba0d3a3e74aaf5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58d95ad760a840f99e5e7d9de2a6abe014d611bedff3a4054bbcb3cac18112a4a2190475446e3d2dbc2c4b988e3d05cf4e7afc2273137d17cfd1f1ba4d593784d5c51b40a06cb0d5cf98b24c4138492bd9dc41cce651d7cb9ba4115ba106202c1cbf29821cee2358413c4857705160414;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8572a4786730aa5346e3ecbf4bca3e2c301900854d673b90b5e57d9756abcf4681e68e899fffb49b6e347b24449addb1a3118121f2b0a10d94c0740d91941f738b9b8869f9f4cb5cc55f4f861b969e443022d62641e76d9e159daccc8406b0f7f0aaa1ea007e0c2d48a24873321bfffba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fd82518a5a2f66b2c41167117240036e21078a32deb0539d8ec4ab13054ce584b922bb58a2c184bf9bc56a71777a40292adfd278b4b7fcc99983b673bb2d220e6f7ba9e7f4be1557777a2b675d04cf49a7401b07e810db6a0ab40b13da4bf082b923f3caf2bd85218831c490c1b5d5c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71ff02999fbea73545d2f83d3ff9f5c1dc400a53421e61d8f48fd2b91765291fd71a40877dab407019b8c1c96ca677e2f7f668cced1a0d839fba480647038805d7b3b311e98d84e49fb881aa3d109e4627e6cc399997fe790c192854d9651db0382ceaf4b129f825bc1f989186199f625;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6caf135211430802870abf33a4d9f6aba789a8e4951c203d8dbfd34bef6df04e33c7102f93ec9fac63e358ee1dfc6b9e0f22e4816148929eac9db2ccd79a4293311784d0bf60470ae098f92447dd2bdc5eeb0e151aefb7a9d769cd627991c743fdd42a153f3e567b4b3da0978aa5f665;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bb308211f5cc31949465867f3368af49bb69f615fb51e30023afd1d7657e10f8754873f43621fb9de3fa8f1fc0ef7d68dcaf1a755017abb9cb261502febdfe4794042f1e60fbcd08ad57f124fc7ae688c6fb0218929aa9bceb9c70eed282028cbe72bb0f6bc2b039e55d952b8358cd4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba83bca73a88e6e29fc7322828752f4f9d6b67a02b3be420c8535d6dd22b90bda2cf39756cde1d9554a715ddcff409c95173f109537674317cf1281091b9b3e912d925051ab499225e8dec472bac5835895259c16921aa1876693ffbdcfe2e95cc2dba386d65f8b7320ab54633b5018c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h709ee619b3642084da20bd1140aab190d96e669469d7f43987ad988523e0164435cd597d75130aea9b9c4ae0e46eed8e70552a451486f414a5ad3af401522b6077fee7c43cfc140e2cfb8f67f664f5cc60fb458af8a2f29d872c19f9fbc13ad3267b5b5ecdf102880bfe0dd849d169be6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15332321a6c878becec523dac75f03b07c24af233f94afff3af6939804ec49512733ca28260f2507a0be45d976ce69d9edd48b49338e6317a8e21077e4c0291dccc2c6accd2f4cdcc062f4a2825d78b6bb485910ca3737952548d409b33cd0ceb9bd6274b0099ea2019d05f0f2d58efda;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc94a6f05419f906c99047a0e637387801f8a5b3e11166935630995f154431231858d5cd4241935da54974e8511c11593435504686c3d6a8cd1d41a927c9dc731c024b42a7a30af459752f2f7364117e55e7a48b53eaa7f770130d7906ab2a41328b325dd4e72d91b168e52e9f4863f612;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb12a325501fd0e7085efa4529f886b6965c52f774054033ca3e59ce11caac8a92616ee8859b417e5e759f420791fbae00df1401606ea8e1aa051fd3905b46a51236a0772c29795a9c1a15667b31d92b0c1f4041881a13ba3e5e35f1eb7cfdefc7ee094685749923c8836c91004b85df13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91d473414bf038c26a0f62651b8ff19bb73e6ab2e063ea18df3fcc7889e3512a109c2056b35da7a1d32e1c3587f912e7729669b85dc635593fde7275d1dd7edd3f726ecb13c63fcf6ec7eca5503946eb85d68538aa5ce06e36b3b2f7810cc935cfd32738f56fdb7f483ec3a1f64a42f8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2d1b5dbb9f5e93343b742ccf2702e60749819dae11498f01fc7c6fb77a33804dd25a944c41af5fc6b218fba7fcfab75a6c820877cb554a038160d980c0ab6f9c5846b48ccd35b02da8bf1b6797c277116be7b1219c316c7163b004be6a49c2b5441c1f78eb16e106cdd715e3be2ad4ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5da31432ee39673f6762931205656b4a8b0df356ec0100874ce374779e06f3a8aeabb1e2e1119d36355b424d51f9b70feb1923680b1b44fafa65594d9705801cb3c112d72c70351ce2447e77687e1e76a7a38144c7849f5b3cab4bb9467b69922cc749b078532aa338bc0e3650851ff70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2ea10617b3221d303777037a52e5f7ba96c09d0e1cd221eb8e8f802e05d161f33978bde158cf4db23d8aeee07e16669896468996c922d9cc0794a8b7550a26368ece12eb52cedf55460c3ecd0d398ec374373bd8806e146f27ae38d9dd894cee46b2aa3a871dae0e0d7325550f05ef3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h131789ee87b7657192236851143871f602a4e34d9ae2ac4cd768f4e16b3c2f5d81a3b344e572eb00a235c3315c29f8ef4fbb4c0ff3030391a9cab6ca78f28545628fea90549f205d1bc18e7038c42ba37fd158bdeee401bfa7fca4c9642fd8f53c68aa2dd14d331267f0a1e626395fbfe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58567cd95fb953b62853f6c0281b78084df7048c079af1c813d5a226dd5a1fc8976b38560d795417642122ea81e504531758febb0cfa98a711fe225ef9a09244c5e3a2a2a7deaeee9afde8a0788fd768f025afe1719c931966e288e05c99e290a62614aff34a93e0d0fc230b85df5d20c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e1d1d94ee671467d28ff12fc25a1036d0158f3024fd8ab4506d1eccb9fa83695063b2417a9f473129858e67dc367131279dae9427275715d38f1a2ee89313ab190c53de91cb009097bc45fb546a130813eae3df6d1873b1bc5293a02ad4326795a5eae43612f0e633d8c7b56bef4def;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff2841f4048e771e3a57bb56aaf7fcd89ad34ffd6c85591bfc23b7917cc5bd673b60592950fe8e5e4ae6c456e889690d03bd1c423247d6b2f65c1b39d0d278a50f8d8a5674b67bbc6084b429335d5211f1cbd08abf77859f7af18edcd2366025d7dcd0ffbb9d863d0982b68d458f710ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h179b44c6169fbfc290334ce265f9db895962e41fe0836dd7ef0152fe1bd131036e697be8e4c5d472521178a6b1dc5e7a9adc58ad5c395101c700f5daaa567d5ce3f7bcd4c6fa554844bed6b39c00a6d0816b05c4cbeabecde35d5c1ec65fd292d92377ea1e01baa429daaae2a11401fa2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92b48cbf640163eeb398980013ec636fb62a7d3eeabf6f226fc91e13f8a7a80a5ad15e72d369156fad36c11693e1b06fd6b0e9138c18870418fccf2b96d7331f3d017d717e4eff423f88cdab0e1afab338ddbad574d135071f33a74469af714fd715d0856fab6d6be7a17005fe4f0435b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he63c2b43d1c7d6b78fca2b2d20a595e49a6ff8ae3543a0a10a03bb96257257c8b41c7c999a5fbd83c1b4a8ec880e89e437cdacc62ee2eaff897eec9f5bc713d3c52d4b48ea1d3ab2f228eccda8cb6362627a0c745f8a14794cc7b6620faa17f80709ba4089c9677c78f4b887cd995c3be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4db63f6324c6a1c73384c5db8d892cb7ea98922b261da6ab519e2cc49284ff4a81d7205d5ea991f0b44278168694ed93de80c8781061558f0c9e66776293df33af299da27c0c5c4d18ad57c8459ebeb13356a5081fe698cb0e3e7b35ec082bd177baea425569cdd3ac9c96449e49bee62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5858333f20563e687da93ecad913ee3dedf0857509058d2ae01b6e78f12e0bb2839d4442ff5028620f7e0e05155659e9588cc32b67b3f1c7a2468a86b9703b096cc09fa0fe694aba8b44f8983d6209d1903f3bf419297cda2564b60f9251b960257b72340141f818ca56608aca8d8acd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda08e9ad44c4954a56264dba8d6ab1b57b5659a4f53e93b28ec94aa1f27e410566371a4d28de62b4a05e0da9828f3f7b41b2b77f9ed22be11ac2775b47c65fd2e35ba238375f3e41b89b430ae476ec9e6e11296a610f58637d7dec884f309298e8fe91a7cd4a8e2cb4a534e1626c606f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h827606b74fa0aba64aa1f7d9985d253ae7a740d9980ee3d20456682b63400104347938ed1e47e76f16b993a5219b1b5e915444a932b1f5c16f5bee8add7c52085eaa06e4a6a45db2e1675f836ca3f87630b1b48dbb0f493a135b650a943eda282bfab6db8c83d0ddc46bd65910ec44535;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3be1879da2d8fd8c27833a5eae374251809e4171eb3a0e58bf7a865f0be85be46a5e2f96d55f6e105d2b6398c7c984dcf6aae8b1a4305a04b93281a6aa5ee7c729d47e34a0febdf23046b6f02d6d0173618c624d77192be647fc0f718fb9a030d882e60d153ec1d7cebfac93cb1447a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f18f5b08d32e3e0d15f8d202e92974be8067374d8a046a35b48735e34ab547a9c858a1292a2fb94d79633bb941f56979ba33f105ad71f646e44754cc1e5e111397b0affdacacb31aee74343cb4883741f9468e807fdac1553ab924312523a4700bbaf826612c14f23fb817d09e7de9dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b1015e02a5b81cacc9b0da2c3dce3ffa97d32e0620c8a9aaeda3f4938ae5cdaed2609fd45c331b65fb0e01305277719fd8c6de49f0e20d2e507aaea44807c8b01260ce1debaa94baa8a11543790692954a9a528152288fb4ad98e92aa135ebd41212fb8eed8a254a22ce1e38133145d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ff59439e4ac7fa67e50cc1374bdde3029cced4b397f807626dc2b29335917eeb7e0d296630516831e3543d671a03e5c0a467fd0bea24e40c77f848043598a9ef0d7dd26faa6350ade0e71348a01db7f17c33696818a7a482d4981991b2f263c2e5e4a014d2468597c162697b99351e68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e96e9a6c9ce5b642f1e642ba0cb0f316c397f4feabb35933a6fa4a10956d319686278c3cbc22750d64b91f7f5e0b1e3c51ef4b4ed88909ba7a75b0881c23079b84e1b96d426c3dc8bc643303ddfaf388ea0e89bb32ebc10ddad8632977ce317b57225d42ecfc9b5d0a0e9e1dccf877d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b22e5cd66747b2c42d840e593bcc0321f29749a15cc980ddb73ccccc4ce92b18c5de50a303feede9b8d968970c341e9d64a11fc98d37c3cae15c9e8350c423ffc9568852472719a67b220be663e00fab00ee7a030d5c265257f9e4364fbee128963e81652e5b7818985405ed07aac4dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25507401a336b1d1038afbba9b9ee72586cf7011038a9f2dddddde477bb0cdcd7c3bd96eaf844c4e81a160f597abb4b4f0e177e7df5ef21de77c76e349dcb6001fa2464bd6d97a592dd773e1b964f2ff382a6ae54f63967a0f437755f932cfccce6ae7c341b318568acae9e0b67bda193;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26625a38d85d54ee17f411c9a480a6281071a0c7e7ea7de05a943a53ac7981d80a84a8aaf4ed46532696629c8b17c6ab4ba4ef8a5c8424dad60172b10adc804adb667d0664c184d56575ba2fd54b45c721b904804342f06967ad3e969f5a504739e5ab189f0c2eb5eed9e6efc04aa9d97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c2b165a21fe1e5c3a40a16695b4d160cebbf3386b41bdefb1f2321638de82c1643fb92f304f30da9de4c8a6c8ef3e674bd4bda83df6bbadb9241c0593ea652555628015318153b40efb062338b7c8e5a69332065631abfa6ed9cff62bd37f8fffd6967f60cc46795ded14a3c14bd7d72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb0d7a2204ee2df771eae1a41fd844d8974f3dd09eea1dfe24014d4e1cf0122344e52c9762212a626ccd18cd13378de6d44b57287d4b0f65120be2e56d47b0b3f07c76f071b4acd77a43cee00b823495c81ec40e950d2700b9dd6c19b6c9e3fa4025cc73d0f0c5f6f306a48b06821378b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10f2e897c75499c056f0169589c55e73f8d61ccba7ff0c526cab5ac85838fb661eb5c8edd013fdb5534d1d3564fa7c87ecb4cd4f0efeaa8c99a181f615a0b26d554a6e78be17d1b94776eace9384b85d7e40785389c01e511d2959be4d39f90bd2967a278c1f6dfb64730e11144cb9624;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd5c21a8d62e9b05cd64bd035f56db4ad29e5f42393af44141c597c4c4c354bf7a0e96d232b174c79f14c82ca420ce97d2cecd081b830aea9fc641b900218d5c2047c3783abe8fe3d6fd7571aa7dba814ab599da8661719dc7bbe4aa5670f3adc738fb94cffd55e7c4100f17e9bba39ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34b150aa24a598f3ae7469ef6f99d5f5e2dfdb9cbc5590e64bcea8265a922e2abd9d7bb4f2636ab27f3e915370855a2064b8a2793d5a39e89305acc40ccf420ef91659bf91d3994fe15ac7a58c467350cab19d5ee070a5c66e6943da993597642a6c08d160aa1a0da28fc25bf755a0629;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had7752435b4402172d671bceaed7448b1b006a92d4a243b19e0a03f8a2363ba32f5a01635b9f8b98f1798720022a7b41bc3f84e8f03b404686075a5b90b67729f069cce92d3626688018ee3a329ff2a5858ca122bc58dcff054c4cefd9b4915d26e6a0b0db4d1ff54a1b84bdf3fc59b70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1002c09086dc97e89b2b46e1483fb5babad1fed9968c17984ea1c9a419866751b1b3280702ed7989b453ab7092f47c6db9ef0c3a55d523b6370d2c9c06c5a63185cdd907e4d53a761c04c2d077bc962e3de5065b6247b5123afdaa2c247dbbdd77c12ca38ad80d6dd371731c3e6b1c5a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74283e2d19e7daa95349b2e13e232c653961946f9245022a29149a78e1cc6a9be3976ade7ef6c583448d10127613538183107f7e13f30f256fe02c1a9c6e4c0537fdeda67b94c55be1aac0a6a36803674774e497f8b0c586b600f1f2242e62a60ad671c4799daa707b1261b254eec8c87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae65cf52d6331c17fb3488e92e909284c4cd48d14b85eceff545dadbff996e90389fd0254873c67743888c95c73a7c6a8260416089d53e1d8b7fb515bda3b45df7e357d6a10c04ab86bdd8a861b2388a247acd55c0e7b4262bb8d4e10de7cc593f52745302ffc141e545ef8206ef9800;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ae16862a0a072329157889f084e0ab74a6856c8a19bf9848cfef2093ed8b801d9dd7991aedb30396619e6358febbbfb56d0efd7dd40bb77fb32f6c96332703181804f6ca6ffdf41b2a71b6b4ff040ece219528d3de0226d2cd739d95e818133d97024eb51fb77cee74b2ef1eea6574c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd1635401897e641b569398aabe6061b539bfde8b5a412642341e2afab149726ddec44177eece1baab9c404aaef44c648fa20e25f3e7b4305636f40b0ff4f5ca00744e6af26c475227a8a3ddefb7ddd09e812de60dff66a8d979c3c317073bd5bfdbb778b95fd95142df696f117df1c95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54533dc6756e2f6d01cb56ff3b2d29f1a46fb65a77df73b1b5d28cb960d9f9ab20530ed332978b583ed0060812bad9447a629b53a187c0445628d713d37914767c60eb8c505683f8ae4fb9629b77a804666a7c099f566a86840db24a4356f518448551ee057d75973c11533924cf9c209;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bfaac41717b8bcb2bc497d59aaaea77cc17068b0712d7a98a3c057a6d62806beaf4a72ed3b32ab1e14c6079e806884e33e43cc315169e4a2d2bdbe8978923a341a9f5155c1a2bdbdbb4d077484d61246e4c42a7eaa4a61391e6e5cc5ded0bbcdb8536a11342ddf15f873f46496a22e95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f3a0c986fe9f79a89ebf09b9895d2d7ef511f412e72b2b86c4b50c04c03e190eb3b370077052d5383266e7b86de0b6056aec039b6cd1bc8b4aaac9df68471bb445ebe9b5865308693f182e728412ecf6a0823fb1290c72308b84308155ec63b06c4c47b1b7681e20b974d700077e8401;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1d2cfb97acee4f3d085144f56d939007ad1607a8858d2ad1ff5e100866a47141d863734841c2d1aba335a47f82db023d9b3590c1d37636f34ad24a8605bec6b6c522c22e4fa1ea137c641ef2f0156e1c7fcd9ecaa696e702fd1806963da64d438970aad08cd5a743f950bba40f08867e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94a70e708eca704bb5a3bb969d8440bcffde3a19228facf74909722df110dd56a5da639be30d6f779ab92e2b079a2720d3f362783b0050be057a8cf108a50fa1d1c68a6069fd667f4ad8e86adaa9a100ad317beb412398bec6011e49331326406adb42fa358f452c802925f5db881ec3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha13f4ecfa9af3ebbe73c1e3e597c84c016d4c3b6eff6dade01d6190f8421dabe15ea8c637e02f89cd0481bc5777ea1a0de0566d1a8e136ebf99c853cef754c45624074bbdced8ba03fc69856e11aa2bc97971f2136f9a4a3e18b2cbec78eddd3c7fab39f54e0c9985867adcc6cc0de8dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0834baa7e6af0e1d7b817a2a403a64d3bb95f7248ceb16bd962faf95035eb8c027f00515a677092a2c97f500e1b74669d5aecf8ac03e95047e0010b9b5ec36aea88299ec38bb8e35aa4acddbf000ece3f76b4cb73d5c4980d23afc86e3df79ad8a7d2d9cf7b8bd45a289a20855e9d12b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha67532a6073cb85ce2fd7798392e9d0a1447992b0588d98f05c25caf45af2d8777b592c17f7a4d4a5859a3a394c7e957307c602d474c4aa7dd7aa791217271a7a17c0499435fff6ef4cec8f8f1e938ee0383b29434aded89efefebadc91f24a2b5d3db54f05d28f36895d21d17277842d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffb89edbc9c4c05b93c84318780d73504917cf61dbe74d5145442e8edcedb32883930fd8589eed9504b3a8b832470c6754af6b28c8471374105f984f610b1de6f066c87b2cb5b5ba1c1c1eb12c0e465b9c5567a42416ba1e88341ed7b2bef726c40ad8e5c47095262ac4d4b6c48ed98a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haeb8222fe64f7388a0ac3adc107c7cf20be5415427d839f8df7f5f3a9b96dc41a38c0595a4d913a75ab8cb39eef389096fa0fc75388f1f13f5c44c7d5d6b958bf4614573897afb361039debd10a08f490cccac7fbadd159b56417e2c24fe96d8723402506567bb3f984761142e4662fda;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aa975ccdf40200a42bd497f022f7ede39f1400e03b09cdae4708d3df59547c3beae629a8ddd5bc7f5251a05d76865d3aa246da4e1fba5a83a09a837325a2dcf2635ede8ce7e917464267442ee1218586d1dd064d3755363d71d2ac77324974c145d4003a749140071e4166ebf7197d7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b0ef190f1d16e626f1d60e094bc5029e3c7d4f0a58e109ebcbf5258f6a4c036a57964008696a22b4863d60eab1eb4e5ba61ca831cbbfc9453c1c6b9aac3d5f40ce23453a58b0e21ed76c278beabd6ba9eea235fa0bc97898434af28a403293089bd0f7fe6289be137c2b5342ad34d2b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h992762c0802544bbe0475625692d8a2ee6194765a1e357aeaacc472e16b14d8a1e3278e3777958807e5233ae73b9e2c3c49e20105d30e0b772e6a02bcfbff29d71d6650fc373a75f13c41ec44b4b563a5c11c03ac628705721570df355162b4917cbbe3922be756d96f148f52661d0018;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6ef794f8140fd45567ced25659a94c4ce03f0870c1505c4594e757156b1c873bae3ddfe1db0def0a21d21880b9c089105a56a05cc584151f65970e5a11844d5fe5eaa506b52246728cbdb820a29643cfd840442397e9898ae4f843180f92c345f4fb73d063c8f7160efaa323e2fcf465;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f96fcfc808c2932d6e4b77e9922da803654e136b340afbd6a875d91c07d7e1bffed1aecf3b95738ca61d00c22d98213aa45973b2ddb0ad0a218307bfa219bb04465b314e5540ef149f3da7cb6e42d9abdfe74d8c3856b7e103a836df05aeacd83aba9eb4d365f05025b406443bd09bbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7853b720e3868ff47e91c3e22f3c97d1ae5532b1efe5519aa0e3f805585384ff4eb029aea037eabcbc575f92b6da1c80dab9c4c49517192c7638e52d1cfac39e0d6dab15d8293cf6b1284427a43abae089c85ba37d46b0187a8c0d2766b562b64cb1782a7af66cf52fbd30052c4f90960;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h837ad05a4caa73c449a029272cb23bd00bd9c456d5fa7fc3f96a275742a20c66484e6b021077caaf27c0f20f849b01d5b6aea2a2698301712ab8bc40dc75fe613ec5271d06a3948dd016693100702e021a36fdaa5213339ac2d4bf0ba273de8bc49e7995735b2b2e91d07effbec9fa24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1067703c518569a6bd05248da163371e5ca32ef851ac3af93d3e7cae56a37084d199c866e46d790d9a6d0995461dd87925526ccf0cc286291e9f02901c693bb6e4eb6bc18135371157614d8ea0ebca5fc53b3da56948f84e733084a651970ed7f7d573f8f49fd85e946a9ef81cb297b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7dad7bb729c8588083d98a2306e2ef5005a6a3d25cbb37f9615040e7f4c180b06a345347f31bd87b8e84ff55a25aa0ab11565ac4197added03741cf9ff23fb9f3d438f36e0440e6bed2345d23b158ff732e913284805eb1703977c37070eb2103a95f507693db9ea7e5223531d7604b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5c5f354878501f00130796e601b2f1fe0c2c6682122ee27e0ff41f3676e498f3a9e957a8f8ee5060b28f3c10febb3f7e2ea80b21b293f0f55a411ddb21c53673d2d14312f518afb4ab7bfa2a6509d6a17314afd1d95112b26bab1aea30e04a7489188938b10c1958abc1aa25dbd3a0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2dc6b81ab58dda34f7fcf94efda2424bea95942eebca00c5617b15328a74ba2552760679cd49497d82ad856e550a96db955281de778034bd067a2063a9a14201635c349508878132c49eebc3a93a5195a6807d37cf305a7d31c02fa2cf0563d69a6538b6d378a90ca26717dbcedb06c9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h777503cc03d390d71424d8dac2ad6c8588a49b1a2c27f3a1756931b608277ca4b0e822e853716523eb2d2200ad3a2f235ee7a083ad559b7fc059bb590a3fea7e42fd190f23f7d8b927d7fbfdd8c3a31dff0b1de39bcd3a891f60187030f37c8a9b91d88ea4b75c6aee6ccefd94e398266;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha67a95c1861d89d6bf0754672689bab5e9b01a6a56a9114d2638503c47dbb721a27d4a325a66ad45fae12cc93f5b4d7535fa650615cd5364bf3ccda41186500636764fd09f6516bfbb4fac4c7def5183dde64ae43ccd1d6d409712268931c109bd7cfbcda7b455452a46a3367012a5a54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h878bb8415b856d25f205b7885959ef7f1e8cc31663464815945ff962c7e8531e2c3462271b035e1394599d3d63f790a2d3ebb4812dd42a93c7274206a3229fc771c439ff8b7f4819acfcdfaf7e218940da9088129034ae9fb94a24d21709f2a4ee27b1801cd5c0af1e6ca532ccf4f98d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2b189679f5ed8b17b3d29a6a66a656ef8267a721db39ce85bc7b24354ca5b336355f5268688c6978617873961e5680fe5ab88666bf482dd25cc0977cca9ff3b040605234530bad310946503d8ed7c1451835ae5aba6a7f00804d53d459c30bdfe4d7f849494e1b2e7388bd9281811ff7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3586ad5cb99beb6bdd8c4659f38ac85333d1f47fe805536373cc3cd7a46b90d7f14bb5d51dc8f315fc56428488c683cdb064f2073674572854795f1f5b3866585eaed3db9805969504b4d928a17c69387d897e01ea9f99d97534987ef464fcc9598070781d399314b7a43268fa19830bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cca12f5a67d6db7405e4752c44c22109fb732cdbdda21b2c1c9984e6b0d6a5f86828a3423449438e1cd16cb32cc0be1bf8a9eec1d3126a5fd8aa0d8ba57b2ff9f93caafa801a45a3caefd7cc9dcf31a8b857d13deabf379ebaf40ce08efa59eb1eb83405663bbe9faf37106093be26a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd80a23a94036ea4caadf2fc151b813b89829e6b6a91a10a037e70ae54f744b71923a463367c6bfda1160acd03c2e88f681e5da84d4e326ef33cd57ef1e2a186b60cb91f3252f3ccc4004925ee5d4dea2e9dc949503f5caf93c38ef0c71013a06cbb93bfb8700d144608400754e295918;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97b131771e745903d1e42ebd2c85a0ff46b7d3db5b8eda71e339501ec0df0d2b8d64509ade7f91ed19ea9420dc71a590ed16f8f5e2e45def81fafd41a1d421c10eabd769b880f836df395a623b38081e50c93067fd5837d493437c04899e68002ad89f12a7c220693104c9eba13694fb8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f8d5f459a86c16f6da35bf883881595123e585d917c3b1e6528e4c18167cb6b232d6cd300a3f32e1de3ac6d17d559d03bfa18e664b053b2a8c62922a78e2d950037ab7050aeb070a7a344837a440b681b25b5808b5d88a915f3fa261ff5580fc0286db986361ccb7cd9e19bcf736e397;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83bcd98450080a84b5fc013272cf8facef192b7645410145e3f3ccc4d439b3b681a1f3e76bccc54cf992dd019764748a8375f22e64abbce5be95f4f02853bfe951878069eb2f028fbdd42c3238f2104e11b84d8ac07eacea094da4ceb8e983b107c87faafaba0f90c6b2a407b3b792172;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d4de50daec4af999548ad8317cea2ce499666d1bbca2fc1081ee8bd40fac9dcac6b13210a1ce62a4b9ced015618242161f96239d5853cc5ed7227656abc6a5411e620ae25d633bdc4060edd8c5e6699cc6f644d514e2d0e1eab56b993d4c33fc8bfd3a83fa1bed8a39ff1addf08d102e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c668f359cb3d585950c3b938c7a02c09c6524eb7b33acae4f406898b190d1f54c5c6012b9b6236b3f813a6402e7d55aa194c41315dca5c53bc9f282d76a813961ff28d4adc0a1d70d401a1de37faa6c5e3760cb9c8417a42248bee8f8e902a1a1f5e84532334020ea79abc90b809af1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h459aecdfaff5c403a1708c784c7e69cb618ea092c020d5d6b5f2168765450a80bf20466cea73aaf9cd29562f6b99520eb53bb618c8db8a1bce8596d509a308b0260ffc3caaa50ee601800defff1686567b669685776930e07c2fe7ae900d11cc1f030f6d78d518e568968a891e24fb500;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecf985eea6a440499741bca3a11280afc7e919bb89a75afc15f3110e215cb6ae621ae5c9de492c837aa225cbadccfd9387677670f671f5e1f0e0a704990d51edcd1e98c2715653a14205bddc1be4c43a0d59736c0b3b190e59ca592cad360a4e32ca24b6838988c5280f10cfc3b4a1ecb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h308c3b5d43087be8b120923da59ca552b2f24fcae78f4961afea4e2abc30a7712cccf0abcf83f9c0f430ea7fcd538e3450daa1ba27c56cbe31115019765cb7a239045a247c295be744beb89ff63620582cfd969abb0cb4a14e844803da807af70fcb55cdc8c5ecd37eea7ecac3c2513bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ba40b18c2bcea59f487ab72fc385b12b841a485799febad802095ae43b18d3cf47debcf69feb15f2618f51d6ee4dfd68e871393d8f91fa01352a9d1ae9496fe1d0fc947eb33aaf18e5b75f1f39c8805259c637b8f9ac1ee02910738061e7da04558a78208b827231464bb48ef7cfa09f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fc108d64b9faa164d3afef25dab5bd23656281d69a5c1f93690d661d06c3cd3838feba3069297d7732a7508809965dba190c0f23e2e88fb9d58cf950ed195e090d0cd9b22c7d2f83154b505ca843c36cfea4ab7cd1828f75f91af9066483cf78851c65124435dde7d23a8704b2f9903a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he75ddac01da5bbd940fd26ab6d0a6bfc3b3ca00fbda8435de19cdf5176eb087a02e4afc5b675c43ed27f560d75dd0a6357462c6037ab5e27b1ccde27bc970261a0b244127838e5ff3238629119ddf6826d946bf2cf316f4f7665e0d7cdaa8d24b1c7325f40854e6d59601289d5513bf2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h187a2f4d1852a88aa8d003c1b184ef5b2523babc87b6b4414f94e037fcc50687cf798a4b2669ef2466e1cbab66f5181be5aef3c3bc14099971f66c110d59ba3297326af99477c996e112acf16353d427a2b1dbfd1a8f1c5b90b3815259da66e623f11d523dbb81cc922d05b27b05e5a2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74dfa589fd052e0a2952f2ce5a9c33e471d08f1414b9d96a3e727053682a0a20f96e14bc8a207131fc675a3dc95717ebe75bf23b2591f56c81db4f3272e3b1e4f9cc68d20a00223124a129a4cec2df6e69cdac6e49ae40624a877172cf1e3af4ab51d5423014a13610130b288fba9e066;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8e26978d7669e36ef0ad38451e87d86d4fb4de92fb31c3771a092cdc6610ae263568ecf27f716d33925b5e74aa85f174fcda14723a34e2773decd6dc8fd57389c0ccc8eb37c365fe148e17092333126017329867c4393c08dc2c465c5ddb7ab1960c3f7af861b3076d9c047dc0e6b0bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f66d93358d397c6c69d54c81b8eeac11b988652ab4c2e29c6fe6341a9678998c7a79677870ac32254c3db4b0df8e445fc5e423929e8f0e65538aeca882ead36a7aea6b393e3a43314e2689f7cd9fcb5187cb2c71fac595c6685e40f049f080bf3d6ed98bc294fa4fa4c6a1b551c865b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ab6f083042411f8e2fdf4c7e440a67e0c056911d46bbdda64caff3971dba62330820cc42982ea3e0238e7f30ba15cb905f3d13cb96eea58e6e9f69417796b7d64ac874cba4d4469c19058074397070b2d8daab84d7b3118ea1a75848719096faec290725d176bb4a2dac3ecaaa5fb8be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34c936c788bc1c3bddfcac310aa057ec83e5dc51d5d2b7e48278e724f8aacd189e0f898ef0e52033c684b7ad8747d792de1a661d27cf081d461480839b67272234b78902e27c991c5aab7f813f01d91ebe0e80cf9cec6517231aa223be7374536b24c1cbeb50bbeae56e0a1c50f26abed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc16fd55a5f04f2ea70e01d867b45bf8b19ce815df65b33f91f045cc39d52a252121e912e16102c7d038452dccbe4daaba8f5425eab26548b3ad8443c93177f043c42ea780d29a526f6c816ac7cb6579bdb8a054c14f24576d3ef57349cdc806e16f8a602cd9b6b3893df13af2e768a3bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94e4e28a80387c88ea1b6f76a69ec60ed182df59207e0faec04b56a34d613216fed2ca96537ea1cfb58b158ff577c03a9820fd5e6312c7a5516f0bcf536abd5ba9481da69d0dad8deff5586c3218006fd9b4bce3437730e4c4075fab25b02d9edd484fe8da0d75688855ab2dc424b5da1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h881cebc7a79c6c2b550c138c50fcbc578ac490c31e241136cf2e3418b493f69bc75e821bd61b621a6cd61ccf03dbea6beabb6ce273b01e1b9b90c66170572ffb59820a9c46497c56ce4fed45df5c00e51d5f5453c24c5efc6ae79b2706183ca27a9f8953b95474b25228895ab6bea5129;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b421d1752b1a3d6583641807bfbe3458a8baa757069b51c2a278f784eb16032a36b300ca5aa3664a2d5cbd47a80fde209db809f15f507432ac66e194761dfb08f3954c5405f08ff0868eac2299776699f3c792a3e7ac328e134e5b61caa0d3117891ed854a1a9955ed663f48b245ff8f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a60a2fe6f7a1210efc325f6bace2746ca3c6efce379929ace9cad9dbbc35d5544752a0caa91ae17e8b3247b09d8585bdf0a5baba5e9cc190dc3928a774f3ce85bbcb00daf9a88d9ba8cdf007fa549f4895d21ef7997c0109525f4b3e01916aaf971b5d8c0c9d2c2c300ac0c9e5737327;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dff0a1bceca887680edfba62ae96cb99256f45a0c0e535f9ab1cc19f536e5dfc49fd7d110bc1f88a733a77178ea2d80627f4950282692062c8b4a49ebf28ca480305cc63577330125e3d41ffeae82a8a57ae5eaceb9ede04d3cf5a9ae970d30cee08f8a47bce9de36bea707030afc055;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h418daa6c4b1daa88bc7961c4483295f91093875dae22e046921c050a97f86b54e6d895b87a60fbd66743966fc235183f44276a833098624b40ac27875c75009ddb8430404fbb73486c81a04af980713189b7f76b861e8a647ab58d9f045d79a594554924fa41a7145a144b16368b3d3d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca2b18ccafa77c18eb63a814a1c530aede5912bfe2f0516d003e6a8c8f97480729caf15e7f9ae87151d56f4c5bf5a4add77f6684fa9ca9bb01029f350b5f5f21829ce342cff9bfe09057570c72dfb56c234640bd0c7c2838eb0ac174126fc3dddcb5c73c9ee23e7b3b9c304e74797ceca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a201c5ca4190d079a27c08ac784e7bf7d1cf538db184a2e85a3c9ea8f10a90c269607079504767a1724efbceac6fe46bc02acf4e9281f0faf860cf8b9489c2a106edb0f177c994256a495e56f541983ac4a9ddda3337effda8a5dfc7731149fc82fb9de82c0377ca64b97f2d0130cd9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f15a992bb800950f89c83e032e7e0ad4c14cb4585eb91afd5f789af70f91004ddee9af2a795f840911e683d4a2bed2a2e57fb7395b22d77595cff7f67f59ec402242562af627396667e6ee5e60981820f855bcb35837c4ac7d06033a32be98f2b7b711f4712b828f5c4d7551b2f2d8ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63679074330716952941e5e9f841a4e2c6d6ff767feb3b15e282a7f4a09d14651c403e1d7924f4b238453f783481da7580a016253c33017da3dd2b7e7ff76810af0d1604e73d332e8a4ea5822b3e0d1442ab9f654d915ee70bb5c2f9aaf6ca4f07ca988f93b0abdd2f11970835a683c57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4cb46c5e98ad42f5bd3f33b2b85a9229cd005b96b089bffe08269618800f0a45eaa55afed59404e36a6a15a4be4af7b372f804cc9469ae714bcdebf07e5daf713d0be925d61b076a9c149334ce4337f51b72e0b0297971d36d23dd0a7668cf6f6727b32c793ac1d3635e8a966dcb69b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h267e88c0f96940409d94f93c2caefe28802d801ebf04a762a2ce5c9a406bd03f42674288895663d0aa874f29ba379010cae85731d685d8cd92217694c1f83ceee7324b339ab187b0a70fe9b81d0ecd92d0f9a2041eae6c2c40a5c5e33a732b96c728e26957b64bf99827af35001aae282;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb73b13036afd7f5d7f563916584b23b52feaaa955991c3689e583aeef886bb8531a0af0cbe09e4c4f537e7413da27db13dc302e03748db21cea888eedaeee558e9489514a27f4f27794694fbf0a4ed902e336e07b962860765f11308f54ef70a620e745055d4057267cdfd2e3302e533c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc421740eb331c85ed3188174c578706980760d0c61e57dbfbabfe8029b259c220bcc56bfb893c1eb3fa58aa9b38cd1a9fa00e3e3e7df9b645032bb97328b222a3c5c8517a0e231de044dd1e5e33b1799f79ba400e80c06fb7a867332ad1d951979c46d9d6d24b109fd10cde52162c6a14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfee7b806f38275414f6b7e16268618d20b13c478b1fda9321311acc8811f9fb80776681ab3f16005459f2f33c9ebd07f4cb33e2e339ddf86b3713fefead9249106cc51b5c373cc0844c7e12e1db308e8ca5f41365f8e773b4fbb2805d69fff5b0716e876e00f5d3b54b5174f41f603676;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f2f7988c3f20e8c8307acfd9f4bcabb0cda4efb3539e1e0099fef1f18f67670ee4731384c39bf69480e4fa1aec1e0a8cbc2936a861fc212fc47fe47bd666fbef994eebe32ceda185cf41192430e7913a8d74747f757f23f6d2d58b00374f94c03f9c39f579177e3187a770555dee2e00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ef113fb766193999c956196db11ded019763a8ccb1c5cffdff752b7974777eee3b5d6f10b44b86eca73a9a9a79ec538fe61ff8e87fce0708c42aa0d07c9a69174b7bb6e835536f5f1b6913d47b9d98ac76ca7ae5749502f6084c9598f78b55055c83d34c3ebf2eca91d8ccaaaab52445;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4daa498816e313bd3d748f72c7a8d65d959a10a4bdfef345825454321660d9429c1dbeb354ec2cf3e09a95cd4d40d5c36fd5d506e706e7c9bb1243c2b10f75abc36006c0fb280df70dfea0cadac217cbab28e504fe1da1add7290eb4a80861bca0a0efcea5b2c6537b4e18e5d91373127;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dee9ae5075ca7a8f496ca5daaeb2d1b74583098bc5591bc511d31a9f19bd413c1f270b1513a3b3acd98dbcf4228c3d4e1a2b7a1db4421380524e6be2a77aa128bbdb86e049d7dcb17e45721ddc774f8b44f8ccd989193f190c8c509c494c9ee1e2ff81552d01a455f0b721d71fb4b962;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5347403d5e9fb643b4323303741a7643a9fbbc9f591413b5d96afe9624d5c31d8048d3a97a1e39b427885022e4fc26f0a3963ffede46e4a4cf3f10c138d7ce0d709ec1d46c75e6abf6406e995e28482f4bcdf68f2216c160124410da9a4cfb84ec1268976b487b6b0c14a76e677575bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29044240e0ace1fa2568b8287996126728d1b7ac663bc20c02c34084b7ab7c953fed86fad004e84a73adce040d933bad804a11fd8f805202bd70cd635c9898fa3482ca68ad7bd2d7a65ae51180723bf474977d952ec9ffcd78fede098e5882ea217eca02997bd88e482e9bf8fb1da68a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h983eec46785c22c2b6a0ebc1dc87d7bb540fbd9d864c664fc347734cc52149442868544f8fb08af4c5ec5a28efde407d10759f7ddcb663d0c26f3acc0826f92477e5e5a7bf0716cd2c4f1dd0a9a75fd856b7393bb19e7b934e65c602947ae83a3cf772acb0dbc92ce0c36398da074f8d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he301586e7a778d5595287fc96221f8b1c49195c880033a366b065de9cffa41a0d83ec98335480d73413c06c8e4859294ab0d78439e970d11cb04d1dfc30a632de73ffbff380f0c1237ef9903fbf22b065992e8fe4b1b5128633074afb3d1493f2718e122705c586657e282a2015c05f51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cfe24b248f255e86d49e47b265d06da61816d0337bf627e58b927a742c6356b87ea1241726bb5bfdf4bc8b7cd2a002085bde036ebce0435d9c9198731cbfcf3b4c1a9b0bcd91c00d754f9724f7af87c8b9ad9c7d1b92cafce4b8e572aaa6cab852c97160f33076a1169404756c46b05f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48b6c70d3dbecd38c874fa8ae3d0d6fad3f0a70ff6919aca5120a560553f53474e8efcabc8bf630d0b3ed46250452a10f5b72022fe0703779a3459c99e5ee414cf95814f98b43f1d7ae59163e4110b71aed5a01f7f1ae802f8fd6cdc13637fd893482ea94e12ed17b5b03a926a8777232;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab0c8e9093f9897ca9229ca6f21db770c2a8417e8af24e518958001bd3ad04d5e820778ae23539c80ac56f1825e827b200d662e8b7802cbe60a78add94ce67b6a8e28226a6e0781633b935626207489aee6130f9991712ef99dbb54ce8b3e0697c4a650038ff58044421ead5f165e0bcb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d4409b6ef22f1258efbfcdfd687186be113b6be3cc292c09c96277e34f744af45f0600b418d3f1114379232eaa1569ed38453ff01e91c52e4dc036c9df13a7d7ccb7f7ff67b6e12c4daa4703a712fd9caf143c0a90599778aadf954f0f95483b9f6be0822e0dd8034ced3c330177cd9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1031375a7e9f9df1320e578ee6f95680a54b9db597ef6874fbd9cd496111520ae04815585062fdf39d696d1bb434173e213ed89ede7b753102af9805947dc2f34efe89ef13f2e5ee39f4bb3eb8dfcc317d780a53fcf8977ed83ba7cfa4266d16f8a84187ae1af941c43325535a0d2d657;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee21d7e9d885f63be3260536493f3ac45c4bb319f9841ed1cfd55fc409269c0090d69e7186024236d71a43f4054411f27cc744381388d468f4325b10b8c5c28f5779d060b6c53c12eafc77d59a7f9dc4a8e2cca35f95b834c8446f036be75a15b6a683766af4c04b016c1fa4277ab9d1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8434088818a2c76a5e3f425dc2d128d17cb257a60d425e2083ac1df907a24c8a912024e46b7815e142a8361687c3ec5ab5f8675c388a1693b9cbd86585042b1cdb63ae840ff69dd6a445be5cb0e1842052caa42681329ef736cd477f02530ff52b36788237ccd1eb5e656224ec34f199;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb23581e812886e981d97f680490d983a369ba1f829ffb4acd1f738c01481159e0553c4eb44c4e360a128418a9310008bd0285f25b0da26caf13a527b210fe3aae4b8b7cea42b73cbf31a1cff36e80b71a2392d075cac63505f5531219b21f6c40a0f5da64ae18f77f584f00895644f021;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88acedb2c92474fb1768d526108e98cb0e528d1e2e4de479a563ea1ec87b91b88c10bdadc60da78e8145cbb8cd9307bf81bc155883e06b9c670f2ca1517594e4049a259dea2c525f6d4f7106657c6fa8da8a31aeacfedb449fdedb0d89593053b8edecbfb64f6a65c4e39e79ff5a09643;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb11cc98cf8f3882ac968d3ce93765d388f5200579f5034c66b62e02e80fe50062ff10239a967eb5dd88e133c199312c56c8b51c2a98b5b001f6701ac09b36f87ff4b6a09dca5ef6fb1c0c1ddfd0a9a6116d60c6ce7292fef863e2bdf324f584fb6a95b762706b736a9a8f81552abfaee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he680a14f8c36b3ed8ba4e24ab269e8e9f20393cd2f882ba0b3f9aa1e174fbe83e543d6681cfb008763c0c9692f8da62cd27f2875831cd2cfb57ea8e74a5d6938dc489ca02060148f507ae6bb2847811dc24264fdbed8a93b0c9a2c140dbcea1122ba15525b73216dbaa42b28b93f51740;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8f79bb206eacede43afbbdb554d27bbb2464e512cd783fd7885b62fd348ed7e352cdacef6aa941a625e6681bb9f96ed0c7abfd19cce0f547ad7536cf082350d8bd17ef6e95c08e3c0c353668d9b5f5fe7bded9d4e57a1cdb6b9e1f5433baebd6075aceccdc038c60db23956f19247845;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h437cbfad3a45952e5fefed73912e027d06a0ba8ba2ae2d11c8eb817a433f67de727d67e676dc1880e3d59c7fd65670e8fd4d89b2f7f6ac5103cfab98e96d1950a21f27c5ad32e932314266137eb9d9f9b6c7b8023ac1c720a63eaa791997b0919e8b5611419670c874f49185494b0852f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32b356037e3ba4cc78ead40c0028dea11bbfae36829089e02564944022f0ba51b88dbf3f045dea4a72d3f56054552951eea33a35284841135b84571142f6d490d13ab46255946299e1e76ed6417f0810bb59da540c45e5222bd80676a03c6096086acee815ead72cf5230e7f3e42f7558;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdae210edfcdb4d642e6d9956f69f30295d0760a8a3824d7f9d7ece37b2f647102180d86cddcc8fecb8edda1a90d3d6818a5e40c8df463cd837af7f28fdeb93e627b8d11d788cfcf695ac14a967f8368e154fe3204182a22ece682dc0497e46bae7a17f79bdbdc3ae2f434e996ed7c11ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc68ffcbdf59910b8517430608eb4b3718275bf8e6a96920341b8ad3a9ac26739301b4109034996c8292b889857f1ffc203952b00b2bf258768d530405e54cd12b39869bc46007f0a5eec26583e8470a81f0d6791bd8ddeb832469aa576f7e2565d73dac735a4380d3c3bc29a11e416c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ac236b349a1ece71461f847d99cacb83d8c8c5858744d47a8be7c8b6b941f3e118c0adffa81390b7b0a387c2549ebb5a53d50dda4920c64304005b27bd6ca515f9a2fd7557a00a96ba0f9c52ed38c0842618ec626328c9821255b0573edd5159daeb7db48fa99a5c365e86bd4521f7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cf90b6c7544e47fa25d813396628ec014a724ac546407121c13b4788b3fc887ad46e352c0349bb0eb91c9a84a7b55cc256a972ed4706e16f6f72dbfbfe126555d5ca732742414f114ccbe837485c86f1329e24953df9ee6d714d6b4761916d3411726da8f35852b00b5003ecf6578244;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b3dfd6e5bec7408966d54842c988e9d5ecc1efdc639717f74a7453de778bba048b4913b924f4e2b1da263c8d1bb009e55e45b36cc869f1f1ad2dcd98e8382a89ae9f7f6d7d3a2ac24484b05acf33e75bf916019b1ccd6a9a3bf4528c0b6163ac7a03ccc17d82857f22cbc019e294a3fd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6970ae915feace5ae47e72644f9be2af7924845f97768fd1319117f885c12de93c4e75b18ed1cfe6f6ffa059919604c5c3779308c127be413c8dfda3823c386935d603f75e5d4609c9c7a2d8cc3e796d2cd23424fe363c98c2fcad2f84d83637fa9ce641c10e2d5154649518dc8a53d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h625ddf4bdfb6d98d8bdd92e26f760a8000ea5d1aa31264acd4f806ccc4206142cd4922ce9bbfe408fea78d32ce69fafafd3bda4501afdfe228480d77d5e174702819ef09c301c4fe70ad5ba02255cd5735a1db3ab7e9ee566964d0bb2b3c44b76c61fc0f25305a83933fab5902fd21a39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he08cfee3136229d07665767eb399882d888faa795aebdb94c290e05bff1d65b15cd99af3c9f94e9ac9d466c453a4e147443fddff0e86a19f666ef557ff9a0795e0dd8868629fe389f81411ac295179c319c6afb7aac8b6b07a5a81d599f7d917ca79196096a4d8784509a0f67662a4e26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3258e1d74ba8c0d41437d03a585f89e9d3fdd5cdc416112fc8496baa435b8c52a00b9390ac134cc1e1137bf8f4071a3e24ac35bd3978e526e6538455e07f3bbe0fd23fd6e5e62bfc5836d62da8d929f249e24f2a63af7a99f9c943d6278815dbd5caaa09ac4a2ad38d934cf22b573fc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4db15c213e9330300bc97dc0ae328689863490daacbff335493424dbcdea5288524789e04d5351a6f1bcfee89c081d7884de940a8b8af6b40099c26012c9d97e8e6bb7cfc09ceb09df71ddc34ec07476473f24dd73c27317b086299cdbca7cfb7bf785bdceef8af560fe7757168df9a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86e524c4a254244eb70f5293fdfedfabd6e0195aa023ba12c6ecd22fdbc9bccdf01ef60fa36e8183ccac913be1bc800d5476fbd9310a33dce4d5361d3073718ad85547a6e03f49500d9454358ef9889988604a090040c8938873216196c175c8546ca6ede06dedb97a445cee79cd17046;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20b25b42afdd2557adbe171e9b17b30ce5b4f17780698661b7274223170dc777a7eccb480f37d79c21f5608e0eb1633431f6a5e0dd9673e36754dd5e07c2cd89bcf03038b7869268e85da301af64aafb49717b5a2a289e37158f79d552dd391775b173d2d027a1df1662ad124c8b83e49;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7727b65d40f3492fb5e614ca2c93881b9d2ddf88a45dd26b04565053e2f895b02c137913551fd3187c63783e3e0ffa3aecb3df0ae2e31e461f94f5e54049fb01f7f2b8bf680b6bccf58b12b17c77bb094cdbc8db408c6dea78db6c95fdb4b0dbd3e77770403ef3cec80b667bcb200b8a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7afcfd11b027348389ed2f6b726d42ac0d1d3d40aef1f865f34c51a22568c51db6b28761b766095f29cf62c4fa2e76a06169f2476c4fcdcf9e2f6040db6dcf160c55a761a06a84066e4c20ad79009926953145c7614ec4e2e070611a8cdfa7b47d9d5f81f8e5d87dc03f6956a3275cf89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1e9130d01f6fba58898c9f05c21ad199ec4716d083e89cc2dabad96d59110d0500763e230e694754249804f00367295260e790050d57b73b7900189f92228678e89e1b54c7676e6749f6eefc39d84ecd04575b9e4f43ef8f6a2e96f3bf89bb6dbb76982ff2bf0089c279552e71efd3cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d58108274a53a6af4cbdca210b9e74e5001597d89fac406c7736b44053ec7d722ac83adb275be56595d887ee891e7e002d2dd524c843ed6193ab2e68c25cd41750b6524e95302568bc596407a941e47b08b9b6fa50148fd99e9c9804d195071910c2014e1e029dbd1795b415ee7646d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8fbc86a729720beab801f03f477dc0f343f7e24f8e681b63b0f977d0de310c117925a89b6084ec9191e7f4ca942605c1aa72680c83a901666370afe3dd4f74677eee63489d6b3f08326e912ab3db701e67b4f7f14f67fbb14c5908ae9f6c9f9ff5cabedac11eab8fd5f89f9aff266200;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56595b793f9cad43076130603cfd91e94f7eb73ff8891d3a8e8655b9665488f58a9b06ec3dab563255e53d285456f926da596f8decadf354d6c2501119fcffb6f9bb74bf4180b0dc7a20047d94950b3b7d0efeb3e61963dbbe6c03b2f2a09a2a704f271b878a497d9cac0d27554d6a596;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b64cf353acf617aa19d4689cba3da7b35c11d1c921a26c38e280ea09faa1409af6beab2aa0474e632c8e3909c169a3ffa183e4857912aaeb579c7282995859bc163c68209efd1651bf1abd3e265d6442997929cddd58564a96902b45abb33dc182921c4a9e769d457eca3cd8ed6de464;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h721305d9fadd1c5c6f3b3841dc081fc81031704d99fc1732a14c9b9ba716ad4867dc15c4cd12c4fa8bf1b06313f5247216d2cab14f830871507f28848edf2afa98e90c210a91f5e5d4cb4f235e5224d40105d5c8d4f54385dc24bf8b890e8c472011b5ed0d3439898e00400053ddd2851;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeb4a53c0540e8500856796deb220d81688a911c9360a49f93c357ed8cb8acb58a7164885259a8b06b605ba04506bb988b5e6e0448d10633e821e928fbe9824f683eec160ecb93ab04fde8ce2057c8a7d87fb5f69255ad7bc5cc0ed76a155eddd62e0bc8038f47858d8cb49c030b48786;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h457509ae4d0c4ec3ffceacce65a2982f4fa70b939322c986b3d42d19e628ece92dce6bba44dd9eee13fc8ef9e337ef2d4cb2d37e9d0f9b0f15dd41b64628704070dd41227b3678e9420ed65f6a7fb923260bf38fa268494133d5879669c8cc02735027efb28aaa334e1e2c66c726f0b01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6be04f935b19f8a7300dabbc4344b3b4104de92d165c3f3b87b5b7fa518775d8030701b2241807d3b0ff39ce19e0abea9267ed61edf9b02f14ca6633bda7e2131e200df7da10f8736ee431c39698912d46f048929931f6a68a7ca58b016204a91b650ad0b4e41e0c0662fc471b331600b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6588b1e55ab5917cb789880d935133d5b59ebb0a1494e7ffdb5bb63e3949b4c641a26bf5b943f094722f4e6a4da307452fc7198dcbc211fe58d4d1b560ee0d453a7f5148a7c7608f12b81af6b3897d18b87b2cd8327535e584ed4ed4be6e03011065d2cc8b51db0df36f8395614030e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4049a9951672d27fd7afaa00ef37984477a315bf1fe4466b443f4930fff6df3d7799555855ca9cb2f0274b63258241aaad57945010c18e5dd2acc7a95300145655d260facaf013a820f153c61f73fe59ad41194851233f358f1e434146808716214b116fc8a94a2f92c02597b0ca9de5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h263cc56d3a6067f508d4c92978ad27adcd701d94c0a3ae1090eca8791566fd831e7ee7b274a29d2a46e02d4fed520a67d192cdbb9b2020d50eee175ddd4bb46c1261f2c9ab768f0526bb41037c4568d44624c5b47a6bd7a32bc87f27c7ca35ab66d62fee6e5876f72ece6642c13f88d48;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heddeebdeb2daeecb5053a6ccce871134353d0fa1302730b50c7dccc683c7b06cafed1d8215ce1798c7d13ecce7b1f474c9791ca126d4c89b5fbf612f06e0d863aaa4edee32811175a608b59ea7699b86d5d6c00c9fa88d8614ca7b19bf912234d285081b34eb4b095b32b9748a45f5d1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5c587ebacb013c609ccadb8fde8f0fe3c0b7afdb20d0fa71e7e4957f042380af12710dec877a5daa3e11ef35af97519d71e402f7442f79680ecc9fc514babd34f2bc4d235db21c5a9d6cca649a3db204313855bf0cab78b3be9cf8150519348902644eee31fe8871d9b0564634fa46cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8963f5750ba8afc048a94ae60614b2fb73d1606f47e171ba8dd37cfe130f298c4037fe8dd4c6fc3769ecc6139f776f4905328427ea2a15fed1611f64c150f37a2c6abe2cfc1cbfc1eb793e22f4c92d1b197d09193bda011af943d53f312365c116b2394e638d30be25150819a1fa87f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab425185d30ac8f7ad083f33444c87177893fcab1f2afa0f969caa8a7d6a0bb49c64d883dc1ede1e6367743d9f1cae1af2e0cb6cf4646bef6cad91c1b7f71692ebf44925ef453cd9848691fa8d694490eb165c99a2f668b7dbbe93351d49cb9eb1e423e9c1e7e27bfc882b96a132ee6de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb609760fb5190e466d2d676bbe76e65be27bba772ace65c8560cca55521d404f5f522855ec29e38fcf285e38e56132604ba28d85d08c14cd8bc7d93189ffb840ac77a2d8ead52fe9131022936b38a8255bfdd713d81b1b255a9dbeb53457e52e9ecef8639b44c103234f0d2a82f62152d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5032ac2fd182ad7215680f78e96a68a27787a77f1ff1e12f43c8d3245e06cfaa1a61d0eeb8879f420c808aaec7e8036c5188a433193f790b330d667968f449d3843ef8114f29a705180d075bc9b1f6ad575b2cf0aa60a3771d19d574ac52419b3365059b8beabc35e08b814d6b56783;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30800161c4ae523bdabd93b2ac950a7292adcc114df8c6289143e0c85b48072a4c8b72c3a51ffc7bd7f32f436328ccfcf28d989a24feae407f26eb2dc27261ae6c0d24557db2471ffca3fde1e22a08788c7cf0ad411ed8c364ca5ce3696e61bb235fb144e820ba6db8628691b4e2530cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d26d38ecac9c65107210c420b43e6cabc9fbb955ee3e1abf8d46e11f0ff276a00d405831126aebb54ae07fcb5f29ad62f65f0dc8b17e0970d36b6850c4a84889e1837a604849d2d0a9e2e44998e7f8126c40a0815a1683e1b08057ae4a55195fddf1e84781eb267d82aa93b22d628391;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4a43d2e12366aae7f0c7f5feefa92aef2780fc5235515efc6ad64991a8c57601fb58ea03756c37c0e7b241621eef6d1940bd59c3cb4934f80b9b594477cf0f55fce79b3fa8b3ab8aa7f002d706e6a2e53a35b271cf36ebdf638c50b6979889c74f400a37ac9d884ff908f8d1516056e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff1b2ce49f39516fd78969904a495762a6d6d2d66cc80ae39979ee1dca1242ef141d0ade2d743a257f94274e64351dea8e4210cde7076ee09a216d6e62eddee3a1399883c2a3f011f8052b7babf95c5ac8b597439cb3f1716c6c0f076de53956079065cb476fe42765515d9b235032e9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h157ce53063e73ac94b999259286616d7e5ed808394b0f22a7250c0507c8f95c16810f7e5c75824178ce8ea6cd0a7e35959bf523cd129482009fbc6382fd3967a844522686965b9e56deb3753776dfd69215e58a5139fe7b258b83c5e8438feeab532d6ea54ce660f36ab4adec7e293ad9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff0eaac14e03b97ce4d5d8ced14aca5eed0382d0944bdd3177aba965cb509cfcb6595c921269d9b86704fc105cfe37a5b047a858fcaacbc6a74f4756f3fd5d6a651ebb47ceb38ab523b1d72c535e97524296899ab69db0b956f88c36669a6cb8b397289030ce9946df9c7c5d325073990;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d449e9f15f2acffae5f4ea8d10abfeb2c6818bae47c9d2c87a8a3a20bc22db8ecf1c37ae8d74cf29d7edd988f58ff6484c2ae33cec6a3f37b0d80534958bb213a730bd9c98bca746e810bd38c86cd307b7a09ea43fac07369c42efac3c3c98e21d44d5c126b022ed6588e298e2a4d7a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf41a9db92e0fcefc5517d9657c7730e6a319f11bfe8443de7c99852d42b0680791c44e6d5ad9bdf3b81089956d73e4f31145230e9eb77cc029ccd8e8a0e49a6a3cf89b610ff0373b56962e72ff3e363144f5d3dfe1b1ca722f3487d1142935117a7427fc5ef771529a1524af382f941d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3c70d5aeb97ca08a3696db25cafb094b22c638e845ce0c0318bd6640119b3401adc6ce075464cf7bc506d6325c6918c29f944cbf6f69ea4c6dc092605b26537e5a6653a627ea6c11025381187cc52a99e2e270946d4897943b6b386ef6311da0788e7553d7d480e16cc20afc2eb07dbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bc8ae031beb5f0ed4720ee60eb01d7619d2642f2cf5d35804141f4fd6a20d595a314389569e91179fb04bb8749753a374f4cea2537defc4c4307d1fad12887fcdb5c0fb084e114e123be735c18828f6b1222e51ffdca512bbc38300d4f6b7e311374016aabe407ed102ba772bed3e9cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ab219f65ba15b7245481b8826e22a1ed62fd3fd445dc244e713ead9adc96e7d4fe09711a34ebe030cf1bc2cfd2982dd44141b6c8be8ccc94fe3c8969de192ead8d40a6933a593bb370059d881f254834b343a18fa045ad9a00fcfd30f6f6d859527e9c30b86cbfa3e512c84670cb8554;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a09c3cdf10b95c74dd7c7b645e58aa18abe792f7366207ef9ef79f0392131d80b428d1c8729a9567fe6b05f78784bae8b26acd7574ff3c493cb9d66b514ab8e7e766c0c64453d3087622900d80e2bd43dd1dd402fc4799cf9d2e1e3f8aaf074691983d31be8a0d260b465747e8195f8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf5ffbff76b91472dffc1d3f151456d5d0913b1a6084bf63f0f05d6e84b0be131eea52a5ef6cf4f96f31ea220615b26f2f294b59b8df3d6294725c3f10733d55ecea73ba811a7cd73dfb36e30dca2a5f0df4863a4c9d2a256e22f4be0a94233684f6ef2723ac1394816088232b9ba8aee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h695c598ebcfad4e4a255aaa6e946988a864741afdce72dfaa43cd06c6d03d22c996532c756c170603c58675a6a1add0db746333405bde6b4f85dd89d0c8fb9c9ce2575ebdcaf9a1bb117f7d7224e3138c8ea268df04a258d162af300fbab0e7e53451e8a6e62b13b0814a03cf69260614;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb276d8756e29cb2779fd11062ce6998324f80219b1b72c722135676a6c8ef5bbbddde762ccf53f90e254145e2cd009a93b360b7fe904ee61b535a557fc058fda1af47b5143d36cf9b71e9e7bf3be74a4498a67c418495bc50492e008150d3d5ea2162072a4dd62142a0fdd387fde82138;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf2be71f9226448ac54f21e8276e09588890de07782abac525d402df9eefd41880e90cfae0c9ef40ea309518d1a7c798b5a07fcadfbd529338686de702e7040e12445947654bbb9c6863ba7d9c54b5f0f29b40e22d480dcc09253438e28936f5b17bb01ef8abf7f8f7c9d06315eb638cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he51e42f08555d70689de277af4062fd7f0cd1e3e858827c167b7c5fbaacf4f4d3593e663c202472963cc3ed809909aa93707942a85f185b99c173e4fa0b1dce1b07382f96ff94cbf2b22cd4b1ef0deb482b4dde32fe4c21042a144613e7235b70c267c6d80e12ff71376a2651e3ce741c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78c4830ee66432ccc1f1ca23c2e3c1daa393310940a3283bbebba0d3ac746d4622c06d76508a65dd21f67fdbec69e9bbdfbcc20da8e98fb26b828989af46c281ad20ff6eba24a498d8f07c3f64a256423d264d4d0c84d3486b242508084fac01330ad26bb6c2c2da7b4bc5626c2c65e4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3627585b7a572fba5e4cb855365fb845239dabe3109de16f1cc94303cd71f325cd7e01291042bea24b0760bbc035e656e6485fece1ab0e3ecd810360ec81be78e5a29f5ce2ad2f36197d5bf525f164215eef8b699e22f1637ff58ca1073cf483c8d486353c00a4c1588b59a267113a81c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4825498760a80eeb2ece3289b361c7ebabbb7dccbaba54e4482ca488c7329903d950fd977343e132638ff982394b25bce621b70172d7e1a24438e28f3f21e7bb79009cd1117cedd14f3bba4e2155b9b3e74627d20b3e4df64115fa07569606f59563cbd91ca2ecf2c913fbe429a0e2add;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h941ddeb4b218101379720d96b406d390ddf20bbf69002bc438e287d3c6f7ba608f91602be215806734d0750e86c5716613c0dbded3cc64f784e2dc117e1958cd9a33c2dd0aa3065caa0a09567c8add58caba7402aeb53e1a187913b436da966b3daade7b3babe0a7bc03cd22be2da79d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda5dc4528b6378f8f5a286c083ff313ea4374a3414107daef92a088a71f5436097a85e98a28beb497bccfa9b794ea459a1dc930064bd3717d45d3e261b1285730f65fec44652cf4a4e73fe52cb86568bbf922a95b4ed3d0c797058477cbd75540d50c8b47fc1d81e2fb0388abf23cae63;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b4b638eedd55e1e98817662a75cf918f0f12bdc39e515bb9d5d497bcd3573efcd15f91152842ea031bf35d8a81c4855c9f1f994d5c8058a8a3012cc44c873e74d96a82d4d8f99a80e50791296896ae19f8f8a126d0992517986575bc460f6ed4fa7e5e6aa650708bf5c6e76aee8f1d50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a06630963eb2083799362886be48d451f97e8c7a5d60bb438795ce1c9e62d7cb18070d538033b604e7d8d6bc877a4cb14de5b2ed34df5e3c24bf9532a6cc1e8aa61506688ac4b18e9b778cd1a5a40d4fd749bc22f60586c0f200616a7cfbb75615c7e3b29666dee703ec894125c99188;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76174658a349c60ac420e708dea0c22ed8b390b89f222ee6f3bacf5558fcac913de4d4d66bb20277481f1662611ab71d633935918ac3beb44323ada569f5a42372a045d0bdf7a2430c0444f66852a5fcb332d36c49f3b7eadf08883ed78706bf090f7b971bd379ef1a3f0b43c39615b52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab5f6736322447db18a41aedc0a738bf24942be367639374d1b25e4afc1bc19aeeb441ccf68a8b060016f7bbd44185a163c006318f49615b8eaa159f818bc341ad4018afff55ae2c0329eb514d4be03547a298822a2e8a09bb48a03f3a0fb256d9b978d817bcf54b825c6cd6300c1f614;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e87f35fb57729849c4115f53bf1a80ec618037c6efda746faac2022827f789c7f0c4f4f9b3673016f5f20387d4b886cfc7ac1798245b570839c3d51bab8d1e211dfa8263c2bcb0128599d1f858b9092a2bd6613e676c2f69ee61a5a291588ebbb9e4723196b6b21d715f8ab24fc27a1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h683a1f9cb3ed58d7521281ce69d1761a3fef34d460b2d11d415544f1747cc7225ac061014b8b616e1fa166d715a7d6569574264af6ad1765f104bd0768837bca67888e2b687fc0bba8b85bafe393206f6d6f200e9a6bb9be86a28260a928698f5fc754c1a624cfe58834957b66479b235;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65e55af937b1219ec3e4a994a99065d6d5b09d021bf59d33393be35610881190d707ba36aff878bb3eebd78fb984e36de2c4aef28de1c013742cb566e413fedbc73aaf78fa34077f174c0b23ba6b5231e99aa3f9c6ac015ca6e3103172a7ed8d810cf5b16b72535b8a7640a2de499bdc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fecb0570e0555d3eb46c38b9bd86a2a179c6eb810256854b1b8ebe0b3368af4e3a67e864812fd8c76d76f2cc8f45d841dbbb129d231f3c7bede229a97e9f910935fb02322905fbc4e8e3682448bad1903c0d7c057bbb2e137edbba3bf37e476bb9b0a7ddfa2d5c23aef567e78243a9c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41532c088f787c40ae3ec234cc65d4ea03afd08b9f878e6ce1a4062505f61904854cab5c0bf385aa8733cd7905b91dc262ad366c80e9b0d8829af43ff4c72325ad7c35f027560e64ba06fab72be3e4613060dd1ef0b5ab2b0d430383756193005d4ea2d94c5f5fb008841e7c96d23dbd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h863f972feb604e95d8c15e66732ad04eaaccb1e3b5bd70caddcc9a06d299e6ce63ad1ccdaf52f11fe9c354a12d2d0bed6b747f18a2a73e5f527a9650a4836e3a88c1183e64ffdae3f291bd8356153d35aad5f63a1360f5df0275185fca28d0fea8a64dc9ea86bf579d56e4ebaa9e9c7d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32235bd7d6387b6a0aa2977da2be76a4f4ebd795c3934efde788b475c157421bc6f5da6bc9e71b2b9b6ab7b59d8b9d845c2919c54e7946bf3b9156fdb906b5d4e25d6fe76735fef78c4f43e386d07782425d57c65c0537976ead519ae7e5b8a54d92df7e4e90d27a493a335d7d0ea03d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e0a994d1167caf5f80da8f0a02e0224e6ef278510ba83c2b43004deb18af0acbfce78de6525501fdcbd1a00822dad015a8c8cd1584faebb51b0f7821a3d0c7457f58299ef0302b360fe703eef0935e5190ee398fe94ce660a2db4c1d0ffffcfffbbd8282ee4b73069a2c89045a6f2d03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h138f7792dd9b253d4fdc0b531cf7fd5cb735bad41a8959c145ec2012d3c01f354e55b511345097700fd17fcfe2b312efd718e394a1e810658a73356698ba2776bca83e18ad6291e25392719ff779c32227883bb8f2299534b6baaac01500e36b756ad45898823be18d3134d18015c4ee2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc34f5ed7a5050fe633f2c5112b654dd2e621579dbdf727eb86ea11ffa786a9ea7a7381d5ff1767b32db62fdb046b920e651210ea9fab2e09e62aa803168f94dd27360551068e3341057c214661d52f2231c66f2843b6ee72f1c6bf7f41b7c46c60f32569a423095f758196d04265e267;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a8f9981cec3182602460352e8b45eac7a79bd40b3ad3c2c8d0adde5205f67cb49a1f2514db24471c91358201c46cfebbcdaa65fded3903de65c8e9c721668aabe50bb8439ec8579b3d6fdda0ff5c2603d9e4b893da1f300e4caa77ceafa833e469290125a52d3fb631a7cb7e4eed896;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8ed60a0731442c9cafea5d9f4af372c001bc5cf7d1ca73f931892f55feb5f20780dff43f7f4ce41c1cf0424e6131ec8e53174c3d1efcf9f2ee9977e4827d5ee045ad9374b848e9e29a6d6795cf77d7dd16b05049d1b2039a6ad6c789c089f4a35182c2a6292e6f95a36d931599cde092;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fe97fa431f51f40f9d3bdb40eb885efde13214be0b187719ef7e3f8bb80d0acd6d3c8cf685ea9a5312d41188999cad713d54a643027aae24c7fd9b69044ebaf31b2e1bf4c12ae9a3f5a3f57e8cd3349eafe7e084b8b691ee8b565406993f85790e79c5448a9674ceb580b937502cb97f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfae0493ba4e6fe5cf7bd36511a54a00d56eb2d7da66f2238c661c172ddebc07e62b5dc47da93d0a712ac4b98211abb047a891ee0f514b0d1c949d7c019b0ccec327072e7a00c9a7f01779ce7aac802ad60cf935316fc32ddf2fa13993a6d0bf2f21c4b8134494b7377ac544ecb5bf6134;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5cf80c104f65215246c2c14aad17289098c6adb98d0490305ec551ccbe99591b9db9f728b2e6ff2fd55680caf3e6e4b21b8115284ecbc3b57b3d35e3ac53365c6a8b551ebdb1cd65b6abe034c50eb54b4edea1cad9356aa7fdfd090527c8b3f33c5e8277815fad062fa9c344f8d30ee9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h509b4dc4aed1a8a69172361d0f9d8930cffe219e4b15d9752fe7868b7da63c3e8b724c4cc0c6dbb77c130ba9bc016f0c5920446720b2c9dba1cfe54acbfbddc81a843258f3876b8e3ad8188939fb62674dbe7cd867d86329e2d641246b2ba1d3048173f44e6cc37045a76b5cdd1b54b9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha32b15c1834482c097df687d8da19096b441bb611b37559bf446e40ade6cc14eb131a397e996a222185b1757ce005ab4e8c32825c5055eea7dcf4d282071dc9050e220c29f4c2fb90cb2842c0414394363571c0d1f4a7b0bee83a519f1d84aea964139690cc2e067dd0204e8402b10acb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf959d43276251ac45bb3ad1c902cec5aecda766c43980c16fc0634d93143756001fb22ae9ebd8ece98598e18e4df717ea029be6913f3036c5bf729f8239dc059079dc165ededed018df52c18a22179afccf96fec189fa71625713463383144a072fcc5bca5a416be02a773056810c703;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h355b464c5e8fb0846fe55397858f69666287b3bd1ae896a726b3508434580db88f84957e451b6e627817067f22327ca1bbfb3d4ec6934ea27f8774ecb58486e5fdb324323ac5042de0fa4eae148e28bf91cd094971e636b879785d049192ee2035ec54bdb6a0b75ed68f37d643b49bbb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56aa019b888dd9ef4816ed54d41a05b1c0e53fa7abe5e33abfcb885c8c3870ab4a4c8cea1a37bd2051334b577e35c744542b1455507fa704367eb2f1372436908b125e918bd00ab7024b51771e43537e146a9748b7e073a5a0d6d0351fbc099ad454573944c003560cb49d11c7a5f87d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b641d748068d54755216c63c85f0f525006b722f05c3c22fb7c097fcbc1e965d38047259cd367d490f73d62fbf4e61246feaff4c018b17c083a721b4d9347da993be078932f0b7721150d21da6ab71eaa97c38f41fe84e0ee02f40db0b016b2caafea9241f8c3e10b218c580903755cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2092e955c6428aff2a10987df9077ebb94a892ebbe0c11e4516a045acd12c03a4272b3f37b22b06e2c46c90f12ffc0811b73dfe7f7d24d1c8fce1bbed532996055b3dd5137d6429138366040a32087bc5467cfb30d3c62f34184dee0a42444fdf12fdf63912aef564bf8ce5c38bb1b04e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he03d86ab7eba289b7cf6df35bd47f58e20563f851500b8bc1569c62336cceb218ee636e8de59717a395f05a0f816642754a5671a5cf369ec47f466d787bc528c02047ce813cd9fbf0339fdf474e154da01b71bd7f5e5909a39d4a25081a539751fd9028e10b4e66e637a94a021776abfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48744f18e089a00fcf2527d46d67851d34769a721f1632d91766e551882838fd50e9cb2f0aedbd3a5df4d478334c020457969526c524577b5886cc2b23c0008b8eeb7edaca5db41397600af78cbfc965c90d8252c62c9f48110a435955da9639bbbfe44e137108277b408511a0d1f6e1a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64a18c2872754e6aebf060173bd7301a30adef1fd0e6a350296c675998473b9c2037a789b8a979768d0845ec452ac89bb98593673cb389b7e7f3201a6078f96b53edd0724d6bec664387cacffaa9b92b3b2e285675855e18fa20715b9cafbf4c34ee9d38cd222dffd86bc53ccd786b92b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d8b5d21f7781275108d0a867d7148ec96437de81a2486eca349493e66cd540fcb493172a43c6e526abcad34ed5bd45172f542f256068e8339b0b9566fd9eb37f0e37c817b6b5c5f464c0cc5698dc82226f0f77b0a6bbbba2f215b6e2addd2ab14eb4ab4be8e3ac50628dcd6b1b78bfcb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbae0e0bc4a815a5d95dd1c2877e55566689cb6c606f204f7207a3ac7c50d1f179a8db61ec68e83398372cefd4f95ba9a784cd3190f9f510f232f1ff27a1ad3a22e20643cfba5832665d24104f997afb4bbd8ac1bcf68421705f381c39492b85623c8040b9bd8d209f82612c070056da0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha147fc7c37b854e6750e30105698d2ba0b0f216bea6eb7b5019a8e97b782e7e65afe38f15a8d8c2c7bede79105ee6fa3c32e4f8c43f15e17022a5fb39c02e6877135882b45a1559ba2c68d5ad72163d3d103f0d3a72978171ee68002facf8204bf0e7a754f5eae3aa2b85ad01c5d5dde1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a2047a31212f4ac268a155393391fea11b807219e665c238b513a45361d0340494196354728a899092911f03ba619f9b401ea6d29192c09d3bf452965ae02b9b07dc3eee7e3858e343cd21f88f31e2beeb4808065841290c3ad2713d8b73704f4c025f1a0c80e5380fdd72349671dbfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa61995236cef1a01f31442befb5e874af7e8f0f43d5e73fdde46688e9d0cf453c3ec54f43e2f13e7efef1c7af9a0da496ec3fbb9d4e8f97cf088967842b3c3964180ad907970a55ec99aa83eadeec485c1d969ab8a24d96532df1efc59b4d4e8cc3d7b1227e64a9b925fb9e3349c5e5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aa50e0bad2a32651f6fc4e6f33e3b4282800026a3db8ec0ad97281cf5c7149643b8ea1038ddb2ada6aa70989f1cf2cb5decfb3b82ae31ee5ae79e5fd225156880fa2cf93471c3678d4512940143332587ab60d96ded7cd47fc3e0b064e93d6dca13c87fe78e19ee1be1988f5a2d12905;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbda648cd67f7a81572a41bd8193145324e2ae669956542e4cc96ea40ee2edfb1981285a67382bb7056d4930b7f424216ef938f274c17d6b25aab068f88326f3557ce5458452976840303212c83fd10748be29416afa43ef570c865d88b2e55561b6f5450193d204d945ac322bdecbdea4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f94cbdb8d610387bd19ec839db332d41b7810fcd26bb630dcc2380cc6f8eea10e1a5745fcde89cafe85beab1995f202ae4a01799c6b583bf17d25bd244ad55fb6102a5eceffde20898844751092263ca2a51c8e5bcb05b9255b32982fbaa121457c09fe85c2301ac54879ef388921431;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba13a4322fb0602a6b3ee167941a02f191e3af4b761440b8b51f2632f2b9d061cc90f1538f552ced5e90b602452820cd47aa8a3b1075a7df81d1f0ae90308df8d9b398847931b8b8c4221b3cbaf83ca3d494d125b04abe85d1bd6f9f6222e126b9c4086b40345efb750f5870bf31f37b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b6a7cbb386982af9823e994c62bcbddaf37869c7e180dc32e0668f63fc0f70c83a5e562db389267a80b8004d3455ff49163dec8eb290ce0a7d1e34b31680bd21cd78ae88af113d172b2aa7e29947ef49689a582bc0c6a9247bc94a2902285d1bf801a4a08fc78e845a34dd436305cff8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b86318694bb69720961d9d2933327fa9f4fc953cd3f2864a1d0488fba930c00d9480a804d5acbfe56403c98947a4bbe5e3b690fb3de1d8ed1feeacc60070f7bc660aaeaeb2f0dfd2fa599a0e321a387d21581523d6437e7ebdad8b216fe7219c6e8f92f5517b0c6e9e3eff7c8951b808;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb80627c49a0e84228af4eb354e8347c4f5e8d0a66311d5d2c1d950d3c9b2d0f05e99738ad90e0392fcd05964bba0ea65a9c3ac93e9778400c9986b49a940d569f3fca8f18460c8f0b7c69fd88b92662ed3ba1c7604853f70bf128bb755062c4c3f9ab2b291a992d722ac5d54e45e19754;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47ae5cf825154276220ce2b0b12321ba23ba73b2f52e64803a0a403cb4527a5176173040ef98acee1ba625d5d33f1143f80674769fe72ea9e6bd4135ce380345c96d93b83d4ae243df11cf6e3559186787639b3a1b8316730b72f362d03a24d9350b120d7aa7406c51e6593535e457288;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf607c283e8461c98c7da588600031fcca749c1e811f61a0ae093e8c8585a4604585b0f7894c84a88c7c7fad672515bdd9d76d68de0e7603394be1dcbc511c0fa1fd40d0ce6c98abd21a4ac1435db5584a804352b27196746f8c0657c9c7b6d002f78a2372e2ebaad32994c992b678aa7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f25fe9796fc9a6fbfb4ef6b7dba9bbca1b5020703b42e352c611155f5b8e809d1ba181422309a90281c931f47ebcaf9cf0ef27ee7374bef28702daf484b6ddfa9d88febe9c8f334bfdc6d0f82cefe4163f0cad053c9881087b5ce29e53a23bf5af30ca93e2c522dc0f42b0d2494cdbdd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h676cfbc232c92fffe02fd12547362de1dbddb7b54783e692ce662c7a7d9781e0d5aeeb458a1fb8ef4e2947d2370a76c904d810126db1e43280794ed1ff90e300c91573f506e54618a75c21a15838d59ec34bc2c48179dc90da15f9eb4b07b11140e4fd3f3acbc242cc5832041f0d1e6a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7c14d7a83aa56bc68bbf69fa396a38b638f9f724383a2fc3738d932ac6e7b1650bcd5c483166de05f378a1be01e8e452509f3fad5fdf8f651d5c891d195e748f4b09727872ec05e3672922385898ee5799cfaaa013e9416a16fef9449960b8114b7da6e43dc571a17f48b521abe24bf9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5c91e6c0b53ab35ea9c393c100ae231d35c7d3a4f15d2139f8fc98e8fe11c7694bfe6b3fe2c83e8657db4b1cf77f4124302484fee02144b82d8e89499b47deeeff8aa93dd39f8f852ca7ce617e1b2b52ef17ba0110e41da5a6854a9b6d49af378feb6603e3d58ebf163d61ef8b2ac49d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h745431ea1a542f9d988e956a7ae0bbd59a5904aa3bc4ff107d986f6348482debae294b795ff79f020cf3c77bbe0a0e9c8ea103b0362b69114db4124cdbcf3c41d82763aab82881ce1e69d6bd5c9dcf59bba58590ac6b1c05c886646c8cf38efd0853e535bb351d196fa36266ecc69d389;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d33563868f44b6f7f7261e7b3f3da83b481e913ee38f60ad40202e372f1f88500ad76b9b60ef724d09c0cf0f8038307e91aa856ecaf9d6d7f9dc0c9901c7bcadd5a05c21595817fb2d46f7d8168c2ab9ffd1fb1535530af20d6f33ca0a54f8c42f1ea4584aae970714418c37001b0ac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40931466a13834682d1163688be885a1c4ac550ebf0b1fa792ea91509e09405244f2fac81e2c634d0a2549e214c91f3c062c4074489c111d79e3a3ca537223584fd6f8d30550d682d52bfb6483e16ca04667ca5ea7f64188e0d989804682412f8961478a9f1f45ce4c13ba5c217ce46e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc3cb8ffa25d2da1a4287d2ef18ab46fbea9feb40a3819922cb5673fbaf229628e4c3eb19e486199d8e95a6b0d4ba1d01389db899da76388228df89ace64d7a88e5b77d81c5e5343cff63ea587a2ed0522336f19b7dc6c9906e89b56b8bfaa6ba5555a6bba162f2a2d36c5c81d52ef33d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1dec173ffd69809740000c95bd36a65ebcc538ac95ff30836e2ae6722812da0f3b701f84fa1c0f2cb6649f09ae6b1a68d491f1526b7d3c52ea6eb90e774a4f1d61db3e3245d6f8855c9a232d1069cbc30ae758e09e72663042e35fe35a9223dead5f730b803d3f9cc40ce72ee9396e0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd3c12997e197f91c8402de2106cf98b49011919f78d75474ae9d6972904fc7ce7878f463ab7ae9960bf1d05c6178c918341caa0b915da391ce9d7ff9542ad523735fb96cfe64b6cbb5f3379b0ff42fcaf8f9028ba45e5e5024fefad3cfe2fb2379c9a11feb47f0a6142b685b135e5af7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2db7412176bd26e1f082ace944d489c5a5f244cb8d1167ff5fad4d8e483cfee864acc761dad9e351343c7980e8ddc5f7aae822f1f88f61206e64ea76ec335ce39456f9d7e5f79c436ac0ad658bd5de971c3cffcc555b6a9f3a9c5d8446e944d942eaec05e28ce5d3cc93c6c10ad416b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8023eae44a616fbf7bbfb038e2db848bc9d593df1046e63879f21c7de6b0ac40566698690c01c7974a38382084ba5c7bc09befce92188a02772359ff4e2e4d83317177a164b6c51b3c98b0967e45172d5b3b691aa5c4c6953c72580ead59a9c30b8758521f442a733deea94d1fbfefd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h695c600fdbb871949889bf00c61c48a1b0eacb91ab00403dd4bdae2ac87058d57c799b319ed4da8b8bad8e4323e10a326a4cb0cf991e19fa1951d2f61fc4a3e8f87e91d743eb15d5822f71f34b78bb540b78b0a5762d318c8fbd98f892d3acbf6e648ba582f7d67cd73d21bdcb2763249;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebb27eee296a9008c2a55afe78d4b23bfd2e9bc442169c559b8f12dcb4284d2c154c68adad83aff9623ff387ada26ac3010d4e1a7d20fcdd1c194377f7cfe4c238f38da3363448e5005b837d811731e40ecf522012ce49fc572dbd48ce821d0478e8082def0d367ff8204853fe4aeac9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd29913ad2eb071b2ada538e805bb015b6a056b80f9bf23cea0d0a1a00d7e099f711a9b72a75e17f75f576ff8395e2503c821b5bd32516b94334e04d6c589a393d53d22babcafa744a11670e3e7a1f2da65dbb00bd2d1cc1a3643529d9df4be43b5b516dd029aa616348b1818305fbc7d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf63d30bfff972cb751f0b159a4b0927a55e40fe9355d3b0b2ca6594e44324d64b782e8f38f5e0d5a3261e40bd50e5bb0c12b023666cce6c9ea197dc21dbb4d7ff21febb6ec7d88af2cae419d171f55a717ba0427e7d7cbf04a248a9aff08114e497d7dd7630929d97c2af66e3fa42521;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80108f410e07a05716ea56bebfb0ae2772422a582b50e9bb134680388660b4bc5283c4014dfcd3bc84b25cf99e25bdf4bd424e11c4a1715a73162ef8c20d48479f647eef2f4c6c4f1f1138278ac0805cb1daea72dec9b038f551ac43a90355de5d2b65c06f47ae5dee6daffd570b82bb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0c8b337279272855ce4f02f20e6b978269d1ba246db592f761117e6b5803dc1a1b958a307bd81334aa2dc54b3deffdeed64172f6f745832677c47316ac5899a6d292fe0a945527611315c5cbcc71230ced865ab9c97aa36e61ca06cc35569a0d822d20930f5fb2c24d32d83b384f266b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3268da953d6dba098f461329ce4e8718014eb0c91fc4196b6c339a142443370419548fb720733fe59f5a784e9e39a27659d6d967d5405e49acc1d21a6a2405a377471fc2802c76d8662062de279601290eb50f52707f8b2d8c1e8863b1f6120c10900a09b1db0577f32db8ea29354263f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h967719c27ee0353e4d71c09305457de2f3b6e3359a3018911ee26e34565118104c2d3cb6b828bee89c87db430c0ef27d8d859d55ba5529c96f56feacbcbb8ae39b361742380b9753ad42390c8e468c0d74316811668cee908e02ed4dfde27e442172edbb097099eee3cdcf7b5038e7cef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcef1bea72602b647d635e0b8a7aaede90100613b3534793f3409e696f11b95185796b801110f20fc1d7b6cf3176bc7a01a75e4ea194bf835fb5b84be3898d64fbb0e68bce00b5fc10ca75b8dc57d16cf5837bcb6fbc479bcfd0d9f645d62730d2ab14ff8f7326cb30c2e0cb824944ad6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6795ae557f8affeff43cbf8687cbe5cf66102179f409cc4a65847fe97d83c4f1946fa20d9065f38d2f5c1858f7af9ca182cf55ffab0864fd76fe9bc60e0b70b9b4f0be34d41ce40f7200890e2397ed8ed6edbf0527af3f552a083cceb6e2f35348824d59290e979357ca0c5f26b0d9389;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3d894f984ba7fdd3572df5fbe5a4f84b55ed4d6b448d4d0564610bdab47df0801d99c370fd92aec019cc8db23af7dc41e8639466dc6d05059b6ab64513f5cebbf87e07014ed04307c21845e1e9d2ac848d753314acf773ed9f12b9381a87ef7d9b196e721fa0591043a2dd1f4afab393;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eb7d210105eb6ca9c68bf55a9ce6c34a150410c410ddce1b93cb29e5563cf5760db03cf9482ca6e7fac788254d269dd7681bbf5551713a32de6b480c96ca73852b607e5edf61b62cda3070dfff6cabe92291bd1e740a830d84ce34621686437a48d78a0be9e6e8f1edb6d4ac8662b5f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6699a8821d15b5a681bfc0932c179112cebfa0c0a7f4f12266f7eb225cb7379552bcc2954df15cea0812c8ca52cbd2ec662d16ae24149ec96dc5d13a1a45291eee885769f8d8712802ed7b9cec6114bb8d50292d279c71263f09af1f001f866639a0ed9ef2e45e8de2116d68fa42b9c4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7558663b792c840a605441cd2b7b427f4dd17bceff00606158daa9a693bad0a9dc9014b2d0b7b1544895122e4080c53ef13d85863991ea552a7145e76b13f093e681e8de78f276443ba2b99a40a6b24b1b58127719b34af588c6f2d58fac02fefdd3eecab352d758008201f38832015e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bdade2ffb52540263ba767f0a3d19bee64228855d6494207beb64cc686eb3eeb6c345a6fa6bb10ea7aa4b1da785d2e9096b6fdb5b5a762fa724630fb2553e3a246424411fa75c8e1314a9c71411d141a79d2febb778bbda4df671c8ab57568c6209dfcaffbd6dbd5f90379129d5b27b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25513188af11e5e4057229993bf092f5a7b2cc7cdbb6a8534359630123ec91308398282daf4b31eef35d6c5d4b78409f2a30530c3c7502b2502b60d510d15c9996b55478f52bb12e07e17960238230159eac1445c4c4076bc2773420d962fde9ad9c46dc678ad722828a7a1878701b82e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h997efd1bca77243b1c02fab3338661dc0845482d8b297b477ff8f48d6946436f2f19c7fbac5a31f26fa98d14604176f35e8707d3e50af1f5019d4005d66abaa957ebae76e3018458208e1239e080edab4566ef6065d809e640d9bd1fa39656f228a154ebf136453c2ab29d828d18a7d8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b30af3cc386c21f65ee39bf9f55ed1dea739274ee4203132d66d9f95f0b9aba4b062cb82e58cac279f253b38693a3039465e05492127ee5a3f9a12dcee73bea13cf8f38a484ddb054b17b35f61db319e52bde91dd615b23126f57d8f07a4b5ca405694eb80b03fd85c9011a8961e3654;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b9a3a4299f32afaf30eeb70d375d9d234a769a6645c14e746f66a8bb2b1301b56b51432e97829afb108e9264f880b194ebc500a8a2564cc3c733cd651c0f23b4a401d8e1189a473c520c634db51f21533c79f21db4218066659b4ee857579a4cb6a57e11c5e4a395118a42a80a5fea87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a5419d129dc2de818e53cac15b08ba2bd2aee9cee092e546030e519c21aecb9c11a3ebb745b2c73fad805420dfb9f3069436e5277ab37b65854a95358498e205656b27d6c377fe1167c86fac3d68f1969c98ef6001fe4b0b517d93ea0cf8b185cfd40d0449d27a561e8f2c8e99ecac4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7189c9f8a5d921f69f023fb17c5319ee0eb14ce7d6a40d852e40196ae160322d7039c35ee777c46bfe842c3616b08951da8234b70540849fae9f5ed786476cb528f58a1e251962f463d720caf2454b6e99c77d83a1b637b75ab7390327ec7de8eca7ba73ebd9c36cbf4054eaf2359350a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb64fabe3ee77f0211dd43bc00c602d0f2ac262bde80794725395672ec9e13478007e44d66d7c665bf71630cc26e90f41b5ddc82c8dd428bb343c830f997964371bf00daa57abc124fec5b78db7f6265ae36d316cf65db156f4b316f44488ddc16a448f38931d1f2247e1319e86cbbedcd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc642faeec065565612721b5945d408b589a5698519b2d8e83ba40555b9c5619061d228a369decbc2fb67a30bf092ddc86c1edf5058f6c512318d81af5f548f1c7514803cad3a94956f10967434ef496a5f1bb8260b76f6b9ce3cdb4ee88695ab50865453c31c421912be7d8ec3f8bd28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f1e1482b27f5b651b3a60108e30953c7809baa21aa2e349c51189d8450e0615e7e98e3a216b1fd6381127a1fe765c49b517e4de2056550e5830ad33ae6c8eb178437ef38eca646e4ed8d9741a459f708f5c63cc4bef2e2de0d9c49db9ea3187db145564b3916f7cb45be41b77c59578d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd5ebb90b9fc28ce9a0d68da70d93aa30216ce689654235a38a782cdabf1071b7a2c49e0261f59d5acebf08709432e66b88d9d8aa4977a57407eaec7f10ffde8fc3cdb8ef384324e1188640e7f3c0b88bcf1d4e88a697e182cbcbdcbc6244cc623d1a1fd312356d5cacd578f6e2bb4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d5f3c68cace070e12d9dbbd4b822ede297250c4c8708189ddf903c775f6a4d46ba90b22da0c4d7ce719b6dccf35e2fd4526050793c56b9f8e796380abdfb0dad50ee79a748e33d418cc45e8534a47779ee6524956077a668870d855bedf9fd7b861571349ceb74454bdbebe475a08c8c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68da9228ef49b14c61942aca55acdcc8fe9df370adb3e964a034f8b7ae5bee6af2daadbe39c31d719f7734456ada556dfe59850c035755636bb0a82164c940e74e0c40d60e5981032994db1927d554061d43fc13f0d367e91191beea6aebe1fd9e79a75ac8ba95ffe9399202c91817330;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0640dd5db7254d76227b86ad49c5d144c1c5eb054baed26a4ec04ddb86dadc9c5cde6535f86578630ced72f878eed8b439a36fb6baff8e4fc1ca77641760a8e43ebc3767b4110654314a2ceb347006aee13113d77823b3464d2b1913e59aff996ee8048579bf73ca14f32bde60cb0b46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51caa1e4c3068b02dc3737a6e48caee4e20874e16615c8b44a8740938d20b43e45bcc8d6c414f673619307f798ed040f5f59c6078341948fe8f5d1af50d0766c1f39f03250ae83c4a441fcc268b3382e3a851652331ee11c37fdf16971e3d6d0fb7e9475d78105ad2cacd0b2aa3c7fb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28dc14771693824a46f03a9760397246881c4658ea5a830bbef7df502ff76d37f8ad157c099e4cab871eb2735f206c4ce56c4943748ff5a8acf0236482e4c8db254f739957c11f42462cccfe724572e617e2ca7fe3ffd9cc4317f49b19264d792d61c2c788243d994fe9d9dab37964236;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce06722f441a9f1279c3679619c33535ca1f7aa87f324652249975c1c33fe495a1339767ce2544f4c8e3c74c23de25810ad55ce0fda80df6bc185dee88acbac63dada9ae57223f8fa33ff462fba74e702b1a65228a1421038cd43dcb3db65242ad8c2d49c4e7eec44646bda1c01fa8b16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4a8d5c187baf4ca1d2bd4e45da0cd664531d2e8cfa3492873611e983ba4d25edb5ddc004b00b1dc761469b1735bc8ab369632880f104f930ffb4631548894fb62a4eafc68e68f0403c6acdfdd42ee316ac50cd233599c30b736fcb7c9b35fc27fb23c356a629c07dc7b3e2ad480f5ace;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9ceae8d0db8490b96c400e2b91c44746003fcce94e5b387c1674c10ae511cc4cb12231f3ffe6e9e202e9501bff530d767fa4234c6e6db8e32208fd30425237da8ebcf419210bf84e91bdbfe5fa6c0ff72795f35f0267c25788267ece4cbe1a2e6f1a3735acc6ddf44782dce08558d7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2343d038a371b90642b0da6f97808309d111b5a011c76db142f62adf4dba143118b2021aa47fcc96409dc8d158cdad4ec196ac7f65a6e00ab25436a2539559118ceb3e916534696e798b28b61f26e162ac290c9cd7e360cef51f20f03b06695bd969fa5c6308142ace43d117866ddad4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ef35acbb634e1b154cb85ae07535a3fc068f245804ea9bda1452c03f7dbcb0751de3331cb74b45ce728d264a71eacd1219df00d15ec1b61e722a1e7c500de949b2bca819e234725aec0655c1c0d75d3767fcd56fd41e5cde2ba09808e1c71f8bc78f2c6ea74cd03ec9fdda1475c765d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h346ed3165679ed6c3265a7ecce2600e1db7685f421b17ccb3f5c052c3765d48c608e296402473187fe38fc85706bc56b9cc1e421d1e82d986241d47d811f397b78a64db54c5ec0734d4dbf170d769a87af933c8997597d3942b0ea354591d99ab2ab012cf53a0a146f5833264571b6d32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h223bf05667b13aca38c2fe0bee94bd2d7ae439b9b655f102834030295940af7358232443d70e7e0ea5a1728a7132104ae618ed3f66b596c16fd144a79bd15cd69ac1289b15bae73b143297627f8fd0dde666a5bee795639923f87a2f4f433307c1157b9b7bbe0503ba41fdee5bd2146a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a9df957d29012179696ab383dfc526aa7a704b505f37fe2da401f98b11d14857140c0bdd2db06212c73f10cb157ba2d3c0073daa9ce82c461ce630663aade25a347bedd37b122c63d7614c156726092a6ee9cddf97c968f6d532ca5cff568f6c955e8593c34e06b75eddf17f047faad9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ac96b3e05de54db8ad34c829c97ead6fcedfbf6075424d09acdcb66216b70f61e8505c56d3d66ab7172322b43e325b463450494a64a262835732e86d39497c55fba2640f43dd9a33e4cffa751f5da2e78a35bd0b488756b9b3b3a6b262b04775d22114dcac56d878255b8b498cffa71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99695716c8efdafe825760d3fd04a46bd9faac7ee4d71bf7bffc942ce241fcca34564548363798b0c44944ea9c24125dd3a5019ce5ee40df9028e98e4dab849368e7cf226088a19370b69b2e83f056a13af776575a66e5eac0cfadd4891af2a17a784e1d477f7429b70b7604da8fb6874;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9f08a4cfacf7fa85180f78e34731d39c76693a45de1c1bf5296e98f993629f3e70185ddde58fcbc3efbbfcbcf8cba3bcbfe4731a65e35eaa7e55f87456c0e8c33c734fe82a9457c8fedbc66645a69557d654301b8eef9c29f93dbd353c93ff89d3bc148b65ebe9e8a653c85edeca5750;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0a47143f4e83dfdadc45671e2bcebfbaef7b41fd9bf181eb79fd78829b11e771b1ca027af740c86fb75bc904cc91fc111402d45687c012ad0d9d47d236dd874df1def4ac7fdf97508983dcb10e633e78ffe1bec800dff628fa218905422ea66ee9afa7032dff17b2dc9a3ec18c63e381;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h753c7f0e59f51a716cc4a0ae38dafdc0638d19fd7c93a0a447eebf841936c8b7b902bdae0c7888906c4ab2a45ff245334da80fc89c6d180d9dc93c7d42a4dbc8586f5684797242af0a3892298c63908d74b26b9d8a99905084f2d83039b6d39b31414b5312a7818cb8974004d28b80368;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde0754a5063ddc09829fe9fc5753f771845ff1e127643d523afbb22b3280b5b8fb7cf4e4892a2df77085405033b83fddf6991240ab3391c0c1c6883196d3f133d72a9663f765220e02cbdd4c7f2c860249c391abcf88c3d6a07357c2391ddad3112991be50f83960e1c7015b6a568d3b2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5df4ff793e2f44415d1c25bc78a779ab66b0d9a8788b358eef82e8e000ffc2e8b8aa81de384d6dc30344a7d92f5b424e73f8235657e2dc466aa7daae64890fe9019402c6fdf6c65cec3aad31b35d37a19d1d62b5cdab86b1154425e22a957a5e00c784c0064f1eb6e814366314bedaacd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfff59a1370bc220c7f7ae450283f9a97ba7f3aa10baccaa48c80ffea9e54e01f716f88f3d195adc0daa37b73240d5765fbb1a5da12d2b4e015bcdbeab74147ee123148939c7da0b7c272357c37502ec0f1ae71d15e5d522acf3277b45e6be9c523bd9c2381d3ed98da05f509008bd0979;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a5fb53ea0e0c9487c30fe48c21c84b8cb453a819fe0a4a8cc0841d02709fb20cd3a34fb245b82e09e8f0287d7879f9531583be0e961425754ea4603ff1410b4cb3a64c7ecd26d011c215d71d69d4b69ef542e0f7c6407964d4fe8e90e309373ce01ed70ee344b5985c7086636d1a1c96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac547208fd6a41380e0b96512d1249e5c32d7391b564c14479fd911b3e53c828422e8a6af1462b483ee49c7d0c5a5de2a0dde413159edf4ba203f1d447de0cf150f314ea40469d23a886ae7edf539eda2f65ccdfb07d8388363bc17ea0d044bc32cedc1e483e6011ccae636fbbe166397;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9b98cd1f8378ff8a1e87154e162dc97d9e9639ad3aa75613b84cdd30b392cd2d3e99b73ff5d88c4069f1ad71489ef377947fb24901e616d072ad10c64e9c068c1d081e25ff63573a110e305aa2cb56b77c96ea0fc9b47c67808795a4aa2a50ac88cf059405751193e61ececfc493cd05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15c7fbc02405bdac9c10643725d0c7864d2fba1a64cfd1c15406f646041c307c9a204cbe0bf6eeffe92ea92e90ccc228988563e9d841ad6ef216ec90601203ec3be42ee93733eeee709471135ba9883aee30c4e1ca41569c11cd4f5182570a2dfa368c3c08bd9078a539e735a9dd01438;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75c80085679dfedb7e1b51edb0cec19590c15d178d4e2bbec1efadaddc9290cdfd4c2e198988ec57e2847f3777007f12240d3c51a109a3861ae3dda892f33cc16c74edae31ba3bd9079f7632281efecebe41d7eb9710c35e745ab240e08c2758c67c32c1fcb7d897a7417754dd8c7d07d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff86d857a17bfa29ea4e9af4417d3f3cb828c8bf104f05f5a3a440a57c63b32489fddaa7f9447def9322c7c14787f089981072ed6cb53f8bfa39651b00732cf0d7a0d962117bcbaed3fcfbd338130c5c006f427d035ce566524dc93c28507d351a638ee9eb84cbee7f9d4ba4357ffd5f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27b249712cd175bc9db6a3c24917654ab079229b727af88416b986964d9fb9bf3bf37af9fa379409bae83c5eb872624dbcad8c29c4beb418084e58ab9b4b295112e51d6720de0d192f0474253b7abec25b6c97ffc74e1a7c65fb7af7ff4e8d50713cb1db41aa114fb8aaa0951d81b1342;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5291bade68388c92160caa3d6fc5b1985bd64e096c17f2ba9e822d3fb320b4ab7e80453951a495e5e5b98158b6615d811978d8633382c631ce927e6a24d1370188de0333fc7505c8ae4a5c90049debc52bdfdce5010830af468a0a0c96c31e80ed816b0e6efcfe22bca62efbd6c89461;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fdecdaabcc91bb6f2d298be0658a95666dcdce52ec962d559ae0000587368db0cb0ddf4ae2de03491e415b7f5faa0d65ff5bb169d150061e0b809507e413148ba52700d856cb5407ff33b8b4de8132f82c88c0a5aa4b4eff4fc3d5f4f1e05483e70c97017839fcb9916af6e973855811;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdebaa5e923ff1cc0217ba74b963b2945718b5745d1bca4aa59d8152d2d0b00429c293dcb5af4390dc17b25ef341d15578fe18e5ed775701c5e998654e4ad29cf07e28230fae4566e2a9a64ca8128de1657d080b7d74acbdfbe94585c588674e3e1faef95e6d7391cf3db69df4af44697a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26bd965b4dd2d83a03bbb24c10853d71e567429c4702e91ef0e97df565706ab8c42bb069a41723cceec864a243355e3ac9bdf4c92cc7d448d1398684f1946a519650916d20d29fdcee062371d2b75029bf26effa1e0499ba53855232a17df47d1b6248a35dca95c046bf422e58f0aca2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e5b0ff8632d5904c3f83c38518cb48df2727cf67b25fe449a81da46ccfd980ca65edd1bad9dd22d6fcb6dd2ebdb02d225c58e2de368088ce657be5e751484115daca5f1e1904cab9ea4d42a447a5d88379c855e122916a5134c070e2678f9662911b7ecd164be321e0477b292615766e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heebeb7b3992fa19319c61c0f239881571029f873f3d18bb5bcda98a7fb83782f3d2e8b2f92cf3a9da1ce94143fefcaf9018fed4a1683a857aceace01eed1133a74c012855c5d1f1032d7a6bba07fdf2245d7c575d49359afc9430e19d331bef199477fb023fd5491f8f22841097025649;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16724e2074a2a828810514b5fbab5b57e9cba1d50856cd7696f6482dba32ad348c2c725d30f16a6c21910b1af0d8237a4d98f056be7019d739d924b1e46ffb655eb5a45702dba41b2f60efa689fcea29610670a80096e2f8fd6145852d2735f186e933e3076c1b349a15fac2fa608dd74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb03bd4b6ef9a4c0b4c99d4a16c5a0c75077b6d59645e58434318dfa6a9264ccd5f241baf03129501d666191ae9a0fd682a7d8ef867029a17b396310198eecbc71f7f690fa619f477072c9905058a4f1352bc60581150db53970e2204cf0db00701190a1e8e67ccfb3aa4720f89330e76b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88bdf4e89425d1c074c037ba97b2b20746cdc482d38e589750799161fa451a6f5e3e973d3dda84dfa1e3094191892ca4b2f2f3de7fbb778eac5777109e379f9d57793042bcbce8bff300e86c6ec1ce985f668925a5209ecef40f59f09129b26168188021e29acef5a4bd40415ab379802;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h611a4da1497e1dd7092db8d38a5d3ea7c33c9fc5593286e23a280d54c52e96e47c9b85174d67683f4754a364310fff59d6a0e7d750c43d5d091bc4f3fa983ed321f7649a82e01337ea70d5bafc22d88910ddc922e3f0943874ac17d46606dac7ddaf8e366070432d7f4a0ba3fbeef15ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b2baf63317e6b11f877cb4072cd7c6f9d41da07a4379b99619fb1f54e5a93721926856fc56e488c0978c79b36c92753ff104a00271da5d998929e0381b4696f3bede0f2101f85dc9e6e33bf4f18b94fc33f574c38199cc8c17e37b64e6aa1b649d0325964fc2536a064ae22269f07dbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heac199cb9d209c0e0f8e53191f077c7690100a58f175886613b457d9ba6087c816322fa982f259f2b3528978deafac73c686c375640dc8411e0cc69559f871c7297ea002423e670b6e2b76d75f27b3f998b7f0f2136b86b9027642d175e9f65b03ad803d285b212e392f68f5d1b88bc97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27705eb68ea9aaf0622c2b896251f42eba7fcd51262120cc37175b4ae283db5b9b61711210900591aae8f267e0a6f1f0909cf08fec5583b37ff26b420224f9283c0fd2b7bbf26d2b89aef8765967f6ba53a0b715d423f8785ee9c796d9b9f71f4b663ae8ec2b47db2c10b7905ae133fbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc62f8dd9bd5ce41ae964bea76dacbaf520b08319d75fdd013fc86a8d1fb128a2bfa088bfc27b605506b42c5c5246924f08a5a8f267b075cfbfb47d10f889cebec115b6c3dd586d2528206a7259fecb1d0b9eb6ed0c5c8692a2b1760945836e4f577129dee759600089fd33928de17d44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h289d74eefcbc1df8697fb72d241c1d219ae3eae0be04fcb708cae21fcf04866d56987636ad70b6ad801934a43ea70c53fb3bc6990ff98ae1de036f7d9f98cb263123ff05046669e58963817a56076e17e28da49d810242395b3ba776d31c15f994fb44214a16894ec2d091725998501f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2662e0134d5e8720c1f03004266fb0190e9ee4bb1c5d4cc972bd1c73b225cc557e39f29043609da5ceb892d0ca10e636fa155c742ebe654397c4875700c927483181140812d5a532aef21041f1e7397c7b645661f4ef7eb668a963fb3a1d50b6a2135148028788e01accc1833549a0f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65888b614bc78ccba7bf5ffd68c048f96f65a99ae8e2efd489b93b38fa99889f4a5ee4d2f7adae9b061b0e31714235c928c284edcafcdfbdf05771829c3501935f401efbc6af33514dd6b0da179153406708a90834f288cc4dd6677f93bf4a474fd3dbadce8c7006ed20014e9b09f75a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf3f1ff0a60feea9c79248cbed7937bb683395c6f015bcd0de10f2eef7c55199016f5f873c9f9cf18d579039a0e1b604998a192eb9bc188e68c246ca75b153e706bf9586bf4bfbcd7bec24c98f462c474c969024d0d16a1cb76e20b36a9ebf845c6df977efb7bde7d2f38fd13b026220c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dd011f423d89ac8c822fe15430aa4efbf359dac695032d2ce6194cb4e06e22798e33b355404e39978af2fd598498f532b02d9b9fd18392404b23f949566d340d73bbd2b15250bc6378333e4f0fb984e5c9d4603940cd9ab4a10f6f714a1475878d13182cf6568aaa26b3720226fe8e9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32dc6e3f98a097a7e2a3dbfd8ac7ecb72905feb5b956309d4ceaa16e9fe3f0df2458692cfcc9ea4828a030dc19e99bc55a5c1fedd512e38b86305c68d1133980aa619d8f614507bba8f6e31f120ba8f54ead8d96ac68b2f75b74acec45d7fdc841d93f1dfa900544c6ab0aa113ff3dd30;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1166c2f32daf6b8d1085fa926862099b44a900a13df9347af370ca92393b6a9510cb476c36c1aed9505dce7205e17509114ab932fc948fcbdd479db27ea83bcff23e51171000282867f20ac31ef0b1242c1f17e1ccd5abde13f660f355dddb0a2aaea05b151d1d263a2031ecfe1a50d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0b448d589c6b270cdb18825b23892e3c2bd80b76a316e6f71c24c946fda33afdfd036e205ef97de55723c67f8bc06857dae7c33e29829aadd0be34d5d749a8a9959c31a9ca85ef3fbaab32632689fe4881d14f2e5511806d0d9d1d2fd1ab4fdfd590d540f6740100dbb4cb942bf48e65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h610fad31320d52520e9dd06c81b8413706c19c39bfd1be68b2b2c18ba06a90e80996b2b8cad6238e63fe06636d21c4578ddc730cb0ae3d181de62b197dd07badaaffdf6e6e904eddb9c4df5feb209e3d92954c3be82f8e9176f1b130f25b35c22f03ad871b070dad1f372260a0d72df5c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39ee9fb8701128ca7f504e3c7f4396b34ac7efe5593a5e666a1e3b42cbdf09ad799339699c6c253f4cb07b75116a4e403c6fc55c673153d0426ac69e3c9ac1623a29ca9800e6c8d99d1990c1f2d60a1f2765c0eda047275c3955509e3bbee8c9362d03a76f87b3396f13e6a6c54ed59c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7f49811c5cc30756f56c35b5276fa23885e7c089f2603c854e8201423530be330585bc60bbbbf69bffdef0025e38e1cd9e301949ff9531819a7192e9a998edc219b965dddfaac19dd6999a6a3678f641bcacf7c56f4d1e82b9faf378abb15888703151fc884bac9ae2bd9fde6a47d2bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4f0ce10df20f9357947e37c9a045bb2941b571443b20195a002b389bdc3d6a3bead2917f9fee128df41772bd500c44df20ecdb13632c8d1f3f1f73564b3bd74b0af3b7622da5c9f68c8873ca2c2089317f572f124a97304201043f0760c0f82d9ca2fc5ca1f4ab6aeb2bd4cefe754f77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f481a18cb9cfc2ca59274de293c6bcbba36bd40682264cc28a68ff992d498a008e7c38a062d09a6c50b417f911dd3e582d6ef41f4ee5dcc81c5dbef1f6b1a99f4b5ff34b0c14c15d064248290eaff5da00861c2bce2633ec2bd2ebc935a2cde4414dd9fdd2d3d73d197ba46650998058;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21eecf4c37ef95e86b6a46a9d31b96a0f1c66a49680bfcb8dc947ae2bc15e5703a970da3c0760bc4d0c9ed89b57735a596d23bee3102ec49f0880bb7c4a43a6bae000029507df8f92caea4894c72cfa1cde4d1c46bc4343e1cd15a7e2ad65d767b5a42adcf604126b938a95a49db1203c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h201e83c2fb8c027b2171baa46b88dfe0c8ff7babd5795dc58d7c2e02f16199781ecb64983ae09028c28ca0810c5b5e2cd35db1e668648da08ae9462a4292ed240b099d55e156ef97791cf837038b2e531bcf6a19df83ad815d863581af86cf401c26b757a70ea0e0aee858733b22e4356;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7114007f70371c2073debd948101ba59d033b88cf7dd7472acf652a3f2fad494fd8ce933ca7af8f40fe5f6aef94966f677f434fac334f0e50e8954a503bb694ace0ad10dd987ed897c105d49bfb4d240647154eff8629309d6d5e3612ef30243b245cac8c30faab7201c034f3bb8c205f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e3eb032a7b75fb1ca110e6fd61a0cd73b19abc2e17ad09c48a7ef205749d9bf003c44f5d9b5a49ceafc2a5f4b543668ca825588e742af0121416d7ebe6b7c144b00405b7de77507b11d44c36a40cdbc3b4c8e53451005e85a3eb7b3d03fc1ed31f75091d22146048bb9c79823ea1f5d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb983e07ece6dc96077108d5d8f1fea2c890834d70308ea5fb13cd19d37309ce21e256b37521f46766c792163cabbb0a10591192caabaecfac1190d6226942142045063ca3c92e544cf3cd9c0ff41063d4f5a6b09301ab43adc350e7fad61db943d82b14b847bd179a5aee5b56d89062e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h969313e28c1f4f18cc3f42ef0c0fa701aa6eee0918930e9aa7cefb8f4a5c9d63a068ecd90302d9a92741fedc4f417dfbd6fcb8fae528fec10dea7ee705d88fbbbbd5a30d4ca3e680f63ec7058ade80b36b8efb235cca3ea13cb552ebdff2d52492f9eeee0bd2e47071f30f0960ae703a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7696ddb90369124f09ff24f5b4c54fb853e273ab6621aa2e007c232eb1a9ccb59dd275ebbf0b94b50aa329adfb7bd0b2adf5194eb43c8a84d2bbbec0b5eee0f02ebb9fccf0647f1102e5d89c564b9870b292a058fdec23aeb579f520a352325a00864076b65cd3fc4a8c728818997af8f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda18204bacbe917fa74ba08d07565d9971637156b3b6da2d8b51fbd2a5e5d93de24c1a4efe656983dce41f040c97a6891a3dd31fd87c719b775a09f7b614bb3115b881457f9b546f26c71102b33ff71f3fdf947ed37bf17ac632a7fde9889871d92e01114e22deb1ce3349e75e0bf7c5a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb2b1161898c84012efcb56aecdb0f427f77b808cd66ac0af321a51148b5292efbd5fb99b1e166e70b86fb706d999c30bf89cf457c80b860ac0044fde6c463e1f3f5909ab64980e3793408f1f5f14f9c4c5c357ef2313c51714a77972a818acd8c15c0ad824aa14fe48d034ccc9470a22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha13ae116344f3c08f6d9441c7b5eb2e8e5383b1cb8f104a9335ae5cd9f2a1aee9f416bb078de78a3b930abf45a3d22862cb5429b312e9237f20e3e2df4458e3ed87f9392316372976844369b733f64f59ed73407ff3cdcb03defacef4c09d7a98aca9c3d6ee4d7048869d2a608d819db3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h493a75ebc521002b742146ffe865c8b24a3aa5cc98b87f0b6fb33d9b959958c9edc6cdf962442e53028bd8fec6cc6889f191e2c9dbc13d2c4218abd67ff8dea2428a6db1edf14600c6c8784faf1f0510368c851f696d6fc2af09a83e5346dcb066e9093c3d5793e4c283add51425079fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69db9df96798aac4843941c3be3a3754e6bbd831e17df6b45f51825eae5ededf5d776b7ed53128ddaa8e7167307b40f2fa489319619e5f6d222d87365e8f07de9e626d43ee5b14da01d499f076adb591d86ed6a89058288d685f4f55d6a60c413965b4483d1a9ad284ddc2cccc390acf0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7cb3c34c5883eba32279309ec2deffcd484f7c67658ec95c73fd196227dbe70a5f4f49586d34e5b488fd84d5d7bbafd4a882725ea8629c0c7e8b488319348d265f69328f59c7ff331100b8b6a1801a709a4746a21b0eac2851537ce11576b3aa65e7dbda56dd82bcfff5c814cab40477;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef259088dac1b67019125e2cd28429ff81905f1135ea0e42499656f6bb48506b978fb21d532eccc7acbe13fa6adafd5d0a362fd94781c36df4a6480fe7af8ed34c268d8bf73bdb1d8a0dbdd6da1258fb845352d9390373394d6924c95eb9185bc67905f7f4a62497ca894d98a55835d4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cdd0ffd3500c53d4fed79d1f875c3fa96334ca1375581810e28d5309b2faf498d00080752acbce14568da60467c898119dbd4fe776212c6dbcd235e486d74ac7c52d080825137cb860aa61d6fc861088a8cd4599b8b4e44d6d9a847e6a54e74bdd416f7e8ebb5853e9c72b0393ab47b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a489c5dfbc01704c1f09dda6b590b301e7630a5fb73722eae334eaa78abad86f2419593edef5f9742c10278969b64fce164c7e265afd03d51944d6f8b8b18f3c27c727d7001f2a63ac2c4fad64ff86ac614b13215370d9510dd92aa1cbd799e7e5c4a14febc152376d84723f8b579682;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a1a3de7333a22724977dda6a1ab92247f7722b2530843353ad4990b30c1f192ab353ae38a9ac7101f549be9383807d3cd2501664c2700c99b4f5b9d203e61122a04f916faa1c051d27222a0f7e10880c9d49fc110bb716984fb57ff777435bc1d7b1bced98a7f524aab72e283ca3f98d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34dc82d9dc3316a29fcb55de2f2d6f06eab96cc2898a1694e94d92b6374bc057cced58d7484098c8122e53b9e5e3ac0af42482f0a09ed4565c947c7be89de0dc408ccfb419e5550ef5aefed846611ef5987abf1e828c1c62a02ab5ff9d0f44249f89ea102d8119f32ec791020763ea8bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24525618a746e1337dc5819ee6adc7e12f8c2821853a30459d4f2f55b156ca1fa0ddd998b037e58c62787299e45f28252139f94bafa220def6f656198deeb6d2a88079aea34c1da1e6f8e74b2930c50a2673bd379317c768882447b708ac6d00da36fa3a0dcd44296e3f983b2d642840;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc6d53f6705364af83c78cb9028866239b262ffc43283e84f0210b938484a33a7bd7097a84575526c707d167de5155cdb7b5c32930a86556f6da5904bc171e1654f0ac3805c123c6473ad4bb7e7f506814ace40dd12a5e54a23d5d59f6a679e2d6996e96168b0faa4ae7e1bb21ba0279b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd41350b6554876abe36ca5701cc1ae61d97cfb2487f9a704c5e16fcbc160ae1f2503db78e35db99d5da199d5033344b2bbf37901d9ba49a521d1ece2b6c88c40dfaf11935c0413fe60b6b17265e6ff57bfda35003abfc33ade45df032a1d23e09495ae96db9a93d9fbbcb34d7326bf26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8dec1775ba6aa936d3c1ef6e48721950f3420e1674398ba72dbfcec44c71a333c4137d019138bfd4637d2ef24153102f4512cb6857a147dea49e1dfe8046d19c26359fb9bdbfd1d8fc142c4502ddb97cb036b7b89a58a49d3b5c2bfe76ad81ddac98c455cf8f2cb82ba870b84d50052;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a141d7d8fc2dd43bde6fea4419e72ce736731d986b6df5b446db78535b9b2334b63d5a1ba7863abc2902292ddc9c5c63f4d0a2036784daffd89af7323fd13f8482f5e3004cf753cba00b653dd8277db6080e6e7ef74bf3b37d78ea6d3e2961e0191745022465c0c09b29cd8b1ad200c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99b6ead51a1ec7ae1e7276d57d3a31512214284a29bbb8ad213cf866e13401614faa22090e07558e0059d3392c43d40afe778bd2e59642e9032b3fd5739042353b3c8203128cb22ecaa88d6452f0c2c0008cbb8143596fcbc7a7e5c2d669a6b6acdff035f2726c96a84d0c420a617be72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f2b08517b9c6390fc96e4a4138620a9ffd9beca87635016fdc4bdbfe397d6b168b078249cf6f7c8afc366eb052f65f3c658655209a9324fc49ed0d13498d37b94aa818950af33d2c813191ffc9c09142b245379b2f19af5838f77622c163b2479bf62e0a602d8425d4692de28cfd7889;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1826de5b1b41edb364e7b2f236876ae111cfb2672d8a9ff07855f89507995ef9840d10ab7a798e5854df8ed96bd9006c2df0834789dc92c2585634bf527613a33c3f4e8d0d16673c1d732502c924ef724de9929eba4b3a98a07bcb3fa28a6332d1a5d4c882359a44ceaf3b32c5c052e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6e08664b1482ff44672f69c8d5942d555440342fdd5b20ddd70a72cbd8dd6a63a27953de0f1ba5002a07d4ee24f6d7ae2943aa2cbb0fd40c6406b56b08927ba6cbb179eab691af6ce87be9a32ccb95362b84e8e4071c8037283f82434380e7dfe336cd8757c09e693cfe90d7bbc2e135;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he24b3f6f6867231ad39fe511fb65c94a8151d541db55e2e248bf4004617ba9d8a3bc76f98fc964c66f5b0faa4cdcca0d4a7acab0ccd88233133d423869edb7a354112a26d5bbc3ea7d51d53b91c47181ac579ae61dba2570e6f2b7ea049023741458674ab53f23ee0809e7474e94619e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc2b0208eb3e6bcedd2ad40885f658ab48247510d703e68a4efc5140f803a825c3aa97c594631d9f0c4a69d4167c42aae4388cfa6f94f7fa5f295209fd5d2b2beb973b8277eb34f2b1eb6d8a957a07c437c2759cf362db78d5a7a535a5db19529359ca82a58f57698bb2a1b617c787305;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb2698bf55dce27bb212a1b635a5bbf5b6ca31dcebec5be73824f051b799dc1763871625244e6e331631a8dc7b50e2520382ffb10d38130ab0a6fdec79ae05057716249531e2fe000753f715d009e66e54ed34704e126dd12a65c4d72f85fab49beb106466f747bb5a83243abd393431c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafcf456b16d87ae081b41fc8d6e8892992cd5097770856da297870e89f512cd5982b9d7596d3378d9be3dcdf5e9bf58054c86443d0801ac05be207f33531c339c7524af912d8f26aec8a21c944995afec8be3e769bc038bb07c9eefff1c89c074635f16ccab2eb1109587b707f69663c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc960cc96198eb291343463c420b4fdbfda65af73b69aa677e7f9a3a838999745fcefa65286ae6bf89997de597690ac20a6e66996fcafcbaa5515a2e53a9deae13e136e58d3263bc837de2644fd7448fc0974c5ff8ac09ce4a043e759b3cf70de809b8a084cafbf29a666b1a0883f073a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf91f2c551b7461716f1a0bf8c2d417b38f96c9acc137b062e97ad752fc3d7f555fd1a8f0a4b291bcfd226128e366aa09e7e001e372195185e44a34625f8171a5c565b7f13634f604a8c85ac7b746f404f254c8ecd20265194d39780500255f4d5ac87457b93eee9a4025802715937947;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62ef62df27ee3b22dafa9820abe1bc0f064682d897911d48f38fd33bcec5bf45536a97d78abc4a8468b62ca514d18cefb8c475a4f32ff42d0c0a05703c8e2c4de8483b1ee715a5d0fb8b0147bac88f0756f507362ae060df1ad2be5e94cb06a91ea8402f6c52dda5f6199fbe3f8aeada7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b05aad5e423a20bbb7a7d1ff6556f2aaaaea66e4b0c9a1fdf66be63044d26cb676fb9810135a3b759200b30b836a8dcd44ff2282046c978fbe50b3b2cd7960824bfce2774ed0bc8bdf88f200780a24f58c872b5f7f4adb96620e20d6c211b2492b7a3ae9f1f60a411d747905b94abfd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb23b36ed9f04d5e9796759468666174d8a1a0e23710ef28453010bb994afedc855ddb3cc6d3c0767c0b9330007ad7b4b0ae7d75c1bf47091b4e29171501eee8be7588f7226cbc7b5d8ef60a320d6678cb3bffe278c7760e6eb38c33dd56b71255c7628d0f5d3e28ac365f50b935b6f16d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9015c29b96d6c2807d0193a3dd58d0be0bd0907bc89d4dcdd3a48a09ddb999904ec14b5dafe6b7e7e0fa3fc71c45b09130149a9e7b16adaa02a11199bffbbc2e4a5ef4edae347db0daa09e183cdc7f08895ad0bed1ded51030aa6d45647650bef8fcc23146273b9c36871c2d0029efc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd832c1a241b1bee9323199105a57c40b653530b626bff9686cd2d8722e671e88ae95a4ac2636d55132db96a59dc8b29fe1d52eadd9bda7cd5f38f0e2d7090ba6bb4750d6260b6ca2d937d3f6419137f3dbbbc610617db62250d61e5346ef8cc85d8f5de576e73373237c9db2a30334f64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h561fabbd52a8ebdf68b85f02e846196b9d21ccc307ad1c2a4a908c8e56d17e2ca23ff2f96afac02b4465cbb9d609cf4a7774fbf343ba3874ea9cfd04dc5910f691ca857b69f5dc5ba02b3c2cedcd5eeb1ce12b7a7b9ae207192e2492021fe1c424f1892ad8c781de0d046379ff00a4e83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bc51a1134f69cbe70ed2d9f1a9096aafe4590f5ced902727d2b7ee2e9e0e1259785e1b5496e6b6a385ad7c8c8b8b0f6f094706b2ebbe37e5bded82af26c35ad4ec7557db1c8733f7a4acb21517dd1f837d30f7e6a6192fc55723efbb0896d5d20343ec2d27b0b7adacab66d312b0d278;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54298672d78f7259eb39edddcf85d6cc9fdb81a62d5a03d1836273a5aa22c3e95749fa666bb64eac5c729a86e2154cb28e9943cc4fa9566a0b3e3a6cd28fbe06b9f02b44fc801670df626a3bb043134da259fa6d9a0d4ae19ab4923be36b1523aa45837796a3ae092582dc4833be769e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf68ddfcedf4a600ff6a8d33d4135ef49c2523254de83873d4588f5be6e9579741ee1948399fda646bdc5ef7a3f254529cf8b55826921234dc3ead6c18b116e8d9aa2c27343f4d9ae0671cbab8dbd754089305d58d386f5289fb4ae00692a5f31147ee8a638d45ad241bc16e9bc310a9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d374912b7b3d9215045fbabcebf15a92d5b0a1f0a27b59bc56e18e2cdf138516a728d906216aa1c77511e7b91deb7f77a15329f1ce92554214e7c632b55756701e628a4ec62f1edcecd7a93e3b8e6f0e40e3ca5b57c1ed2b3cea0d498d8d321e1919cd36e1daa78303091dac32cf38c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23612e15f5bb49f523b546809687487797fff3160444cbe6b8b3f552834ea6a7150deb7f5195143824c93fe838f6a1d5b2685ea532c2ffa95ddc0e21d7b923461c878a923c4578ed5aa918b5f5c7aa9c8d6abf3a68a7e6afe42ee7ad1a3ba4cb7c0f11d324770784219a9a1c54434121b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha84bf6efbd611752c1e6b08642c54973ebbb7c092b15a0e50311a14e7ebee421ade2cbd654f1064ed0283a05f89e4c4a1c9c7e2e214ab5c87aeed65e898cd01f0ee9215c6dc40942c7ba59bd185b584d553b46678f66c842d54c35fa69bc36fd1205dae97b4cc42783782a03da25bdd6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd83aa949fa4f8d9ee32eff10ca6ad9187f5737cc8bf29ad786f44eb587c33785fbdd617113677b862f177766212af17d395312614b4609fbf2a0d6981f41627474fe5329ed8bb18b194d56e5268f6e40f4b6ce2296e0c434dd2abd671abfd6a768fa3317853a2d0dfa77c51d644baa60e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h478965b495162c95ea40e18c3e7ee59654f4321a47fffe2be6926a8401d544d22fe77091850bb712b28dcf9b1aebe5b2e6b63531bcce1cd6a17cb46a5ea361b72fb8790afb3647eb03d8f78334615903a6e7729eea209b05d1b8545cc524acc6df077519d2278ae72d6e6f2ca6eacbb93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0eb32ff94cd0c957bd3c0e17ebd545f3ba633604c07df3cb91359366933e78282a4a01ef96c7e17bd72c5c6697f8af27931abb3020da2991013dc8b092f2d0c4f33e6f1bee2f2895fc30fec8d3960aac632af160e78def158481f9e2850848ff759b4d1efa5d5d2954a98d33c6a67735;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccda31da0afc5e34f35b3509e842735e2c2c9ae2c2efbdc59b5f7ebeb83ff86a6b674853609c39f4f69e366e322deb112455232af4fea075df66c4e480b530c7e4830f54dfbd97c0e5095b864f032965c770da1062fd81a00984e1071aaebf57ce48f05f8a78c56e2d2069be107d15e6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb980a493cd00c479a6d13ceb2e751e7f4403909b48642081bef6cbadffe2c9d12500cddb4c8f965b255780e39a0bb8531ed92b9b91d6ee316958e5cec02a7315ae735dd640f859c360e20914b93aae47ac708b7d41878b11d3e3f04121f2801a7db82ba78c294a86ebea541d031f0e6c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2ad56a24a72f78b1e2c648e3f0af55bc8ea1e196a4b352e7cbc84752fc6f2ee72193bf9d0bad9143b5dcd43f2eb95a7f5a0ebdee74f135c03c3e3a1d9f18356e07695e124ca64dcb82999dee10e09f410fbb3ae759c18a8d3d7c12ce66c57595b68ea1ad73a550911b02ccc8676bca08;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb77f02a35fe9444ec514fcd0769f6cd201db5b3c75dc9c12bf911519643a68781cced8069e6302041573e1d4d7e0fc533d22efe90cdd9bac7b5402d9965815c832e1266e9e6d8106e04032777a37a754b124a8411cb647c54032f71aab7edc6c7ce5792d8b5da69a18e75a77a3798042;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47666614395dddc0c008f04a1a3581ee2ffd6462161741ed5c70042e196ad18f067f0fa2510753d104b6f57a132069f3feb749a3a263893c980bc7f2caaf5de86c3f2a66ea5b678d75f2a40e9fe6bd27c5aff267388319c84a1fcbb480a59c4fb55f3ac72bfd162592ee137be8d5babf9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3755fef3ccc6958c36d136bca1520c2a1c44fe80fe121d397647e73d122ad2c7058e4498491e8a17f96705a01cd6cc7ba0f499596aba610ca31682f003ad401eb758d804d904a44085555ccf7dc7a221d86f88823a7da10e42aa623a7be65cc5e6f67c23a2c828b2ed3d651afdfe7579;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde9216d2250219292300fdf2c48527a913e6a327d013bdf02764f173b708861dc2289ef55b8ace6d4888c7916e4b868e58b30f0d18b39ec7348ef1e7a9fbbc3af3527e3d199ee8ccb6d1cbd65de05f5326624ab30e2bca52201a7348cb4e530f420bfb23d1ba52dad0efd979c4b513d65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf28cdabfd73550c03b0c407198ddba599a1db3544dfdd7733130a25229cad143f210a4bb54998b3eb112481cbd5f33788af6d524a9b0f0abed2c314b1848f53b84c1c297ba36e935f8fdaa95360df84153545826066b1c1d3bdee604fca19a5e285b4dde6bfe3e83f9903b91a2736e06f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h615e9939e2fff93ce225015149a8bc51ca1ffb7fe9cde9e7ca1ee5bf5258f8131b0331bbdac2051a4b2c87d873f0b640bf69f6d5f26471eea86bbcadca7139f7000bae83a8f16d9ebcfc3db6259dfed93a1483e067ab1dbbd88ad279d2ba55673d687de382a14a8dfeee9b557a6b98a0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95fbfe65c2e0da6c301d72d00c33546aa6910e1fb44890fad9c647714d4b6d7731184122cca2a03bb165a947cb96c82fc11d33a7ca2834185cb0ca9a38c4adb4d352ddc38f1aaaadb5080249e6bfe6ab94680610b2f528350241d414d7839159b4da6033fde1e2de12146c4f031f50ae3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f3697831c6278cd2f7ac741881f654a35be47b10f7691221c74a7483458155b2aa578814833d5d2598ad4a777e75fff7b46e8821d5e13fc9b2b9a47d82d71bb03035675f58e01ddf963ee81257b25f4c40dbd1467dd105d803b035a620011c2ca399210404ac36c9edcf844e56886a2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h112dacc3bbcdcbe40c95f4a8aa3043363509ff9ce005a6c42a13a0390647166c53042882d68be99d35576924c2a05c31cdde5784642a51b65a71e8d39aea59a8ca27f2986f2efb7aa7a76a9cc3f86bde55934dd2f4ff57bf6998af83e4d049b02d15e1e691685b5658ce2e3bc5d53f475;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he63db9a3315cd6184eee80179ffefbb04ce795f72d898af6d5b99bf4e18e20bc65a7ecaffd0efc213e60ec791ca1dc54f0266944dd50bc21d840a0919231ba5d8b15dd1c21bf269268e46acad278dd7f76578f4285a204cab04233d7bc0161a92cdba4d57506eab304b37968be7507676;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h738754042f835d076a04fee1f1b4417bee907f03b9d38551f00b864db00b7ce93221ba1b0188e26b07ee5343c7fb50316c2230897bd4a858ab6c66deb8f38e9c77cbe4ae88f196bf8a491369617ddec930ffe3078f0fc472f6d9675cc8928868ae3a2322c2fb0b628972b83969ff4eb57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h437d19b1b5144565c8f38f000a5d521438bca853535cdf82728e403863face2b6d3a0296a85cbf1de4fb0d7ad7f1c24469660e87afd2dae9f0618f9e2293f80fd62f6d11dffbf0160cbc4e48992951b5827ee0ac2ee1881ba3284b8573cdabf162a71c72395c5258923a50a2a8a94e96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb86ffc48dffbcd2b53dcdb73cf998ea61447eb91b416b09541a9df9f8c9c0b6be1f1a45136918d57f7899529e5cdda1008629daff0d6385de4da51b8245371b1227da87bb17fa90490fdd2ae504bf4bc1158e11df082b3b9b062a83fafe0607b47607fc44da77b64ed245d36780e3a3c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha61427d2f4d93757d69c7b53c57fb67cbfe4ff3a734ff78fb9fea653d0c46b928c95dcc37690a55258b118f0c7d67a69288bbadc4db92685b05fee34b4cbafb18084c6ec528fb4495d0b01f7262a72436a09033309eb16cb9d89af8f591ab4d31efe3d3b1448dd6865c88c780e62c1d73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf49aafd641c8a8a4231279834f0ce3a8cbbc00488de6994704b6f528aee01e0d1b2f746101187141cc7ddcfe70868766cb5441870d328d8406763a9138fa175f0da1050aca8dfd44f1bfd8a48a11869ed50adf4df602ced4aef9e5d34175e882dd280f98ccee73a08cece20bae23383fd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc865f5d91733198f8ba07647ce81760a0473f28448a7579c34bbde0b1df88b57d8d43c164989a4cfcae22208dee29797fad569c8badf6ddc253950b92fce06d4cfcef6bf9217e54fe899f87bf8dc511f65a2df99715f99df47d93d537d573e520e137166953988e245043347aa018ff4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1756b14ef1e7ddfb8ba483b2af12a6f3ba8715111af08e72ec3eabe5897835ada72c523e222a5042ea2fe316dd0734de9e4fa7495b42a3b72ed1fbea5700524170cf63d5260b610994cedcdef1e7820a69d2f0e8c838d09c5ecf30ac721b1166ff67ebde600d1a3803c00a59046f26b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9996001a57bbf5d66f00d943b11a98aab30acf1d1c832a3890c47c8c37f067f773061fd8ba7df471021f259e6eaeb8f232c4c29c0da2a129434b4b568de214432778c5b2fe32f327f8b79b86533bf4704dd782a5a72b22d5473b63c7e8b08b0baf1c68f28333d2c0003682961e5a89b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd39bb4e87cc2f7865799219bb933ef59fd964d8ed388250df3827cc813f5f97186bec20115e4b5334d2e034fff774abfddcbe164f2722e25ce45bf9180c62f7f44b9d56db9711ef7103ea2db2f97f2322fd81218734495cf050a1d726b49da470e8e73844e946f65b99af162fba67b242;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he56abf0b364152d7a9a49fe7af991a50ebe488eade95184e1acb46d2ec0ccf7cf797222f1ef749b68242bce25d80133fc517e11381da3f4557d0dcca3a9cf9fb761fe246972a9e22c82b7f344d2fcb0ed8d3a3cf5cd80643e445a4002e2ba7794ea465550f8ad373dc09579b4c861a515;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h385e2f09f616233e897131b0dc3744b45fb2511a7e016f295277d7c6dcbe41749e8193589157a75d0e41980c27b0a7bdf6c3ff0b19bba73094ff34176c8e196915151e792b43e44c1f09b28f70179bcffa7767f3443fddcf5eeb99ecb10d529474bcadc4b015ff6d365aac37115bab6cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h282df150a73aeb97ca0e7a4069556f4bfa9aac2c69c9bc576c172406b5bf15b212e94bd4535e51d0e21e76f1d12a0bcbc20b67d2067984189b45ecae799e1666789bdb44d05d46676ac5aec06f0091c7b485806070312acc73c34280a312bc6bfe76630d050d0a22c6ba16530b2194199;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h388284c4ede609fbaf9d1da13948b863efa6511ff2022a9a2dcfa7a99d7755bdd23e8112b89bf311b0396e5a9dacc96150568d7c0737138247ee2a9ac1802dbf60b22161d3bbd161e117159c8abcdca96bbd7afb50211dcdbc21f131eaf933bf267788627ea64727fc2319d43108f6f46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96ad80cc24180b7231db71abdf5ec1805d0e5292b3d7647f63494b410cc2192683a7f7fa8925b3280453b9b9908776bfc8af4236fdb5591e47b2e006361d0da307f0560cfa368201cd206cd4a308d85fca9f9a3dfb028acc868b04a9c2532ac950eaca1a49a5497ee721915754cfc3d41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb70ed49894ee651f21831ea894414ed8154586411d63fb02bddf385d264315d9bfa7dfcc88443353e48522e73c9959936ea7c8e02bde9cfd38a36f646b86f69a00285e3d072072f3c27453bd67af62be86e2b0bd32e7da9fb9915f9c66a6e4e0b3a80a149dd368d2d90932975c74222d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24fd0958943ff1b9ec5d0de68d7a85eb8d6bb2095b5e10de0011d302ffc136fdb672687f25a4adda3bfa304faaf6bf4592e03190d67dce5e4a5b1adb3d73332e7984e874fabe80a93b7b2b007530a39ec7c552dde1762fc767f00420765e82abe332f9fdf46c7d33db641ecd01e8aa83f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92df8dc17a70303131c5c4d28f4b506cbf0f7eb30566ccb277e47ac6d026e1d5589428a7d3874355c33bf57b7d86569deda2d1700dc96890d2d5c23779536d9defff5eda53d3a2a7dfffddcecac41388c3c7abe8fc59c0c1ca9887e91475dfb221ce9362064e445cc65a704df28e41f62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dc2abbb7cd9542d81772a53f015f105af601b8f248f32b502c3f9bf38b66bed7d5a6477d84db91dd504ac091dfaf164a04e077bdaacdb60af11e07198666bcbfb52aa5e53ad00b997aec3e4d2240e73ae809e21cbc3f1824517538d514d5a6d5f329e6bfdaccfe5b5aad6d8b5c5fdf8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fc1dfbec2371d97612d7319391b2abe6e186cf06271b0833704c6dadefb4d319bf711f46e295f3a172ba26a644ecb8dd63a57ebe7464419c6838e9a9281aaabd63fc892e8b2a50fc4e103834136463b4f1f10b766f53c579f1e561e8f8bd33ce1293931b6b91360307d34d3b0a047891;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf129a22be034c4fdf83c99a336f5159bd68aa5c23bdfe0871ae8866cbdfd5e55e130291c19544ffcacff4c2127fbc61a08f28c69b1338ea086e3fb2178db175b7117069fbd5b3b98d3342b06e2440aded5888c23a3e31b25b73baf6bd877ec9e777242ab2cf05185cc8b3982660f5e257;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63f59dddadbdb94529a4157e6c22bf3a37674ff19806670743263e184e354314cba5a3b7f6a9fc5a546925a20983bcc241c201e1ad77bba754f08e69091d0a7e2d80a64cd56f12e63b9566f39af98801267cf92a5b840138ef5945b855ffd7efb565a903b2973179b9962baeba26274b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c449c8bfcb3e2008f01336917b593fefc9cf76d5da5e2e17bad411e9f01f1e28c8394271f94afe4f445b5f023ec12429e98704430edad60de18a0846378705c45122b27dff812d9f041f5f97b40ef10b5636aeb0a9c9ec9a5a2962c1963ce13ec21532fe33755b157aa7a32af5af69e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf327d40af1f803dc3c63419ec9df7d85dd3005e8fca952f7cce17d751ba9a403d2b77d78bc8884a49af10668bd8998ccce550674d8b2d9a5d6f481e315741df611cf08f8657e613bf4d609f2c4c180ee3df570596a9008071bd34e91171cbbfbaf278d9142f363bd718fa777d8d7b2106;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb42b9f521f849468afac7ffa1f0c25ed97fd0e94ba3f645da076e0707c93b28132f880199684f8c3e4eda9305b41fd2277f39c7ad6929a3d2b8c7a34d980a149e459b9901b94531e8e51c4df7b60b4e1340f06a72a10d743ed183303183b04909c13fcf70d94de7a988b87349d9bca855;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc149d8c74141635a4799e6480cd8b0d3a2339ff3191edace66ea3f631ace1ba7616759270f18344397c19e22fbe0cad4c577f9c9be4c06045c1fa56e32e7ed19a28e077429f9ef0edaa5da4d25ab3b4fb9cbc92a414d05f4e43b44391b3e5fb750d65f89f2409afe5086439a300b82fd0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90dce3806636d37bde4932e329f5d7f7ac83da7e064fb5f241a783568bd906d0c7d99207399857b8a006f7c1f80a980dab25e4f8d569db00a4f36496483ffa0e1621172e9142aa1bdf6e8f836503c32dd6ab66734c533f0385123070a3499dcddad5ec1f69a0c58b234342f1255652daf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71c95d2ca8eb4a1016998197b4fa7f4382975264faef9aef43e3578a1c6052487fa6ebcb826c70b1e3d9717d4620fa16f84ae8bcd9db7a13eafe90809f066ba469b4864c677f3dbae1a828545b6f1e5d1031e9714af1fd820816d823f9ec0b7300cf883234a9272b87f1e35385a540b4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h932636c8ab205575bb066cc123eb3b4299630139a49362c2db009e56e2c47bec1449badeaaa1308484e7dc4dcb2c3554da6e8e633ca83f09d94e89aded08fbc6bc815556a0a6f30c661406f8ae0692d280289871ffde5b185c9081b09ba1f303b2d49726580359fc6d15802a1d476125b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27bb873a81a5ac4b32dadebd7a110c69834bb7bebaa7693135f1e9140f92550079bf2087f574821d962874cfe41273f3251251e40583f697f616caf2806c05fa9444964bf277cbf9f0dcfb711acdb29887b97b7051e053d94ca24f69a5982d1f3e0aa6749239812ed4e31df0d65e1a299;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90834df9edd895252fa57f1ebeacb1047231afea878e1af858e2a5f281efcf87a2e322699ba11531fc19791c8909f81abe533167d4d739c59b774ad46d0c4149a32d5247972a80a56de264b1bfb371fccbd0a7ec8b2391d63d52797a00a9164e1458837c43bbc4ff2e19b4f1ecbafef74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab0f9d5f5853728c357441ca97da203f2adc4feaa10934c04c32ba06e3289189e67acdf21fa38f9c10380bd4e628c178a42e94e48a430602d549ab89f7929652be9adb4f64eec21c8cf95910f5c3bd5531c10035904a506819f9784283109adc106f2e20d8283809353d9c7161936ef1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f4534a64605a4b3b132410c0074acebadcc9dfb52e3379ddac2f0cfc6f3796c472955e0c91ec834340bfc615b0e00bf8947100efc45c3e79bc46f612623cb4c5f1675038c3b74d1fac7737b1cd0f0f9c1bb7eba02cd5ca5c83dabffb8337c79e1814b8b7abf0bc6b7287f6b2e894ec93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd41db53df8282faece98914162eca7372180c46295ff66192a73d8200820efd002f9df38f348d0db11159247ba3e38f81fbf632c6e9c70ba71c923550286c2d287e7a478b73a92cdad10ccaa46d4ffeecf8b1b395c97a56cc5a84ebcd730cf1cb1b2801bf8c79d3e721abcf9f09e93550;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd66f4b61f773cd81769d8ec55109631f1f17e033f602b78b6558f6871e97aedcc8d11d81ec608848ff91b56992d7b79d9c171ecb5f9426dec29d231566d2199019be77f9fe50312ab405f1784b29bf64c79844499dd6705fb5028fe96332516698f5817666b9c2ee32802f9ddeef60985;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1be0c34a725d9f8ee17c291708723647940e4505d0ffb722b9f75d2be69d159b504730acce14f903687e53688679408cf2f681a5c19506cff63ce3c1d109c3129f7e8fbbb7b9c6fddbfc7ae45df5673ae6b7186b69d7285cdb839243e3b8939c1674c07b23e142567bf9ecbba748004;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e306b6e5b71b924f1e3edb0bfeb576290fa011e03dbc76da616712123a3dc69f63bf0a44a7a780bf57d7c14700788d80f1453dd481b58efe39735620313256479f55a250a9254774e3a3ab4358a9fb28a35af78095157d406cfc68ee0ec392ff53d41ad2c5adb7df0db5412d991a3030;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3faec7f26ef2ff01c5c14277b27f69b76a265bc6d462ea082a0f05db5b3adbf25a8938bc56b1ceed0d5c33e0fb635951aa8d6163039cf82a9c871fb90f4983eb3439939147a857d7d23c35ffd9904b3c7376102c0fa039f1d0c35ae67d34932d7c4becd33e5760255540e729b01264a0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h314c96da9de27ee73d0407b6f817673e33d85ff59ad0cd33d914e3c0587d1321ab15d6f8b1dcb280a9f2d93ea3a0d02f557b14fd2c84bedafdaee8198a4edcac60cc55aa7a7fae8f2910d216606efcdc2abbdb9deb5e6a85bfbcf7419276c2e7544639aaffc382c6fe844363443c7c62b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbe4da5533b84a7e1f21843b39414d26cc850b19aada44cd4c2ba0caf23b47eca7e40dfdfb146ebc4dfa412170210775551c72f281d05b314aa85ab4c10945f8527bb02e0a069c24c9856c6d731976f08cb93eefd8af432ad3b38777cf170a54c2ac2106ad89139697409e7d69f3c4176;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdb544d7ffc4ae505ee49777b6a9881d8f19a0356eb74d79fe47e5e385b099ef6af172aceec7088e14db1f514756645156b30ba4bfb611a894316c17dff82c179ba8d64586c54a065fc310a0d7e85a111d4d30172280fabf4595ef31c1c702f21623b1f4b5656efe8e81c49fcf7f036e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1670203b320add6964e826faa193133a16a1dbfefe5c3433a5742ff667fc998b7a0f68d2e56ec651f62f61113be1a435cfafe563a8f8b738cac40bfcf42ebe93d38d73f6667bb0a75b77ae578bbeeb7f18250d546649eb37666d26ec25f5db684accd9706615fdeb7fe79ffb89581956d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78e28e2fd5a8f21b5a8d4b2d57137abee0da413e9e238b5f2ab94068b67f79c6ef50d032416482b61a7fa298a30cbf8c9eeff0eeb9de73ecbb02ebffa951aaddeea153f52653e988f1988378d4f465362e82c203ecf821fa61264171d5299a0e5891d4788c9276ed47e8a0fe325a14923;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8b1870129761fb88493c94878d0c3025059a8e322032fd692c1368c33ce1a39df1ead4529982d3787667500bdaa33bd51cff7614d7fe22411e21f206283fac5c25616f79f6a3f73909df915c247eaa135b36c9c8e88987935e783447cf2a5fc75cbdc06257d5470192b98176412f28ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd702cbb4ee77326cc511d8a3ebff4ad1ba6cba6a232b74e977cd909b42b519f1a457800c7b7794fdda2d030a0bbfb57f184867a58b3e902a64c482162ee0637e19c63bcf1d1b4c73bbc00b1f2092b94423eadb925100b61b96a2daeb2745054714e2743b61636452dd8dcfa0ae5f42a02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7423e724010483e4ff09d0f494f66a2baa1b6946818eb2b82b50f5bf09d096910cf30c6cd67cd720000a7d1cc15afdb082dbf06b8b6c2dbafc80c4becbfbcd4a77088e778efc89202479b596032efe2ef3090aae4a8f2f625bfe32b3b10bd71f42586c1bb11cb377c07cc3decb4ed0019;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd97b929737129c5d9dd5b200ab154649fa607a6762f53d568ac409b512b795c84447a9803dfdfab85d49a2ffb9365c94798125c5a4378dab96aa4e420f0e7bde4135a45efedce54e0051b70a164186f4b1d7bd4c839500d149031de0bb4166b29c5fb19ea204af699dbd9760af21e887;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5f58c9f6b5aa8fdb6c921d060de6736b3eb4a161e7919bdb64dd140a345518b7cae23dfab13485aae3164e2360c00f4d783d2abc3545258d7b03363a1474a12111acce2aabc1f227591679bd6554ba9b0b1af376298832e3d4d7b2d435ad8143a79cec8061a508ddc5af7a8415a0b7ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ee6b8d696898f631445bbda1236836f7160161b0ef762588ccc69cd11fabd8459c0976a1e113ecffcc7c415539cb2e39b3044885d70d2c856bedddebb24fa3acf400d00e4b8dfa4feca1ad3761926fb4025fea3d266b88ab2ab5273e20e8ba17184584702d4d38eb89231e0c519bce9a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h866fa498d35f4cc9270b44c44b9c576b9cd2e656f32d1426ecf0a81e8370119f3b89baff4c94ac3f247f3c79970d81d4d517d2ee1aed9e558053b1ef3668222a3b8ed3d8f763f45d52c2b230255810dc8cec8930391b43ffbeb56ad9b4b5d862c1a30c5b66f008b789f4caee5705b551d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e7bcbf360f75aac7730c2cbb154eced319df2b271fcf137da4f2c27490b69143a64cdd0debf388aeab0b311f7a6be164ac9b1783f0e9ec6cfa24f8083f8c0ab0957278e117b1f8ad047947f28e5f63a2e632957b5c124181fa2717361c43d348d553393207ceb06ba66b0dc1918ddf94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b71c22f8ce6cf1a3963c84ce7e6a3c7ee334f5f6d6e34ac8a12fd85ada74dcb2fb9cdfdda8289e87fbebffe6b55cad0224028f388e92e9b9556a5c2b545d2a2ce8472759cb2568a46918436c52e5918dbad8db8eab3e74883b251a95925106878be292075485dac8276bb6c78c90768d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3161c6939c6b6e57ec80763bf22c77bb389dc075484b34e4125d3fe29a38633f7637fc0d21bd1670af881f0f681ff65d98d00e245a8008f5cf999dc2936ea983eb2499f82f98a571da08a5a3917db4e5935e10bfbadfaa12dccd82e557610fb7d03e0705f94ef0e34a6a966362ae139bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he795ca2074ac20f2d9e2dfaf421c08ad6c8d3ea21f6a3c35fade4bb11660aed56bc6998b50e33008d9b696610abd93d74afee7d0647d7146c3e5a527d1ab4313880147e6de1e767335c27cde97efecf35e84b239cc797432acece278627b580e53c6bcce19633d43343abdab82affdf1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2ccbd6c10a0e1d5ecacc7a1c9581df2f6f7d5ade07a6a28277cb82f71776d88ff38a664fa59693563d65932199110159637b69d07125dc96e082c20a5b86a185ff4c5e7ce9b48620334e078eb0b60bb45504366e358e2828b13d9b9746b80a93213b23224d66d3a4316b2dbb2fe4ef50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72be635f3425a8e266e8643f0a792febf18b8d2948ba9a8363a19a9f585f5706dfa65466b8305a9f8af09195f8dd5134d11648deddd2aefdb1b36e88dc154ab94b93e4c33c78db372175510f511f0442c2a4c29e14e8c144d878dc0f1c9bd418fa1fdb9bd55d656be693a71ed93fe5cc3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc6128a02d6762cb37cfef48101ab11c55bd7170deaff8352e2a998e869909c384aab6b4d5140e49f5bef828da30c0a91ccfed239a709b3483928781b1b934a63295efa7ee34b85a07574e92e075669e93b0111d66cf119c790370d3404db6a5bcf0a851960e0ad26d71dcf2ccd0e670c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81d3e17535515f4c17d31e6431ecaac11c07d53af1ec194dbc03d1f0c9540bd6a1c80f078fae68b3af43deea6a188d6b1a3345158293c609701d1a0cda92053a3697d89c74129cb29d9b5a26a7ccd93a9f83fe842a49fc4f037aa77340c789a34468f99ff38a26644ba71d46e00207e4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97ffd7a9da612dbd9e9db80c7a9b4fa851358ac42576e1472c2252ed6d27990698705da1ae5f1850ef55b63f2c70dac0bf5bd4d095258c0db2e7cfe174bb0d30c7b7d8132453ddd28b6e1bb891999929e162f33ee17b3c6ce28c0607174efba406498ab05cdad10249fd6eb561747999b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8694a5be112c08c028b89dcf50a595681f6b13c652df61d8a379e3db4e93d8cfd523ccdd544c1d88a48e7e1c481ef6267c2a873ef3b2d20199c5eb395cc5b664ddb97ead02362dffbd8e2a6d4b57f109601a161b789bca3e3fcc75c6ec701468981c3396562462cbe7448c3a7158262ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f6e83b1f709351d727b80f61a3638126ddfa5a7c3626d0a9309524bc84cee667ca1ca234f692073356a4cf98b1aa8657e3db87601c59a1f5de79238a0eb9c6980feaf84af0d446fdcd819302bdfd42b788d31468032ac977797427abec52b7f1c004e1906e2b31f2052d0eab7a48ae7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91efb26684a54f37c8d9890a55cd967ff9e32f728498ce41e3829b3f830397aaa1690fbdb8d2d9e025ac7b111332c423415a8afb8dec50b781f669032fc018bd1c7a0ee9d12f9258fb54297aba34821c1c3c753e37a2d593bca0ee911d25b0f6c82cea1b652cbba1638c4db3b80980f7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673d83a8625bfbe730ae43a6a89ffd56b89ee7e84f88abb021d0069741a7da7e04074eee42d7a0700f7b0638258ee7fec22c36cde4ee5be5fa811cd9d7e819dcf9dbb24ae8dd1962096e9876a38d7541d1e5e1527ddd498e2c6153818695fc3288fa5741742b5932f1e0e6219af2822c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca400c47098cc99ddd19a5f5a2fd7b4fe23e87c62f48308050f8fbb0c53ff4235283d06a3ec7fccd44a11af0adce7022d8ea82d21378034a1531abfd4731d76a88bad05585e12c60e04117851f28af8acb8270eb1483872c779bfdb3f537a1af3aa514696bf0409b78f2c928304ff9e8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4a2a8d0120391d2343320ee49e7e3438b402959b7038e0017b5c630e4d01832844abc763afec56fd68bf4854d2ad915a10ead85a724e88773e928e6c4824541a89fd56a35c33101249c64c5a9c168a70b1d7ca393f4a6e9930f7afda69124af198717cc0603712f60666e9d65e3fab3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1c92d60701a0800723d8a7cb2bbd18451bff2136999cbb21cd544c23d581e66d20a1afdd3d774788efa33730ad4e389c17a93b3d4e8e91897c2e6885c78ce693fbb42c403df1b3d4d06b17efb4dfaf9c14b93a614110d249a662816b83bbd5c9a6e0b5f2936f20e4a3a7b9432cfc1477;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h717fb4daf1f1b66708a7ec3de93bd5a4fdc032df0d4cc169cd0ef00e6e55bfe645b5087da8ae3fb1718eef12dd8a8a02598c554dac588875b76cf0fd1da893f2a7fd112310837765754ea11fe561522a540ae7a0c89be9826ed87f4317b82d71e8613ad9c079a3a64a0debc235bb93ef4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76ba4f4eabac854c6d4dbc7a62b9ae1efda53529b91a41feceab01e9ce46c16ad2e48631c76f06932fce2bf5cc29d0dff7e56998aecfb5b53826ec01cd7e6ae330ecafd8cae6a2d003ba96aa90aef764cae46087adb8078bced18a4addec3fe31c3399746d11436a5578daa505a01f300;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f96a32ee3f24877937650677b809952fee16bf7b9020787efe5491b36ae402d536f43b6d0a86da6a4a8d5f754f5a51b25353bc076d6ce97c5a590a1be2b06216b29a7fd451e4cddb80e1c1d93112b2b9275edeb3f93fc8f3d42579c22461c8ae9e97a7b9994d095f0aa0b606ade42ee6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39a9f64f73d59a71607992cbde12a78397dc1c8fda1e5e5b86a5badb7b80c39607b70cd2da42e9693ee9a2901b31ab03a874295ba7df119c168112e2de61ef47828b1fc8603195fbd4141446b1b9a9b5030ee5b52b604fbf5ca379a2236f08b5aea5d6882a1103b91fdbe0db5ddaba3e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50f8619d60b737a20a8ab791f1fde6766905e7a99586f78ae8ffeacedafdebb83bf05ff8fc1893d50e3f4d5a9f9c4e55a9cc9a2ad18448fb04af00b9f77d95847f2612be6daba42d6cec1b21e55af88a3ca537e0d2eff8691c64a1984dc6a8dc5445a86412d51cb0f68ca7ef68a2bff9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f0c400a7df0d314e1eef3a4f1f1577eb67672eea28ddc2305e7dafac85ba886a8a6b4b98f741e595bab9cb5effedea550f8b8e73b7de54e313e1ad5e5f626b592e06237ef94dda204bc32b420c4e1a413bbe75f00b7dcb13b5f9ae089058b5be7a57faaa094870610780c2e3b2dfe583;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda5a517184d32356eaed4939fa97bc74cb844b651a0e9187859550e4a0270009fd50f93e0e2960bd5a0320d2be1d8e36cb67956cba4c1bfdbb78f0567c0188ee76971867463b40bad922d6a46ec988c685c303c404b7d7bf9dab4b02c9582f7ca28eaf9489125c93adc1ad68cc499b59b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b336516463b968c4cd8adc85da425129c10b1e199dc7563e1d4b79a64bfdbb4a72309af044721253248d6521236df640f718ca085f894842c4138c8bb2df84a4c68c11bdb308464191325851454890a48342d936be3e587a914669ca0529503ef2a1a3544c07e5282bc7f1edfbbd0d2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h350d926de3ea367cd160e503e319f60241358ab55ad33077c88d3d4bf6d496f957e2375b019b000b8e0c9766b5f09a9d6325503cf37e30f2ef5d8e0e1942e5427f4944520f28ff14058816c6b6a0d2824f9e9b933858707afcb3c2a8d78d8861b54721bd571f8b068688cf9c2ef9c5a85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61169faa1780fa189913571f88c2235cf9ecc590e0cfdba59caa4c9d098acddb4a4ace2d9e1d81d859257b17c08a252a315aa79a5a8cca7aa5daf8032c0ed7ca4343ff3f7239bf4374a06cd291096b09d5681537353659d026417c46c1e4d79ada06f5042e902c64952e508975237f3e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef507f8fef926677beb2305456a62f17648beae21f6e61065264174d5f349782f89217b6841eed709e1ff24b5965961fcbcd4d0c6eb7afd8af07c0608dcf4ab4ad77153566cdabaa863a801ca75f7e55da79154f78ff5467574e12ce8bada8d1f4021fa52f04966a9b18034017f761cf7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5166d0bfe8ac7cd80d3b56de2e969bd23817a45a7a95be2ffd31964ac2d27fe3fd98b5892364717fe2b195a4b872274270b785427d222d199e6a9c8b46147ab08cc4de2f837a5f8a01470268a8134ebc3a3e973307f777a86a245a1f1257031d85d715b687e36a733ac5c24bc35e32fe1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha920a70ce78816efb3f0a5e388816c9b324585283baa23306381726fea07c1670043d6f444657a84369f10683a8ac66f08fdcdbb822d762d8521c160c266b3cacf66c91c5fc71302388f2ea65bcca2f9fae440481b52ff77d29d3066606e8e23f6095aaba87e98456d580e409ca0d03de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8806d556f3f8f74f7b1e02ff3a4acae56e443d05fcd7da3bca89dde42430ba47c563cab738356b75073372da4e38cb827b304e8769982dbc5cf121ed2350b84af2397d7c84bb77b73a16447011138dd954bb6a195016aa8fb7d92c8c0ddd34e10a77e744c86fd12def42442d0e9742d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e883e9f751f1148722814248b19e449499dc8a136329b3409bb37f50582cc77ec06f964fca743073c5b2d2b093aa1ce1f959a2bfa9a1dc79eeb804d26174693d9cf35204ee926391fddd7a086783ad1edf814270c280f344edb0652a535b86549a10b4ffeecb4497bc215a423b9205;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc251b0a67102c3ffce887f6f2ba4e9015739e4a1814fcafbcf1ee1101d96d98836f4f7804caa001026722a5965dbe56006b03ca18c48331bd0fcf6c13d2aa69de52ab1b1a84630337619be5ba57254188e8ba03439f111f2b1b0856bb1c104d8914b1f330fe82c79f43d944745058aaf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b93edb7d86285e9e6814adc5ad7187610a65ef54961f50c6ba1bb0a06e9b47b9cee1b70b2e92e32eeb246ea5383281fcc16e3dce3c4ee4268918399fbfab7338019f5bbd5cf98bfcfb6ffef25e9e8e4d75903236f276e159c4c40ed7221da6acba2631ec02e4c736801696f5abe091c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h991ee94abb67f4b597726df68d8e1ed13015854929b2bdbbac7746b8336f3ec97061086f31fd2b5fcf6c128ce327d69a01b6a709df02a08fb26b34c908db1bef8f39f66edae6f4d633e4389dd909ee5af4fc2b3e4fbe65a9b1752938650f1aac89f07a677d17c10d9dda90ab7bb05787a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had944783f3239fe35c70ce5b5e337260d952be4873c90dc14a694770ee999a6f5d48bd3b624b22ad8ca0eb4e218376f361f167536e2869d4995c38352f8e8f37c8657110ef2b451fc9dcd7053fb34bbc2dd01a3ef86cf1803f52f5295f2abeea2d6e481eafbc6f6238f2a6e00a3a475a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d8f026563f6e51ce1074b0176a0fea15fda80a5d4975574ca66ad1a49aa286f3a48c02ebd8f4dae208e438239da3c82646dc17326fb8fc783168cfa690f00aa2ed3b728b65c72dd9c432561ca3e4709c727fa20cb318111387af51b6c51482765cd70fb49ebd6c919259ee466f736d3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h300137ad98230e57560fd52412489350eca690d4f5576437ae71cf17aaae00d55a6d0137d881c7d55fb3116a89038e46cd6a2ee2051023bc6c8ffe98fed06320d537226b5f764326e16e9e2a45613476c5b424552c155d1ef91650ab9fd42d6c6d473503212f62a0624bdc35448550bd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec1f7bc5c1e3a6e4c2ff01025d0474cae88ceba7b828a62f33237215c7a27a5c33601a84c1eddbde488fc0dba454f70b64acb00cbcf6eaed997c27f53174120a0515be1c008fb2474979aa7e61b697ea66b89872f016eb83066a84d0b9a757fab395c6f919d3ab5e35cee0906c5adf5a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65e2819d012ba591480232bddf9becc63a5dede27af4d2b9cf99bb148f40258c2ad0768cb22aad153dadd62af2ed0086729cc91f5f42656932bdea38996624b7cc9f34b6f6548f685df2f70700bc908dcbe8a6b191890549cdad9b361b5a10982ce453d6bc634ee38bed6bfc8fed12b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96b0e05c5e952995f25aa28ca7f0b14a96e8bf3eaadeeaccb903b5fe938a548c3c096db802382a0e331a6c363ed9e50c506cdb3dfdf7b6036ab71bfb1d5eac4583e9246f08cd7e69032474e785fd1f95e7886e28682bf2ad6728cadfece2c427a43e72780b994d570b8caac11daf4a072;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb706cb9c97653cee6b7bc7e4fc9d4c094d0dd3baed8a0ec5c63aea369e1670d32e6ff6ea042c0b2bc76a2f57267039bf21798431a1be07794db47c858ac4bd4f84bba8db5b6e72ecf2f0a6bc8a0525e8d3ba495c058bb997a48e718a9ee7f3a70f0911e886e1c2f09c83d0bd4877400de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe03ce6102491b31a6d0e740457fb7ce3905e97c4652658c6d300f33ad05aca4b0e6189806eda0dbcf7577d5ab1ab278444322874f4311b6fd705d644a1e267c49d9db06433b2190d4b75bf1ec7d5b36af9208b12c9518b69ae2f7b3320803084b749a6679c4d18e9483784e9e60dd8aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9cd174fed3c130b3da6f17a20cb96f1ec2f59169d4e0dffa09d8d14109ee3ec8606e243a1d3ad5323143898cefe331972b1dbe86b7ff54409ea36e7b6326d19b9bf7024ac1dfa6a321e50f42f448dc751664f5ff942147c83268aa5bbf5fde10b97ce8a48c1e9b99bcc6d5b01d29b7dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd068c720a9506f6c546064fbe399434d5f68b7a895d5b7ea0cc9476bbe2bfb3d11a215cd756b3a1a9bdc92f6ddfd210b87271e718d2a8c3edc9863c47e3b96c1767ff5170a1843612680a2f07b17dca9f2fcb8083037dd58e4adada357208e87de36563afbb9539ac8a1ac7431e7f501;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf552249534f64aa33535bdfce48f798cc1da02b6f09fd3a0e0438326205abcbeaf3c3a2e0e6111c64ae42a642bc48527d76933afb6291460cd335bb6db8f7d8cb6e9791fd7a4f6ede57317064c38203ddc24528205eda478704e5d9d4bacd23f7395d17e09633e40389cf24e2411d9e83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h640d9b4ef095670b7eea24cfeede926937297175060bc8ac20e58576e4454e9278d6d0697e157b008d55f99d0eade7a6506377889204f6a9936478435bd05026784a47c183f55c6e55bbd6f013351504f2ffd32ddd078dada46dda3650e760673db7f23e922908a005806ea3b5237c956;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a76fcab10d25a0262aae6f61b003ca7b8209126e0950df61dec0aa240eac389d90132d9beebbc5a20ec025f35e759c448ebd48757f86f13a240fe0a26f65028c0c7dfe5ff2ef49fba57d41f3dd22fb5bb128eb340bf121989c92042632d7c089eb82b4df62b2d52932080097d42497fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h833319ef7d8f6cf77de63694a1ad729b981f1e7b95f22d83235f9bdf17228bb219bb9bf5a2fff81b70131b30479cfb9794e4a41422174ace1720773f3cd9f27683b4b6ac8baa8f79e3e1fdde382b06fdc18dbc85070482b1df3734c4936be6dde1e30adac90097436f9ed174616c2da1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9642e47945227081a56e300b1af88c0b5a97f15276d8179ef10360ddca0d72830ad3bc5c3ae23d7fd48a3ce338a16880bdfa68759ff0bdd9a04b154b96917a008ea587780cfa5757914759c18971b9e989041f8322b1fffc6442d5631983f99e59801befe9a4bb353c7faeb54ed2b1b3c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd4e1813102107d791bb186ca9bcd4f7d3d8f9336b9848ddda513417302470401ddccb5e330bfa7480b3c6d071ba8e44cdf59a10a4b167a2f73d3d19458878b8c9c995b0c553696d10ef3f643295037afe0cf8f2f7610c87bfc69c560977fc81e2a77b00e23082d9952b99b8dc67e96ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed42b437b447c21f0f334edec3b8a6a771f83cf2c275a55c92e8baed33b2c090cad508b086ee20ada79b09a2d88c61383a9a928ca30cc3fb15ef1a5345a5a1720e80912df36233b4d30b210b2eea5a7dab962d5747d119c0ecaede561ed3211dcf72e11ab6147375fc36547f3e347e4a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h934802628e4d949af9db35925a64e773ebfe3c498b80cb6a496f97e2ed4a2d286bf3bf86507d3a289884d0a15d5149d00babde0d5821536df0b0aca8d6e27e564e96ea24d79e751da7810042f9fbdacef65c48504dc1e28b1019f63fb1277294a7108f0669408db39089d1858f75e638b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8467386f97849399d92932ada57989402ad606c97249113eac703f62986588bb3d2b3a28c36100b306f038b45def62809301f2d53d18a38d3fc1aaea3706f8d07479a1a8f5c3efeac5c343a9fd9430e1c7c928a7f2163a4e30030ece43249d2cb28fd5543ff3e91f532951caff579b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3339e11f102d886d85feb2b56099692ea1b2931ef07a97bc60a2d12f205460006e0aa249f1c123c01725099e4a8842d32cefdcb7302dc07ec4dd3f4664eeec6fd52af6c541e252d3c642cb793214d2468b6ef54384d0186c177c267e749a79aa82d61bc3d36642e9488719604181d63c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h969161345d0bdfe4179ec23834c353110116080d098e9f04a5033536328072c04a047e806a4f32e94883111369992f15c8ca2cb47099df8b32b817254de81b878b765bc1e5b481841b2e72881bab0e28ba4db63f81a3bf108a11fdfed1fe4b01fd47290043aba7e724f08956e88afc95b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7efad8098348ea50b0bdc63a29a322bbd565ae9c6518b77a6cbcb68c54f5949d351f7744c37c40623fa43861bff2f76cc7b8b5279ee2ca4230558c73f163d95697786c003c868af66bff3bf58a9f9d7f038528f04b84ebb4882b1739eac8fff7753526d3482931cbb96ee8904d31b78bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb614df0f5e7bc5007ebf905e1ec7464b2c0e7295b6f9019b1d8ab962e257875e70201a4bbad6685e4c49a29f4e048613cc2b5e0cfdaa26417229f9b1bdad00ef7219f579546de5c3730ab1593109b8bfb78010797eaeaae10f1644e85e4f406482f10210fb11bc31bf91f6bc512424db2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9070e8ddcb886e9de90c124faadffe2e6ffc3eb40ae15d672539b11f968504f6ef17fa4b07f5ddc632971c56a078caac995d044a2173ac5988f446284a553eb01997aeaa330de3050d352bb71cfb6e5a6d925efa4c226f889736e73c98401d53f522fedbaef1b197bea06dda57cb1435;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb109a911dc0860ab24ee10019c3660480206e257d9d3bd061548620c955001cebce7c6783570541eabd943a5e0a9407ec699147e902e208251391d8505e14e3ec3e69affc1824f23bae7ced9832b2d41039959adc7855ea58ec6a87072960cdb6bc1fd98b7eb44d59a0f40a9072f370c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc18116244ece28795d51ccd18870f9b024713e8296aacc66b621285ceac97dcd2d36ca2cedf526d4c288a710830bd444d0039ce53f77d1c9b1fa59e6f2b786009c32c6fa67a29ed611452d23303ab775b185f9665b28b759e6390a331a99ddeca5d00707275001fd23be54a5ba4960673;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7a4171e06a2ccb843951bfba61b84a36ae51404b9bd20ad8337eb94705c256084cc277ceafa593ccc54ecb00acb68f2f4da2b714667aae995888221d2586f107e2740c7cbe8cb4c540c134e7343c033ecd97266402770fd18da3a2206fc5fe7987545d8b20d1535613eb5f28756b3225;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3750132104e0f24b8c75ed88c25f860535f3da859562990ca2442783de6e22fe6663a8cf55d637ac367efbf64d907252f1d347d3feaa4dcd949175d288f3eba66726f0569e45f646b3f9340480d67d7da6aa8ac2146743bfaa4e4adb71be507e1f2acee79c222fa83267dd841d1ad5081;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36c4fd3c4649edcaabcd6f00d3c043e9bfcc48550f21972ca2aebc02ae44617fbe597dbafddb09ace3bee50689f7d8d91ce78c1c1e059ef29a194af3ef6917f66feb009e0af78dc5a30039f0f0bbeb39ca1a0dacb52f1c7c2d5fa889b3627b514a9ddc66b23e5ea4ee7bd31366d4da5bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha34fbd747e344b37a156e4625d59273c6cf2733b45c9f6fe266d81a9b344b9f5e6ad5779bb331aa8770ad15c8b53dbcf188177807f8cf75d02dc42fdcb11910fc6fbe7225a8ca15846e0fe1003cc0218a6f0e0c4d25a3576e54c804d594dd0132a770913aeb8477733a092a542889c1a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4402ea099763b39ef7442b8383c0726b8f139d8460f26032d0da92e64edd1001a69098598a89f4091f95bb0881055c14b264155ad993a549a104caf1528475b7dee66529f05a2a8a83f0f550d0bdc0ffb5db0b9645aa66fa08944472fb5d3912e4aaafc915f580b8d20c0ddf4d8793b0a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b5744db9c835626140f22d8c98642f86333b212c76c5745700acaf1d9923079e64ef95f0375c03ccf584e258d0e0aaeecd4cd513b17284275015c561048449c45a794963f552d0049142e7de2c9ea774af711e3e3c7a30cd10f5834239507ad68eb516a4f86e3b6bbd0c1d968db8906e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0b5be95baf6e1ab7c03094dc1d6806f184ad8db4388c967eb878745ad976011820d9ed3ef74ef1a1ede3b8fe6d97a215ac60a3f467f68eab7e813e95e70d9159d84f2ef0acf434d514482429c5577fd001ea296b710b201a74fa7b838f70450737cb876858e5dd32a8f7b178536472fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e76d251507e693b20c10fab3932ed4ffe7313170e198ec09ef1b175f0fa94c213a9ece0199495fd61eb0ea6ddfb095cfd6e6d07e67d8435dc06198998ee0f6b73b3de5dd96e760671f4596a8592fb9e1421b504b1e35ebd02eeaeec1bd3f6e98a6d00f368bd6e6e8e67bd1fff9674746;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h315ef9ad71bf5e30e18e10085b32bb257902787db7107ba260cbc289f93ea691685eae740aad5873104920bfe911366a1f8f554560ff1e8d1116ab15c9c52961058f79adaac9dc9bc57b8f3b7f9fe2ed507ee2ed70fd8d095fd0205011f69dd63b41421b15dd935415aa6a6c0bc05fa00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h422dc3cd2d7c5c6a2001c6651dabbcacf4ac59874e0ceec109eb0a6980b8e49b8f0672223ddb55664577d0ba1f1bf42e48dc23eb4b35e8945d6723d3168012aa5f9ae849eaff242f21328d6057329709e5f77d52fae375f75106d2c54d573cea5ee0644e32ec167ff4f8236fe4d928f3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e57a00d9e247766b7f7ec8f06dc087ef584661e73c5738c68abfa5afd8101d3ec1151701760e43e94c048e591bc79fc0ff4ca9670bd882444f4d01faffeb83e31ddcfa356ef5bde0bc7700cd6c4c5bd5958bf4be8b1fce5c308ed7bed10ca6645d74c72fe544199325ae4adbbc129bde;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2f1cd985975bd63cf1f0a92527b52f52778a6aa10c9920202ff2c232c7e631f4810db3b0e65020ede915668adae05fe422dada1268b785375a7cf5b9028606d8645067392b1f4e774c107483a53661e39d82ed79cc16e6db410df768acc9b5b402c65a491cc5db5c458eafbfcd969920;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3298197f9930ffa4166a98b2d03019b0f21b59ee9342c152735a7d1a04c5fd68c0ee19542dfb378e88ea0207ef9f6a49cd5b851ef0890f98879a4353638b04d9e45f59e6002bbf454f91705680a32f65d96e15ff675fc4e63cb6265077c6189cedb1d9cb864b0d784f9a10b21b51c865;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ff2021e525be9b70319b0bb3bf173c0de2ad66e54a5dc8666a2c56d67f89027ee02940115bb22f6b0cb267b58914e138386037e18661bae7a1c526b03d85e0b425695457b017125d6bb7167b02bdb83b31815faa03caae0624bc9a9d1bb4c08ea6a37bad9076cd66b2e29ce7303468ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d42e902c00409a33f62f12c9c0fb82689f18c9ba24df992f2420cf5738789a9f434165b3fb18e970336a016778d0bac1cad648a39d5b0e8860743782448907f892fb66f25b936ac9d6e79711adc7ca96b80de921ba1937cd3e69fcb6646c956863b47e42b20d26c9b43ba5d18c0a565;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e639bb535b4c18fb07e75fdbd73dc2d5abcec7fc4608f9a9380f91b5c000a9dff59e526ec5b7fc5e04eb333f33c1269c10734f72b79afe7ca9d32ff5f29777a87515c1bc22ea4d649c455e97475ec1aab9acf7d352840539ac347257ba1be03fb3601d77a3457f216c8d9c12798be633;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf48373dbdae0ce2ade6efc443ad580102497ee568fb3a07e2f14fd6f3a276d55e8bd383c2f4a2ac3c08b43b6f21dfc3094159284e85f9224d954d5a885cb2606cfcfe0fa1c739158d704575e1ea9b2943353dd07eefaa376285fa1a8392700fa7010a9e2f5935f357355028670ed7a2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8346844e5d35011104042f90c9faf89650d0469b2c3756b640d3c6417e6fe8145e07eaf6b0e3e65f3b2423ebfeb2ac47002fc2008591316eef6bea2aca841df5f9ffa319bddcc2a0a31859eaef9d82f542433e34eb65851f5a9bcaae8c2c2ec5afb9eee92976fc86450dea38f2eb5ba91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b091db740a00b3b4193ce4b6706ed39568030fd00372ae1842a445225f458941333d24ca101eeee17b61ae0dc07ed62c4b151e05a879eb0e3ad61774f8082a5f6c2c99bb103ed48fac9608e463897cddf339dccd5c00bf06fa9b6b86d8ad0fccab852a4679a87a5b315bcc33b5522e59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3da5ad339435c4c6073f2ff8d081d2d39504d5565c37103efbda2b330d8c5d9ac55ede309d511b03fc5fbe7b4c81ac2ae63b714912e6416fa5cc229044501fce5dc00f8e4f95dcae3e857d09537d97204bd61b136adc90ba1236c9efa10d4557fa784079d178ff3869fe1d0d7fd143820;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h451ead4daef632b6c60731112994d8b8001f4bcbb267c3603e527c1746b6aa0f3fe5de1b79123ef07ba33c74d60882dd4eefad44bce01de9861f2461e4b7d3fb5f6efe5b8f04358a3e19b5064eaa96aedfab7ad720bd4a32a8316b8082cb1b3e321a83f5892b0d0115a3800a4af2ce8ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1246da51371e1db433d1ea118e1c215982ad6c582fc2ffcf83915ee09697aece1cada177e33124c0ebf78f91e992a3d32205d468751753c3a7ac9fbd882e8c9c744f07668983df0d750e5e2a634588653cf849e3329f70ca1a78b0bd6834df1b9ccb41687c0138e01da5702a2624f3f56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae653e94f1bb26ff962df04b0f39eab675cdb326dbb1c4374ca70519dc3aafce9a1374c023d21433167405114beceda02c776b07f720ceb84ad8b5a07a69a01f4d0f14c0fa7c4ad25dba9181640e9faf6ef7fb88b5db835d50a20ce3a470e70e247ecd065b3e71d4f9cf275b1cf0a3b7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6b0a3245fe3fd407779fa8238a41af3f84848c21bbdac12747f1426b29ad0418f9fbc48d76b46a013cadba3b0b297e4660892e2aabef4569ab8d96b15df7601dc1584def4d3fc5b5c62b2706b08598b38a861db68f1749724af12bff3fa38744bc0624babcb738c5fc9e7343a1e993d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab29619095e31d7e8c90f4c5c64b5ed0c11f49d52cf22dbb09b333b3743ab39bd2e6c6ab9f9ed44872323ffce00749e7a2d958e96339d9ef7ab54a22de6765d14fd40b9026e464c619fa60ab12bf4795edc8ffee2e17951ba6e8a54aeebd3a9e8ed4bd0f65cabef9e106fe2f0638446e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8592e4d0d8572c78b318d9a95231e9501c74d8fe09586ce6012ef631e537a6dddb965f8465b723400d8e8a682a2213db5bde5ac4f3d5f18c6335198c1fb6c59a5630b29acb597c3a2d07b83bd22ef1e3c26191bccfa20c4a95a04e572f6e132f275d0f9989fce22639c1e99c81e20051e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1474b7970651c872527f3a27c55d48f7414c9dbb4ea32a42665c050fdc96811844d84cf5a9d1180a1d3365dbf26d1992e7eeee3dd3f025c51ad99aaa5d58b4fd95dc1d322f913f8d69de30e2a756b0ae0628273dab5aa8e42c6046941e50686727642139d74fadd2579c63eb5a7ad015;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb26782fb59182085a7eaad7ca1f58878397fd460002a5a05d2345f85d6bfeb758e7228c6a52c00e23d5d75d3eeb539c3047580f5d1313f07898f0e31bef0ba2304ed50052ff7d8a03a8f4763f7264ce5169e40ef0181506cb2b674c8e103359d440c5175a28f0ca7edf22b3b7df88e36e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha260b3b1d9e2db55aec0304a59af2bc8f0d10cfa07c1a4d7a15e7a80e4646fba727a39ef2020c0e4367fd4aa7bdf2d0672e1eee884610e7c4c6d347b304fc229bd5e97d9a6fb5319a629cdf0248087861544f4e5f4259d5225a8eb1191e996a4aefd05f5b6444b16ec234f0f7405d56bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12d08cd7e2c1a0979270614575a066d75fc8d00a079bfdc918009723cc2bfc08b716d1b0f69ba014d543e0a708d63899ce8fc790faf56d97beff1723ce30394b23950e3724d5d401b7ce8fd88fb35d2ecb6b6a058f1dfa4a95e2e076c124830f6225b215fcab941ab2eb57b46ba3a22e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6cd396aa4cdfe5be7cb2456099f6acde0e6af53bf4a562f4bd6c832553d6df3aaf7c184a73d53b23cf2a32ddd9532bbcf6dad3fd13f470c8f7b94f3f9f31207f5527822bf512862edb8a95936de0e536e34a0fb5a4fdcd9d3719345304574c6c39d26d44193a67bc631cc79ae5d2dd7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c0b7ae42ae7d21a572d5d860c3d68ddad8b913157983cd54cfb983563645845a03b206c55c51be8c5aafebcbfa5d6da234b050c1cfb2b31df4f9d9669f803ce80cf6597c2ee42bb1aef05fd53ae5c21406628dbbf8d5a78bfa2db4e11f8827577c72e118965b0f33bcff58b95a6c9b9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c05f5d7313deb9484d4b4e73391a77213a635025c04f070ecee9be8b437bc7129a39332f1984e921a1823f58ccabbe06f14b0165cd9f090c18384f58cafcdc147f81dbce6a2a5cd9f7a4d408e2df097bb934bb8d3b3db661e53bd89aad2393fad2b99ef636d0c632e4d5d5225067b2d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h741be21ccd980e4f6320f8741b11371e3b7d928bf25e8de691c9744b916b605a65a5027b91c15b51f2e04cc30720fbbe621e005133ed8d4b5fdafab73e84cf7d14d851109bcf89b7f77148060cf0ad95bd7f7a2044622c5821c5e9f5b66b06fe5a46177ba82da5902da92e34a84f8e82e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65a8d3a762e601dd5d158e1f7e98c897871c2f8adcb9e9f835615f7941366a3d813fae2da8bab713181a4131a784dc38d12d7c742bbc76cd55a3a70385ec593143ca914256ca628d12da18a0083d22f11cc2bcc77c27995da70859f3e71e6163147d78cae460e292bfff35486f413ad0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46f9f796874a634dc6dcd1579e1a4fc5e2c41c6db5c7676f520782243cf0d5068c4e084608221c46b08912afecddbfca4dbdef3b0eddfb4a60f686e67a8c016dbe86f3464be76da4a80955ec14e6997e6d48f8452acf6b4bb1505c5d0d9b15be463c5756c56b66a446e032002fb123450;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc10b7a40782711d81f6b77fcf0134080f0c9dadd7bccbb853446b48e853a32dfb732339d38feac78c783d86b9acadb47e5096195190df5bd47c4d24544e7a5d68781a3aaf1afd7e0d8ac1f5c9a1f08b1683c04ee734c8c476a4b00957f05405618591dad90468afd4d5e77722b224950f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h666b7658f527a20b2e4d48603e4ed028c612c0683acc1b5ddb8ec8db83da2e2aabfa92c5d8486b059164e47db365d2bfc813153e7cbf2e8b66dad634dbb6996e7252ccc0ff4b726128edd5bf12dd81c7afe97a01ea3d1156814ae6ebc37c799c55ca19c6e4337fba72bff709b16d65031;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63415b59b60d71ec42d1121e526f1d5e76354800377e2525878797843aa3b5ed1ab37a1f6e67b9effe6121a9f495ae01f614c3dbf2b395f791c4d15c9a65ff9d55f5703d9284c7da41c1c3f4cc3958a9545d843c2c4233e4a2b30c26798b3f652eda9a47aac1594d3fc2caab16c0cce5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e6794e9bf572b802feb9c39710a0eb5e7fc329955302bb6a1dcdf6970661362124517bf787128afb20b3a68d6592a54e04dc00d6e623db8a604d7193c0156d68df0203e871a3b4d4706b1ec42281645ed640b883e9f885ee9240e67ad68db72850dd7e834feb9ef87bc48a9ed9700d92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21047ed2207413e24c16f23b45adefbe0b78a21735cced4fd9c6fa31116436329d1bb7b7d5c66c40d5d39b1f572978348f656332939050737700dcda37650ed459d775607c9966a2d1c457d4347aa71472612eb4120130ff634894187e2f8901ecdd85b09337cd6f669437e1051a716e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h633d7bcdb20e111813a5c470fe798e43cc35e328f2f2a638013c59562468ba4b5402a7fa72da267aba7442738b9cd71f152d5998a85c77ffc916f701a333148c7ebf0d42a0df8908975318a38cfbc969efae36a704bc67108b9533ac10592ed9fc0ad215c9d6f1fa9aceb7ae1a211c0bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86f05b955fd9cd4574dac1e19232504d123586506e8dea903782e91bf817eeb7fee0608ca34cd0ee15943f6bf3e6a300bde3c000ee4b53c1afc08832e627563939951239ae86459cbf9ecfbc4211feb9e5e269ab47e8472e6dc26f4fce2f0c867aefd303243982deb9d96e8f9c30ad585;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2f2c32073111c49ee2a5cdeaa876aee5558ed0f7fd55f5083b873d2a533436c5ee9e39cffba7cc9d4efeba1dac9da0f614e9207a80bce6150cc8c0eabf84d1517388394a2709bd42a5cef92b04b99a4a70854e05097327f3c4bf6c1f64526a1c20efb948e05e9a9c0fd9c3dd8275494b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55d207460a3bf497b4732e0e1f7134ac001681ad049b11b1ceb3fbcf203dfa21dbecbf1d33989913c15553b621c1bcc6a094cdf8f331c62b2819ea5a312eee4522c65de09835ed50221d0195b5b3fba602827b9996926f75ce45b44a59d4cb103718daa47cc5f0fe9aebbbc0ff435f4fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a8128d53dd1024cab074b0f06ecbd8352fa82de611b23862763b0c040ebdbae6bd887e629454df8ca1f883e30f43ccaa8a137c6d8c71863e4fea7563d1e4d174c6b268651be832b22b0f1be426d80fa501574786a788b3255a1b655a0b6c03e497e6c92595d993bbfa979968f8102788;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3abffef4f23dbf47fca6e22f2543723cd7b26fb42014ffc756f267207202e539247856cffc229487e8c54df050493bac49a59048bed20350efe77263b259f338d2ce65b943dea6324430fc5aa137d486beb0d9258be8f8245abdbf47c51f986b3c797c556b34c0432a97b93de739b9b5a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dd6cfdb63054a82b5aaeb936560c8637d67de96e2a28a4454a7c2d041939f01f5ea2a20e4f684d5a28c3c1090360d7887432dea17981deeae5384afb8c49c561c27089bc71099fac492875f7ee2960509bf5540d5cb3ded299167ea20640d2101ef9dec8ab28105c1cc67b532958fd12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9935719c28ad1305bca46671fad077e770fad1956342cf6cd4c86462e2d6cd5ef27884c0ccc508f4b638c28258a9adca3f1b4f4ae2bc94a202c6599f8b7c034d518fe111db14d8e961b9c5a4fa2ba5d53231fbe830d3cd3c0a8ff67aacc0d38be07f9702b66b3eb65acc748be86b96ffd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6db1c9f738ebce5b2094cff5cbe6968ea02b2bf16802f9f5f938f82f5b665e9161a888812cb4569e15ff97b5951cf21e0e7e00effd98ad5404e2c69e9dc7a701cbd23e9afe6157d2b2d338f13476b64ae26e9d8148f85f8868adc268ba5d11929b64d9038d0c98440b3620b861343c830;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f32dc3c1fed024fbcfe2a3dcbba9ef525719523c672d2ecc45e23e152be33df32e85db14ec50ebd75cddbdb410d0b6f24a8bb206688cc0ba4e9fb7ef8dcf685541b9c9c48c7e5833c3a0620f4024a79d6b3ce6ccdf06ffffe19c85b66d23b77da3e2b66a3e9cbd99e6d2ee7c4a9a79f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93d66d6ad3cc8d88fd010a52c9852b2349d379af1f9acf529870943e6fa0e37c8a2cb70e7d30e4f7d49c56597e4cdef81de4dbbbe56c6570d38ae0100dfffa8afcf0e6b4e2803fd3c4bed627b96c1a8af333214757e5f7165e502a1ea173f73387e99004793ee15393ceb156f4ef9df84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bd5c9d4c1676a57f0a04b3fb8507ca6b07af264b9738fc21d565b973c475d91bf68f4bb79227faa474514d68e5c8bf9198599ad40bc5a1662dee750af9255dd0af5b9b3477686870b9e8717d6acd580c5e0b260c88eea886fadd61c640d60de96fd0489e47fe48e8168f8c3351171ea4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d4c5e63c451da28597553135212f9b4de99af6d248bdb213dad650b3e2237a80c1d2c33b4978907f25229a62709fc967163721cff0eebd7c0e27aa3fdbaf951d9c8599686b21c6c3c3ab28bad46d6f3e054772f6144ca0b4c0b314a75bce1340234a572e470347bfbc985eea36c2cf70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39ba4d2262b9669c58ad5f4df7f065532f617383de9aacb868067e3aaac472675e25db5b2e7e9a928a074c53a00757ca54c23d36b6bf5b9bee01ce0f15d8e7172f2d11410ea3e8b44958c7201e5808dbdf7166c9069d2df89af405ff21e17c4be31ba86c156103016a4a712ff6b99ffac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc3f3a1ebb9052509079b3eeed68f02a563854e5d4291efb6b2c1eccf213867121cdff7a40547d6275c1e7fdbde74f8ca15cabbd5f774c1153ab6567305cb62758d55e29c0007f0e9e72b692c892c469b00897c313cc7144131ba9f7fe48d9ab9b0b99ebdf88edede3cea59ba384aece0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d0894a0189115a1b480545fc0f52ec2b56b78e1e0dbf090fdbc3004ad1c3b9ef9bc8550e5cb2d2582ab61baa90357ac0a89a4e9f4bd01e505c921b12e798d6c7231d645f83a4e9d689cbda1e3b72ccf5ebadca154ebd9688852013659658370c3c75233ff67d5797c8d2892cf1632f01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88bedf50f91682870370a0380694a501b8cfabd56ef9c93ae1c94a63bc2446fef9aed883ccd749270ae5f70128993710a879702b2bcc76c7ba0126dfd6cf68d3d7fb21a7fc7d0c00eef11b14086eb0f44a609a04c2420471627c749d36faeaddfbc7bf04e33601a764ed6abc74296ae2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ed22c669021be0d2908f3dd27017d34de8a40f29d7aeb2d9c4bb541364bf7f0df04e1646a8bfc834e8b8d4943d377fa8753b71f1d6c3cd162649b5fb4bd86ab9483e08875718d20c146fd004b40aa35c9c9fcbcecc50070da0e2dfd874318b0a8242fb0559f52d6c2cb05853da71e988;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc82141c0f2521368168936c2f40861d0a66f1d80e9db9fb1b1a94656a107c89e29b7766c37735eaedc33f495d236cc1a5eed714055669db04ce423f5c64a77dab27c977a411c13f16c14351341bfe1209d283176194f1605fc15a1de16bce9c79176133a757a3a84b0a6632ca01dcb25e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c29ff0caeea2fa9dd9b2937d7feaa24febf7ed5f563a4f0544a835758c00331f37d83e26f7ad55ea81f1d3b944229e13617f4cf021b44e5876603d23ea8d1ceb81781bc160f13f56bb2105dee4e25258f7ae4b95c262fb9e6d911f1dcfcb077cde53df3ce9abd3d3601bd8e014267e83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a5bebdacea32097f8470a1aff386c3415849e15fb1d22ae01cf52359ca3e20b0b443a8925107ef80240285d12cbb43fc63b8b2a318ae657a4a10b40f724a2e35fcee9fe4a97efdea655142ce83bdd144e73e3c773d3d9a404b862c905b43c455fdccc607f5530825e4eae982ed65dbff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e8a5b50d3736c95cc316eff2662e656741abe9a0cd6eede4b4f98fef197e7dcd00f3a6be7b2a9fde0ea5e3820f29f01976c7948989ecd427c33868617f34200b358a823f6a981cece47b11603c9586f69d0218611c500d2c5fcb197fcc6d92941e8a7ed2b41d042af2e6119a94465b6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97cc062cdac09b2923ef309eb30911f4371cb252ea5b1630a2ffb3deaeb96342ed7678374f6de7242f6103da43469dc86fa65bedbf97b2f603f8c365c4f74e289ce2d86dde84da7d323174e587d0858d48ed49a29fdeca6e735489730c64b58916f7a667861fa3aaad50eca804f81bcf6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h132d3685b61eec87f78a505ffd14d93fe0064ebec67cfceac07e2cdeea65f69aebe0dedf98b05a60d5457c04c66cc36a516f96e35738148c527aadead6c903f98c0d7f03808a2b75e035f43d304bcd47979b36acdc81c8d83c963facd419dc18fa326d98f2504dea0f65bc7d5b6524163;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52890b9fddc346a022549ed6d73c445b4a3c27113b42e02d8aa0c5298689a81d0c3c686cac681d29eaa7d157a600a4ffe38c82e474723040fe20d560926b93c7be491da27cadd81e06c86948d845c1da6a4fd397905e20c878eab9e19e58319a91ef37cab54077a28266f789fae0bf614;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ce3e53109c31de6276c3557eea5251d5fa9c0d99e1cfd3c6a4fa0b3878a1d709b12ae367c66368aa92168e72deeb1837a57d552a1ba39b3068355dea0ac8543a11f5b626947d804cd5a5f86c58d48649e55b7df3b1de48b91312393d85b3356d68a5335db7de075e07524eca5ceded50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedf8c83ee3165ca222f4dff756361482e6d02783c87dd23bcc1561ca2842bd09b9e3d49304bb17daa9432d4c2f33a280dde1b79f49331182cef54c4e8051696b4a4a6715ab45a5bea8e051880988e4bcc3fb6b6c06c301987266317571bde0494efe443d5c6c934244052e2e72eb9afd0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11ca7c552fe3430c243f6c7fa0c01a9db36a650338b6c750ae9d23e84bce0302cf2023f80a97a85303fe6379983c1d8635d6ea0a76b28ea9b6a3fbb781e58abaf7f4bffcae203aa19c071c1ca826b86d520ece0bbee8b4637befba0538ff1f228460a0799d39519cff1b202ccba6b33b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he78dfdb1aa1ae9bec00db0c6a47a6cd97cd3df3ab02722e955e3acafc108d9afdeb2d9bc651ee181cfd867827cea89142c175018308b15e41acf19851def1a2b56a64ce1bf46d1f1e01f54bf02918bbc7e9945ec4f031e967292160d7af97b8d95adeddbbeec4e067944f8683422f5f14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4ac9cd7da0d3863a5b617077c7c432a7be0868850a67db241a67e65daf8ffb462222334b431ec87c0ce1086ea18269420278fdb57bcc2d092383419d926e29a5d2b2cc3748a325921a00ac47ebbfad5638bd4764fe9b79bd9dc686bc97b36e8309e2e554dbca0898cb839c7e50b56989;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc89f9662352bac568e352da62787673cfa47e6aef3545c7ad08831c7bc192279356ed4f616182f5cb36805c2b9deb11cc9655c30c7ae9e3684a9396d5b69930418d5dc4863d96a76bd9f07dc1a1fc11f440a5a36acd80b999ef38e85d7f0cf60f599edf0f1a8ce5636b825f621ece094a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c30eec42f16028e98e153dc43a11c18cc72a46a861b1dc173d8fd92dc93d660278d358ae3b3f718ef23cf810ee28a428c1eddbc426e647c3cd4030296a7e03346a6e715c227ba5869ad2a5cfb2bcf93026a844f7306041ee19fdbe6b734c07bd14e2e6b81d10669c215bc390558c94b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c640962a123260834f6cc10114f37dfdd369915359d64e2ca618a820b0973517a48042c9249c7314de5b31aeb59d95a235bbc948cebe76b3594efa88802df2fc1e875aea6b19af82ada4eb70dc765f9a0c7ba5ff0e374715b84a7dcaedf6e6b84ef6b1d69a329d4251193b1e6aefee7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha573b34d4c2ac05b955e2c4f182c6cacbfe817934d8483f20643d2ad0770c3f4bb92f2e17bfbb2ee9b97f89b1c1cab1914a51e34f1673ba967a30f157bc6b697ac4bac0e943820bec68341964342ac133bb7ad316372973e926d5f9a0c59fc5b5ead18bb0e033b5ee91ff7bcdad899067;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d17a2cd15757ea4e166180407b58edbb27d476880969a6ee95e052ac769e350ca3c069d841118bc96e448697c7a05a9bfd3f9886985ff2f7ef001e2cfce64a912e53f6fd865d24d7c5fc4d5ad3a6552e8b6cb18a92b4bfbd5d08aca4df7a60a4c8bb83b87a32c92b75b2097c28c85efa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc27fa5753bff50397db3d37450cd5a1a76903370be89eb0b69237766bfa7456d45d96ec79b9b72b8a8593a1944425eb5bc7a8806a3154c498020a6c846bfe19e0b4b44f95b4aad27c13e8d3d8fd0a14692b517e9745a321bf1f2a366508aba484d4af7e53a0dc8d619bd5a41df302cba1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h248d13a3f4103afd2ccfbdd2ea71447eb8740999bf9f63e72eca5fea22d8ec9875b20806392b2df4fc7b5b1df605aa2e09525b82a1db77103120ed7645da61815f7d63d4f9ee600925cd74e2a67fa40e4e95393f2afab6323d9d1cb0c95345dd7f97b753de814216fb9b0bb4d5884d972;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb58d8aa7ccb37053fec23339b4dd9365838bb9e63e4e9e7fa78e284fb798aaba566f74168b624cd26ca7b7f543b7c80638f2c89c017d7e85e5fd10cc7d3dd82d52aa9c7ccb922dcfa447685bf2a486f6036d166dc51f8f21b96f99ba831d4111b0b548fe4439171f8507b33c724f3aa9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbc83fdb6a8dec04e62a49a96770e94d694e240090c529a84fe9e10866c810f259994c7b1264e69b9646ab769f5616e7f6100292fbdc34be5ded0ad205f315a5d14a8eb2e1a397c88f4e87a11db40b0bf12b3acd3c9a6ad1516e0c6a2a1c29ae9e7ea0f4bd8e2119686efb3d67ec27b28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ecdeed8babe417a0f7022a451fec1f6f93378254aef6f4a05fd8dc1b232065383238718208316d5e117539b939fe3d4156c81337d6ea7661bc0450349a360e664d8036b1486fde9d1423a7530640a7872529ba52d723c54ab129026c2cbcf2c495e0c08e5aec0627ae8fa3ff84c98e3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58b7bccaa12f5a29377aa327ddc3805e88983aa357145685fb8b6ed9748aa704f36d44e929bcd9b5ed214dd77b8743f3f463844629fe9aa6d5be9fcde3fe71686a889cb9b174e09c20f42efd12a361e024aa527ac5ee6b109d150ad1ae562f54da801e1891ef28e4932d2ebe8a0274f2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he196cb3f25ec06ade7a56d4fcf99b5c1bd963e5e8f93ed3d7df13af16be14b4ddee9a58be581794a1cf98eec1a84595cc75168c09ad98f62907a7292062db8b37adf035198500ba0d9cb6f5d75dde790926c703f6cf684716cf80399b2aa2f31ff8ac95ad05534db7f14d9a5e334b50a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48098dc233c028e0602d9df4042ce0d937127db1c53bfaff090f17b39cf561ee32f7a7572ce814069ec20af8f535f90942d097062d0245f06e248b1db6f60de56f09c02ec189c55d80a02616ad2b0f82d580b2a1759eed01544d0cc151b93b6ba2afa18841b885d9ab49e0c13e75ea5a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4c483a519bd8cb4cda3319c5f71aa5839fcc15a77e81b449fc0488b9c136aa63ab986365b42ca40c85a0d280804c399ce0daacb24186bbd412783497347203340c1e2c8677f3c97d7ee6928a9790de931ae0261bb3796f5a22452f91a6099dd41a39d3c23b141197499b6505c02f0826;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e08929662987334e7583231456d9caa4c4c481254c2e42bbf3aea2b1f99417e7ab1bfe8b5b56330658703f237ecd90e4a0017c956c6737a2d3148053be2160da93a1fc854c05724e11e7fc16d4dc1dfcf5057136da4779eecd6a250b58efc93af3ba6e5418b3ee45af9e96acd9b57100;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h271ec01e2ca8b0164d2c10a3a025977d0a4256fc031a57f2d9e9c522abce252887ce8ca8f5c168faa1276ab900208dbc7bdf0987614803ba2291c6c38a48c5a1ef5de1708bfc5eccc501f2a2fb02e178af0b74e599f5c271460c334ebb6cc09bb319bb5896532c779181ac7a8594e5799;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9cb591ac4bb6406c33d0d2068c89ae58679bd5a272544487adac39ce6b9ab0b168141ff3eefdd39064cbffc386eb8552ec52b28d7f4e7fb0ed7aed620b9eb500332e3ff2eff6289dfcee400978ec7ed15942af7adafa813ef7fc6f9488531a5dc7db0db44493dc04b8d1f0ce6d37601e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe8d70395dbe429ad9c4c3a1642667b9fe3101c923257a4bdc1d9ae9fe0446650ece1c62201616b881e561003b1c87b910199c98f7f090c7f1fa99c84adad8569ae1a0708fd8bfde6611e35e192d8ab81eb95969c774bddd44c323a9fc92c8f8e7f79e3602852f71310820b86e35f1b1a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4118aebf1ee3913056027e2d1eb5c013c075e7d38c8efd2387bd403956c03bbbd72addd665ecec4a714ba4a984b90c58918d0e42ac258bb7d4b6cdfb5cd5b68295ca9b23351f46d74f1d0579aaf1164f96360dcdb0ea585e8f57a6d68c6988c26f40ceeab7b3fa77bdc51b6c4a2497441;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d82577d7ff0e69f9637ec49c3022f770e7abfbb35932d967efccae60e5124be953818a120125431ff11c370c0d042da062e9bc924e11c0afbabd08ec79af6a00ad36b547660a38a768eb334f64e7aad0601e9a34b51e6768a4f523859b9e011146b6ecf6b72e5399e1182d1a60e31d93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd901a8c1e4ff2ca327651caa742d95c8c9e1fc2514f8ed82442ff0bbc6860f290fdc6d2bbca08ad9f78327dfeefd060239ead761b73d0b5c16e7dd504cc174294ac3bff723c1bd46001f17c1cdea58d34b0f1223cae0286ef355d2d4715e5a50771a117030ec88f9e25550c189e48ea6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ef2ab169df55648d1f1ccb671ca62711f62bdb4961b498235e5a9f7a67e7abe98f51ef7d96d86695d12514b4ffd26fd8e32959ad17790c96bdc78d3bf26d31add0ddc592006eee84fdd0ddece8b5cc0143708a123ee064470526761952805fc4419f6946c71ffa6b750d350749eb1460;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa0736bfb5700a5ba1aca727c0eb597f1350a5b7ed2ae6fbe909d044f5f319bd7e87b53013aae606e9a4587875a06e490de9eea49cf69238776bdb3f38f387d5adfceb1925bca4463e467de0bc9edde260f977d41ca405662bae459583af6d21d1dbf182150c9bb2b4cd17db7839b7de7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc98214aa734d259e27744f21e654d09db2e9d1d43396ea691d3b048e4c00cbcf2f7e5294524bb183c81f289d6afa3392d2de8b07dba284874d413a6c705c68e37e3109c110d3e2d17df4888dc6aa90e8a978dbbd5e78ccdbe2563d8b2bef493289bd21af9b44f9766196cd330e4944e67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd009b570db51569c08bdc557ea2a74d34e2c4fd13582420ba654ab4d478a016fed261b95688bcf084ceab469ea928903c0336a2a94ae4eb717a09759fe453185d896fdf38e2153f7e0310a7b7d5cdae1b4857ea239c75d2f3345b05e704ee11677b87f0574c10ff9adb22b3963748570;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he267908d7a99d70039a408f500545f3fb5611cecc1670e188dee531b986c0a4307d9f39ab0cd7e9d9466281569d222392e840694a23e0c62fc18fd538b650247cd5e35db015f8ade275066aa99c733d7e411894be0f569a7a254a3aa3aa48ebb3e2c841eff57ecbe7d0003317e6a0bed5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he995fff1ef9e259a5829558fdc9892fcf70177e8a245e0ea7a6565d9cc4cc17af61e6f2c0f99a93f8d5185d86ef1d8c0b327e50ff472dd7ed82be6ea3f716dcb42088291dda4c15f948e334a9b5cbfa5bb5c337d5ab3e6cd1ac49d70c54c07416c20214ffad5aa11c22f3d7cbd257b892;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50bc47ce168c6baebd0dad8946adc1572ef4e9233eca6294db041d8fec7460a5b05407b40a91801d394c093838213ea70c9887ac392b5452731223bcbf474d50a146f35e9cf9cb31812537018c97958a7d2fa31110c0ccafbfc54e008a89c2d97d64b8240a132de84b106825286c8c86f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf1517277fbbbcd3eb9ada3d36f207a2f4fa812fb461ab19aae7a196ce981fda6b338350bf63a3f1fa7b99de34301269d457851085f2a69da38a40f6f3711e6cf64a718d052e7829b5689fb6f0773a67b07275d45f7d5ab8bdba3c9682b85790407d0cbbf10bbf73922656db4a16eda89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdea5be73632beb59d4edf1c3044af1256e126309636aefd05b4922614445bca2677685a1ff92ea5d82c8080e19bd0a2696efbca3f823b1a2e9501eedf866c4750d535a06b128051731eb64ec7ec8810a69e216bd0a99154ec57798baaeebea93108e8d37c9b305f3bfb65d085eace54f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81190e1d309aae40852cd1aa16d53cb2d5753bfb7399d7ca658040b5a5022e5915ec879a2ae8243ad1495c612cd7a20ff586e832ceb054dce4400894d9895d0cdd54b26946f54e7e06dcd3b1da9b2fa0cc3ee07f276fca2e1165a70d56cc16721aad9d732f7d4e84055d313c8f26acda9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h972ec5da2f9c5c7dd563a9050b15e94631b94e411ecaeba22e2d6952567281e70389f46b79b4db522c1afc4a66d0f17fbeb183c7382aab5201307f18dd3f161b5fbdb28df8b8f2063282ed951e9a303f3b8387eeaf7aec8fc56a3e5335add081fa8e03ad0b7e52d49f1ab8d55f08040f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fb489a4425e748881eded2cb37db0981bf9922b4cc3a042763b11cdeea4ae1930b8253d4c7abce8851fdfab5ff55bacf9f77ae3ca763a4b73dd38088ad8b0a845017dfcb25c3bdce91de97c223f334c4818d7176ef62b185ca1f0bc53d2fc9eb601e27269c5f7752ea1bee2e91be7cdc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h435f9b18491f7f3005c2d267034b1e914a3d9bf77ead71807464242de0d14380867cf9fce4b2cc0ff2fc2fdc8b1cfed49ffe18a9b5af9449490a0d7efb9d27eb5b9b383f196c27281948e50f703e8e90e3f10418654c28004e2ba0d96a95ec90f280a2918444f673a6b748e21c3d6ae0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64871745c27655ed51a452d62d583e5224435392ed59a3712503d47e5b495887b5f75f56487214f8d30a729a8b23d510cd5942fd148cb3f4d7723e93c22d7f01a313a2d0b96846ac3d140818423a4162205880e677384c49ee4a12aff612377acf26168b9ef3f1a7d0b6a077943bbc691;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd16c1ca5387c120a9202c10dc728fbd701e942d9d7236348f493d57b71d9a13500dc6be81355a07c1677e664e1b5b089e858b17cc42c32fb6db6f2556bc1717f98f06b0886332f34c45116e6ad86f6bf9a00e60cfb25cd0fb366196a20606881a0c83ec4e7eff0dee1fdca09defa1f6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf86b96c59a92d67ec6a3e4c00a7715cb091e7950c74f468ada1e31aeb4cbb2844eb45dc9fd09c247477d7fec29d39c7cf71b5c50d3f10d71f94c7586ba5be1cbe44424071635091ed5f52822e514dd324c8dca9041bf7379cc6898af13fff179c43f3d6daa02c76772ce6b9ff671a1d60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h483c1191dee51f4bc99029344ee9ca64712576a2474388732d320f05e5d375da39b3c7ca32f044d2a15dfe26aa0fbdab62b349d7fb1f2b4dc9d53f43aeca5b7331424c70b2834603e140e803515d78560d4982fd4164db0f29b63275b955554a4388f384ad6940b942a25d486208141df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c03a584d71c356a8ddb698d1da7e7af37479c182d3aaa1f3e9e6aaf51c37f6a4c49d5a37ac2b70017b9c8cfeeb88dbacf01f4b78269d716fbee46faec691c6a66137ab2dbaa557b6cd56a953b0a1564ab314e32dea4904ff500b54db25e04ee565b700c3b69e7b5ae080ae1bc9011ae0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81656f1c73cf39ea86f5f3233dac2d47aeadf6fea07c5b6afa87defb25d359b49d431c2f6dae5b25dd8a52e7c9bf7d9bb26a0512f313477c8979447298ec3cf66d14414841d5bcf8df4db129d6c359199f98b490c89b951d52361369f93a3b1306a28407ea50a45aa8696f1ba15db2619;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfba4d1ed875b2dc5d51e7b20d951a181d17fab3d163e793bf96bd96521a1762b9a0e1f18113d15fa6d912e355f3a290fab6ef7ec76987f313a241f0dac1d9b3e4e32f00d612cd2aabec7776649ace433df97f5ccbf0213f38ac7c3a814de6d89ff96f4585b8d4f00556b36d35eb61dfef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecba4730a7a4614cadff654eaf728fac47518fc304badf7b5161c2847fb515903724dd7ef58d388608df9ec4fbb877923e6980436cbd6ceac078c66b6b8e45c6cb2c792dbad760bcb5228d4f5bb7a905f5def0d8a0f56363c79a3e62e029db918c59d55256f3e4e6a8300d9f4cb870f5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dd3e0a30de87f9494470a1babc6a027d51b3e889d30e54f48486f5d7e2f52933294e3fbe0421bae6a24104d83d0a74ce41d612ff46391f9975f25dd9fa15d057e16f3924b137b19ba7652de55e9e15bef8a4ccbf0a4e5b7eac40baca0e462231bf806649e1ab71c1f84f299fc48adeb8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9913bb9073e6947c0569ebcaa2d22d944b7a8b1b27a08fe647578d6dd536a8e4f9d2b3c2d4e3ca4d97963d4206fdc542d02e99cfa0fc69bfef9fd6d8a254b8179136bd5b14dfc48473ecaf769801ba05f1d73607ce2bbca55b88983f820cab5bc951fc55bf89c954a68d1b5d01550553c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cc034715fdb9386fe1542a43624a96d62072347f3e6ce3c75def003dfafde896beea93c5ea0ca38fbb800c8025e81e132bc491ae0640382bdd3d6cb3b72ceb047ba77660a44e54425ca4fb439960593ace1f5796c30086434334db7457d3a0eb82e84ae58a00fdc45f0af0e377972a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5788d1faa112e710f6fa0aa34242abc0b62ecc114cb37a1889f02d9b7337936d6870e81bb0cc600e992a2af98e11e86394f1d027ffb7c301ad062e8ee7422fedfb875b2aca803fce5e82c546f4b5e4b6922f62e6c74c3aae6db0cc63ea2ee9c7065d530c3c89d65dfc46f008ad921fec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h544f70e7faaa64fcc1c70a63517528131acd9de57c347b1df5a1f9ad45ff062a6cdddcc405f9ecce2e5c29992a70c8a996f3c602286bb8dd9234a63c88e54f94dcad244ab3eb0edf154bad41d60c7cf87890e166a202abc1fd6e8bc3f8226a2b5ea57bb55dd9d4eacad68c09305c29fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc03f088884f956090afe69a89c76757f40229e73a990bf00ccfda62e7941c100537263924bebe753500d3f78b53ae00fb634f9664e80b7775f7511d4fc073bfbad66c1fb00654794c383535b58dcbc77f4e90a0555d514912ae8b57f924f5c4e717cf8f9c8d2c2ec8a4ea2568a71826f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc34931e2d74613364ec090255feaf2df3ddb72d8c16ee0e0f8dd8bae624f444077401b91482b601a590e05e5ace91595ddc9c3d6fab773b14bfa630f3990fabd34a5fe0da22cde26fe23865c8509b864774e943f462f1f6141ea441a8091081c6de14ae9aacc8a68dd64fe0a5bd346abf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7481e0fbda457260d6a0a2f1aa745aec778a30cd54d5fb37ac296dc13d91114f52baf8e598ebe9e1a44839b52d49e89ce0f9752e2f2cdb0dd402ccbfe102f0d3f4c9014ff0a3c2bc23dadefc580da7825cbfea04b82a9c05732724ab91b8598f9a245f71eafe77cd3b78f9ec63a683ed6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2083ef30786ffc00397ed3cc35437eccf26224709915aa501ff6b76efda321e87b27aae6289c81e181ff6b9dcf8ab425bf12ec413ce2b69bc181ff62f18babf125fce025005c8f4f69f0f4cfa35a245c56fa9afaa7129a9f354b0ea8728e8ab71df28fd0938d3a82392d8a44bb40841b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb97ddb1dbcc63475ed36636e439c08e707792cc67a7d23cf8c82a77a8dc6f7e36f4ccb551c19718f43b1c8f80e25bca6d4854b7d457676e7ab69e3a8d734c40b7646e4cd63c794f73b23a0327d554ac24ae818503a22cc893566d27d904fb25661016d8eebe2f112a39aa4d391d352f10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82b6046e842f98ba3c35735806f47ae8e4f91afa0203ad0c34fe586f9635e86dda00a01ca4ef0f662d5abb0749ad2bdd1547852c86c4684285d8c2f7a9454c584464bf20648f8ef53727eb8cc7ea763322ce4b650cd412ab17dd4f577853c0f3016f863e5720731706eac97ca364e4410;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae1967aa369056e47b066a5163261d4e65fbea7ff43c57e7d6d18fe77474dd4b7bb0ad66a81cf699f606881d732178b5b4e502004c35a92a64b13f6a91a4504ecb36676b0dbd9dc2c604921575412cd0c844b09e8c55da5dc8c7a8b46b5268f68190ba8db811f9b54c982e95869f647c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9329de0434c2f0a31f822a4bce35ef5cc5c06402e3b18deeb1849c977e36cc45eb82d75a42403ad8f83685483261e6c4437d65e450b556554d346b60c94b6f8735c62b41d1f4f8e589f5ac7da0bcac0a1146f74b56cdf8c2616c319739396d923c7e1dd222e8339c4030fe9bcb4abf344;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4690896dd1fd4ae8aec6c233410796d1353b36196c98b14569fb7e6ec5b3cf224702146fb0a2d5f1d2914c40b7cb47b95b8f46d14b97e8d02a4e46efacad99a39af5302f0f1a0295fd7bcaf2dac17ac47da6582223f6070e837b755ea160247b0d938d1a1db5ffeeb62444849374e5de4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba879bab2de1e862a51684a7f7c4e0ddc364bc4e8c4db5ffc548feabfd4c48cc39774a5f3edbf29c9971fe3732e311e94ea58ad331eec1de41b73845617a8d14513cc031c6bb1982a43ce1c00e7b786bda60d43e830897ade69cfafde7393d67b02569c0ff974915a9965a4c9b529deb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h332b3f4fae17e5183c3c9f486965fc2b50c2aef308e4b913f71b1cbca0777dcb1276e48aa843d84d58bb5f7ebd20ce35d93dfa968eab10331f99311da1f21c62dfd893a8cbacf99680e7ffebffc2b62ac06497cf5af74ee3e3bf0325d2643cb8dbbba180cd8f4199f5902125b5d76899d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26bfad330982dd7e491a3fbfeb703e265a2e83c94ca8039d6059158049dda2d79d6cde1410881a44f28d832bcf350179d1707278bbd0abf58234e2a805249a8fe5eedd5f37201a3b5ae9723c4449edb10b5e2ba7a16a92a2844fa6e57141e28a9aa18d354e43c7c71d8dddf421684f591;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71ff7a63f15cac880b8d6e3f335cf6b4fe76f1fdb99b748883632921a1b9c9fcc606fb18bd2e94a60d780be18343e0f5b04fde6061ea9222e2366218a5409dbcd9ac78cee32c106c177c4aa5bc7d4223e1ef0e979bc8a55b83564560d34df388cda8559b4964b2eafde01bc938c8ff6d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79fbfdb5b7f5f670f3afcd3ab57a785752cfa7b255344dd6e1cf5581d2dbfeab2a4064eae892bfe1eec7c46f86e5a96fb2f056b410bca41f1c043ce9a2993ca871bc53f754d682fbdcd13a236c025b1aeec138949e0e039a7c64fd74576a6bba8c1b6de9de7008775d651e754b3f9246c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0451e39dd8633bec22624ff804219c8c44ccf789e1d93c73ae52c5687206235da8b5d6bdbe7dfcde7bb4b0ac6dfef8e842d64ef5502f645d75949a7dd051ce2d000e9f253b0b700c2f378cbe579dd71440f77901c8a1c846dc9ddffc33e3d701ce64dc4def2f7411296000d1b2145945;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he02081f01f7cda47b6c091c68113e1b45250365c88d0712d0efd1003b10334d06cb9e1f1ec1ec043094d98ea8c3059f6a65249b317929246ad37cdb333d29559dd6f5dd7827298005a752ea8c40baa6436c575e2f7761844b46ad3386d2030771c1d93c92a0dab3c4d5fb89810a6f61f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17da0b99b87d437bd2d77116895094e68925163509785b691668892c7757614f96137fd506d3341a85d7cd90d2fcf4b2252d38b1989db21d8f000a9c9c61519c67e0c6929a0eec43fe6966ffdcb0660ec2f62209df6b70946d7f3072440103211692fec8d7f86999f510baf760e5d4bfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9547707ed63a88238963ea05f7b7beea781f21351a9ff75dbde3839f38ad15fc2ab79358cef282af7d8f9e5fa6aec8d8775396cf1362b62e77e507bfda1bf0a8ba34a5bfef026b1decf86257be2ce89e0093e637abeeb6fcc2bc14d693e7b8ddb418199e0b3ac0c1764e1f47092b01b7e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h126e269281010108f9ffe9ed0bf6727c44e83396a4f0959a8c313781b2ddaa3d4d1bdb5c44a0b7169062627bc3c19b4fba253e8e1f5a7336e4a9a1264fa9e2a755ab4a3304293cc9d6b0a3e0ccd568dd1e9535b9c61ca177a7bb3beb4e93c586ab0a1861350f421ffb12172e77c81e4f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb923eb54ed8783ea9e421c7cd166735ae158bd0138d9727cbcbeb8e53e16ec18877d339c288d2b2a67d3c3c610fc22088dc2b07e58d7e4ce6c2c552a3a08b8d60403659aa3f8f62b60766e3239fd0f28f1b91defd04c60a08a5005398a2b88f1b8eeb06c5be16c712f0dac11afd891f88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c52db5babca9d2acee612ae402453c6e30a94dc8c4a5340b0520e0a1c2fddd0a57ee0b5f0357f221318cf068737c96306342785ee71f5d22245b46a26c0d9d57b3a55824b86c2c449f4a4282583a50858a614d31307a93c8ec27c365093c430008dbe2163e855795765806b497e11a7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72dff4f03dd1f69865cb1ab45346d1afed67a190d056d19895757204dcdab5de96085eefd59f76505a9c265a6ddfb0c84504634a255c644c7cad30ea115fe7c4abb4ced9b0e8b692b36032318413b174728408e5f83ff378f7e1e4621aaf137c9da8f89488d8491da2e7977405f08693f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcac93e93a25596d96308611bcd6a3650fbe16d56ee575865481dcca520661d3666ac58fed1422fc52e873472c8f3a7c2bdc6324853ac5f608b823afec488056f1eedb710f918628aea00d58f07330f267a0505ad4637adeb728aa46114db0610a03f85c793c065da3fa59fb684fed5d43;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8859022d0166341ad8d81f0be727522dea569f1681dccacdfee723ce00af059f0cc45b13299f0a491911e255ea849ffbe4691b4b41b16cbb13f24b6163445a964e34d31e6e0586802ca3104f2c819eaca063b80b861e5ce149ccd1dae5e82e77fc131854e7150be321211aa2041bfcf2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h549967b11027fcf6f7f1005f6fb5b6a74037ea4c6ba49439aaee3c466cd46381fbd72e0f40cb11833b3971cf5b6028d2a4822a326e5ec92ce6f3c5fb0556c64c65442548d6cd1f1ddc58d300ba95f18a56269c59ea5924dbc9862ecb82a2ea106c6613edad36735b7e599446412bdaa3c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f47a2bb6494740dce62251a5ef69e5b5b4d09b6519ac8253531aee467f42c5fe3054830c8a4b306382cf50abe82a7f133545e84ff1b9030d79384b05a42fce48cc6f89c3151ef12f09567bfb752186c4c90aaa9cef8a1f96f8f93db5e975d4ceea1fb8371ad5f7196c62788cab27e7e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb299914c3d168d2ac048858a7a2c3848e652f041a8d75b26298aa101a3f4df9736d646775a7b837874c1b217607cbbaa555708909eaa581002f0fbfc1ded86c5ff38da325bb069d9d0edfc66ec30fd64fbdbbb7c3da693c0b7b53e5a7976668e311ac545b21a03044c23645354c788737;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd84f0671f9b5ed09475a01e0a95211cf2d03f525a666288fbc1aadf00f302021c5a20ac01c6f0fc2c0aac05d320796339721e37d72ab84144ebe6219d5dbf4f9921e1bee34894902736a713c678eb181ec24e317921c7c9af16302938378f47286254dfc0adc91c93e6680f7b1d05f979;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2f3d6cd706f11bb0fd3d435518c00942b73a10211f39c5b183762fc93d7752eb8126b0c710766d1fea6fae4e61e99dc52f32735c66755e5e13a47c91a37c0b46e9fc0df8319fe6686234fa1a2695fa2c21e4764e47960801c8bd47290eb3f5a91cbdfaf105e31714d76a056852f7f949;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88bb5063208cfcd663d2d23624c8421ad3a87b9edd4f635e894a9bfebeb48ee6abdc7f8721f89af292d0c600478594054a994c7dda177daf8c9614d7c8f1a47967342534c3fde0af7830a6ba64e83e30ee16eb7e4dd8ee95d34b650dd15c8f4c975dc6fce79136d89ff164e462575d7ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7df617e3d9df2a1b9a281d31eb511809f6aa7722eb623c71f699f9605f1a162c64498589edcd419959ec0302e5fa372ce9fc542ce4d44641a350eb098485f2ae0b40de710de9a767f3138d9962f2bd978b2594d5b2df93e3b3220e21c695113db3faddf60ad4f89f7ee80e019240a3bd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2ac967980238a56960f5c298e116d25b02dbfb0744d855ab3dfbeae6b448be2a85ff1e72f772841d297be57870bc6768f11924e1df7a8cdb33fc6e2a348fa7f2e6fabe179d290a1e1793855d3f6aad66bfa11587a978e42ce44380d175d82216c43b21dbc28698d9772052179e5aed9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h359bf76de8128a217b4466e9cacd4cdd8d6605f215905ec3868936d3d06987baa183134a54aa0761d8a987829bc459d918c1c22ecee810a31e564c855e056da0039d986bd873949451aa821656ee533f5e247329ee3d2e87f072d0666b1981bc8eb9d19107587374e4611a2a0ca90342e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9fd87f31c0bb976848d52aaeb89b0407b9fbbb6b4633c4b23a195b87aa552fc6e471ff466db8fc7b8169528999296ef0380aad41dfd3d9de41146805aca8d88f11609931ec506dacbc58cb2cef9ecf6fcae8d217055fa676ffaaa48c2d5d760652c4ba0beab2414b63fc3e928650e014;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32198126ff6783e23d946411342ee4217dc511f825ebaacfe3a0a97e203ee6d2b4e02b4801bd9f318ebd73d2742ab0cd4b7f37b53de522fb277e74c6a39e4012c2c1f89937e091f83ecef1789326d8f02fe91a6d2b57b3b345a590353a54e68bfc692e107530256ec86100332f6cf1d25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9376916779e6b678acd2bd3184b3d4bd62e8f00b2d855bf4dbd2937edff82e882776021c84eff8609f37704cc3d35f895c9f41a2aac9496e7933a7b76e34d0c1997263da0725f64fe4e0c6776fb52ec6782ad56409002b35321c02d3e60bb3b73dc35a5ce033d084792f7827db860a2ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc02c2eee5f59499ab28e636d365d859ef669a20cafb5854f3f4f1888488ef799601cebe5decbeaa835d1277c15fb7322ac56821f770fb4167383be83a94555b984550fa2f9108264648100f828034827415567c63f80e79db6c3c39ef87ce3ffdbca56aa46f41b483a5f33efea8edc56c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c6329226c6c357d2b0a237c860910c69fd34f2aa1fa95aea156b6567f12cafa48fb337b93f192e4cc3ecd6c15adda720087573e9bc33ec6432e40d9a11d0cb11f0f4b0fdce74513c2118a1903876125d012e057a2544a71f69b6e8fdba6cb2699c330a21ba0b16c7c1e38dd555cf840e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14ccfb6039e411c2815ad57a950e4ece099ab4565216e0d873f4c1fcfdfdf16b25282aadf87347bcc3e9cf0173d0f81cb9e333bce23afab04568b7183fe12878044726efec9fd2a19833ae7865284b7b8009633ba7184e7cf8d0beaf1282a248a52fee62dd6980ecbfce886464f24dba5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5e725351def940eea71a652b77bed461ae17f1980132331d232b3e3c5ba61e6da088b4877704d218d87b7fab63d5658d7eb22560c5fc5b56c8ed7b48e190c32769ef5c919d54264f085429a589c94dbca4e58f9802de61909214d13bda8ff9f46e02fee2375c3a3a7653461808938354;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bc3409bafab83fe748e1dbdfd8c7974230fa8eabb9bdadb8721fbf67e683170f0a5f48daee6e60353b88b1e0f78dbe248e7926a704dc3ac2561dab41a8db745fca48fe42a9699c3daccc01c4ad344d95ca139669d11bcc08fe7dbad44947ed784e416ae01388dbe771b0fece25565bee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0c160aa80cda609164f596143beaee46b5037f456ebe3bb9c0267a3fcd0bdc4ca7531b9b0481c53123cdc1140a54ae5e94f694eadc257ffaf702aceb4232157d015473b084a5eb0a024bb3027310063d403845ac2f26a7f7f9e60b277582055efd1345e95c676bdcc3e295cfd6d45087;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h465a1d13f4df4bab91be9ad473e417d00ec8439d3f44d3b38caf6a75a4883201703e302c2409bc82bb063dbbaa048882ea0e93a2565627d92e9131d266b50aced7051b55d34a9ba91c7a01c26b8fa070266ee7adc205a41617f381b5a15f642e5489b3cec40ba2344800bbac26b36319a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48caaf9bad896d460b67b93f3742888f47309c59463eb92ed9c95a9753b1d23d2fd57b8ba806df245ad16d7132b5f2c597612dc8b65053f8e50d59073c593149f5572c76f351dc9601de321a41d547c04c2630ea0446cffa0467acb8ab798f4552d7b34ab952dda3d9792c1980af1f218;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2baacd97ea27d4b04bc7d7502d75ede3a5581f66b83e58f353521205c9b73a0f82c6a277118bc2550ee7bb4a04c4010c363f36a20c8a2e7f1498fd110fc985ea92493e505531733a9fc8fd1fada8c99dd70339b4b614ee8b810b50ed725df253436776f19329ba767fe5a6384b179c4c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f17b20621b80dd947e3234f3015425fa4efa7616a35789a92704aa7a31b52a97f2482169c62d41f58c6cd800c9150563a9b9f39732b2c7ba08759f9c1c42e5b2a8f7e51f682098c4e20ef8b89355dcdfcb4c91148a7a140633690f60cf423ad6a990d65400d7d015a02447d1520b5b3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb21fb61daab5070a27c637cceb4dd40016b6c0c92ff4b1f508b89baac88a91ba12cf334364f2f1b1735ff6fa85559c95c71cd9ff867b05464ebabc1daef2dbd6d831a3836a1faf2b1b71d82053a3ea673f0e814b5ce694369ec84c1a82100dcaaa342d67a1976f0a99b468e3f141dd77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b4b5903dca3b57a5900ab7343e5a9db951d0d0a1d08ca0fda99952a3cc3514f5aece57ab2649bdea0d9fc1e86354cdfe55924b12065fc5420796d3e5ad0cbae62093ae5afcd8f0d9513d6defefe069c85903e3e4d693a53cc4225dbaccb49cdba4cf1753fe02728f25c169b8609dfc01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he080541393d341f9c46fba7e2894e2b331ec3193cca71829f4158a1b35ff5d0b9ee721fa213a03a750487451409b7fc2c9f5fed3f2ce5b6e4ec5f49d64409fc991dbacf90ee2775a470e2bb58d1f6b73e3aa17cb6eb58a330da17371799ca1f482884ff169c027b406b01175cfdbd9410;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0cbc5dada25727c45262b84a46dc555842f193e5c5e0c24af22fe59f91303b6e712ed855b864eb12e9ef89f13a184cbae13e2bc9706bb47f6436a1dba8b2f3871a0eb1d242e58155a4b42a94cb0b2a94de49be86b467d2fc40ca16944088ce4104a3fe1a4fff52e59f12db6704df651c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haeafd504d648568ac4da1ef1f6f339ec34b0d9fa30dc4862a35f04159d9bbc1826ca20c68326e21a394080dbea2e10c467e880b40422fae423d983081e6b1d78e2f3a7bd18c6153b9d660107ae14edf6c7c296c6bf998ff0946cf8f524029de54d9a368b7f9ce64f646a74495384d3331;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec984e3018c1b0d0122431358114486fc9b5154b35cf0b29a326420a089aca445a72a0d48e3c0b0d552f2a51a03a914f3b2fa3a5b934d98e28365383361a258ea16ff3ed1c4478ad49e40dad847f786b7578bf059ff93a5788044674c18d366f941296c2d06e7bee5adf6c774c3d0c561;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha181ce22674edf39b5ac774df7249db0f72ed8260fef8df0f2a43ee2c8372d6d0149e413f8f5e0db3ee5128ce7463b9bb5e5945c25962b0db40ab89d5be839b654de5bc3b004951376d7ed883f453b883eda592913592741f3b293333d876921c4a6323f5bee7535d8705166a79f69046;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93f65514caedbeb53545d299e9b656b173f6ee37a63fb68bb77bfc01eb5524dfacb810caf0b3b40be021ab3249bae9213cc0fc6dc54119bdc54075f17c43e22f120f74835d05034099989ae006bc89b6485f16408425708a23446d2601eb5eb9ee931ef711e63966bdbae201a44b91009;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb49b1083d41dd7130bfafbfb42ec57d419e737a820c41efc9b8cc855587c99f6cae01b6b1a06ba51b00e54e982940e7aeebc6beab79f933fc12622c2f935c497c70274735ea4d8ad7638bf33a7001464dc0a56ca887ecf81ce5a4a6aef08d98ceb44e83c688b8c5ba8d7eeb2153b68f42;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68e97a03ad1b471666c4bd77c0d126f5995f2d6ae86072daf932472c894aa2b685269d909e4c56812cb49dccacdd7bec125965341f31a9ef1dbec7c2302fca0643b60e151b0b48ded1f4f8abf7cf0b05f00099771310727fdc93696a453cc8d5228ac93f09179e26c02888ca23072f229;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48feab6149752080df42a199b9b5d8ce88d1a87ea6e4e1c8f30e14b1a931f042753eaa2163aaeca3eb75f790075ba854f48a7f06be66a9defcb0260e97cb9a99a4462edbe7fa3cada1575b460b84a6c59742b50a78a82c255fc25531ef23f06cd27e906d8aecdbfddc13b24d52ad86395;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h294867f39102aac315c7d48d3ac41d6338255f7acf2bd230d82cb6269468862a68fd6ac273b836e3684220fe89cc1925d06e35b9a920a74598764e49679b7e73ada97e2f01d738b20852302c9ac31fc5b48c757c6dd1f8122186a172938ca730495a80f1318d0e60488066b3985ee1355;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2d7ae649d8401b800e767f7a1ea1855b95b335b068aa217d5a929f2e022fd719636d66bbc847df6278626eebba1b9ad33f89d3676ff25b66cb463f896f8a41f0f31e0d4fad484a39e0b47c98bccfdaaee016b942371ea4e4f1d09e9b43839c42c0879c50d14e23496eccd00f4f56fa22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10b01597d8e8aeb80a92793a9172fa1c36c16ae68656696de5521fd42f25051fbe7a096ee59bb007693f34e74d862ca786352a58914c17d3c9dd6ee47de02ff9eccf8f53d05410b67bb632c58da4e7eb2d77c240efb3a1bd1ab8c852d6010a4840bee28ed1be3997eb30313aea4cc42c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a94b2c39d85040f39215e52b816866437e626e3212fb98694906795ae2848a8f17bcb04e2d25a98ded5ed10097cbfa81b8c3f43983520cb8505756dbc59836b3dc79b0f0d77d88ec96e26426ef064aabca24cf56ce2ff1c093fa65bbf79c5773121adee34a9a8cca2b285adfcf193a7a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7e506b013019427f1cc899afc5c7aa10ca1f05a05dec325a04a1b67db64788ab854408d9cd2dfe9ccf39861ca3cade214f451429c6e65f22499b90848d0a0b9d8e7ebf949e2d4fefed888027be70898e13285244802c7bb0ffdf68d41b2d2f21a0e52c7032898ba1114a1a8292b9b7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a60f6b4ce7b6b6ae1fe315653a9d5af0917e3b50bd9ef017e693dcf91b02c22210f59a9407c21203b8a171447419b58e877c1d8253d15d80c7a3ef18a7ca3f9f203beab8a6ebe048401497d8178069f664789f7cf2a8b3b95ecf86f1dfa0e5e710aacaa2f0b1de75811bca8227138401;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbeff5205d895ba2a8b8ea8bcbd90eb17e8dbaed29361eafff301480012eb260a9e49047c2712edf530f85a459bad860cbb5b6e7fe9a4e348843b890ab9918d2bb798adc625a5ab0917a479e904ffbd2af4f26d4ac1225fbc6389e98e7ac2b9109c8a42af1c4c6fc9939e06e267860ad7e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h659640594a872fde8ac72aacc0ae5b888b6dfd4f2be00d8c22c7936304cf4a571303e6653b49533e69789eead937b6b5d5f9005316dbecb7a105da1ef1fc02628a5f71b72a6aeebd331f92658c590bc0aa7564e6724fe46a357b3923b8f037d8b57ea0800e62ffba07634ca25b9770946;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14ef20cfa060b03ccaa3c880ed17eca033f359b93300ffcd176a3448a1d14742865e73a4a2f3781251916775a5c5960f371c1645096d85af3f2cd65e025d4ac67d308ff1fcf16ce5e01f180facae436e7328cd8fc83eb58eb2f28445affb2aba2cb60c0b7c05c2572f3558ff9a2ce638a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d4ba4f87eea3cea136c78f3d3667cbecdfe891e7cb34cfbea972837099405e2a9bdd3e6ff0475fd4c8dae4bfc064594adaa03e5d2478353f6cd57f80f0d57c92dffddefa5fc87705310455c87e240383e0385dded607e9e571eb006149de3512a481690fb1595d5f1af32bd3970c5131;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde260547eacba58239c325525812bc6d1c0b9a6e149e90397a2fbd9c115ea5740aba824e53ee1498498699d4a79bced70c6b8f05f210a78005e91a5b83afffde1b2d573b782d8c4287bbdc4f88c263b0a517ac3bcac043cf8bc1c7f26f4aa83e0decd980a8db2beb39485f8d7d648dc6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc18969398cc7443712d55df7d1b74b176701a01bb761ce8a8ac74e733049c041e5c1c0a9d6b61b00ded36eae2fbc6bec9f508e4163358d69f3085cde0b05df13245028fcdab10817b1370b3a53b3bbc920daadf46a7fb0ed4ac30d928db67869de149afb57f5bbe00844ef2abe0f02118;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c2be97267457bfddbb7cb94dfc67ac4a98714ca241b4424817021a210707126c546197e85dadd368c2773f755ba2d3a4f05f1c374bb804e5925638ae8d1e0c031a6203116953a4293aa4f1d49713a857391425f767c92bf1744b5052dab8581de43375b8fb1d6bcf56412c2ac8a56385;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4645caa67d7f8a052cc6e6f557fa4af914198403198dce1b118038879f2d6a0cc11d637cc370b3dfd7bde15ee818fe005ad852c76fc2b80735d58e9061ada1ec0649394db0ec266bdf3f238197a24441e887a8762defa4f75c8c8c28d3665d2d277ceb715da508141a9327e6553599456;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99c5502dfcc8176ac641cfd58dcba923e8eacd357279732cbed7312dcff122472517daf5c39dcb2bd80b75280a91e08e6483b46551d0bcd1050a0bbfa5f8ea4a6b3a0e41bc791555f50992ff4bfc1aa84b43639d9f45fe09370e38af58d62becc138cadabd64a04d7fdec946fbe99c3b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd306b75975e77b8a8d0a0017255fd89596babc9704db9c9358bbda605b58713184d91970f8104d5fbe8abc4c3f1a935e5f38ed4985c0ecd8642ce33ad2e283fd8a700ff4798165ef5cc87a71ae1334ada0ec6025143dcd6e464365d5d117548fa7bfc3d957272f47d7eae17bea748ad5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2bc248ce04f4eb86467833d73f96b57a2641ba15b3918a7cb4a79b1bbcb2f5d2e1bb31a248d972653e970b1a63af93470952dcd12b862ddf719dad05b2ae168e47ab1adefa474d6ab38d19c3c7944fa1adee3b56310ce8f21a445fdf33d9158d4d9fdccfc83ac605afec1f4c6c92776e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h140de3dea386c1ce9357f697d70467e475c0dbc6299cc75bf84ac23f3f81410ea9b022e2471c1d9e3b208e40ee12d097cc50771300e82b52b64966bfb9b71d49eee22255e6dd95887accf7ba736be7ceffa0a7f4532de5d773fc5b912253c242ca92cb7ceda7bb896691116297ec01af8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e6bc376293c1f41b474724f86085ea621fa6595289ef111ad6fa58cd450d08b6072f3cb10396979a78d8747ffc74fb61663dfac422af5f21cf571b141f89b8ad8483d30dc4944842372c5162d1a5935c51f0ddc9a4117e2a148534e4b3d4149c40891dc1e3c830bf47dfd7b05a7da5f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fe2ad06465fd4bc777644d5052452a802ff6c6f9338f4411c7e7dec094096c6ab277b75abb08982e8150be336d732194afb332e46ff169cd6f8feabd12893f22ceff0e262de3d79ec88e76cdc46e99a843714596c22d2f3fe01009cb84d12322b207539a4d33dca5b70e9a3fea5a7ee9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef91875081d6fd2d5b9df99b5c82ba653404adf9902c9da497efa1e9c68c2eba0dbd08a943000998382902ca9e788998137328dfb0cb2fd1d362c54e21d69950a4da9c3efcc64e0478fe88b31a3a925a8d8f6ad577ec6e6610fd174b7f67ffc1aa8fe5fa3b22cfb93849d2fd58e69fec4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a90f6594f4f3a19346ba5a5dd037e2a6c952d7844576fe6641d088208193094746f430236835eacbb9153d7edf9b46cc03006bf0137490ac89c8a0ccce0476e24b91352979aa6af32b59984c61c53204b609f4e18655e854e315e45b1bd8a305480129a8cbade74b889194e54828b8c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17075bda9adc6b2270b6201996e4e46bfee786144563c669d477e19da99531090153b835a6b93724fef6a04f3373ac12f488443daa56445f9006af8e1385e0584bb3c7ad31b3fb1a5d3d70c980019cfb862914cea5ce0a82a96a94d611290c622d516f82d8eb499d0e9165ac074fd869f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab4b9cf194dc0bea626b8b05095896d77f33860e078da99470d3bc99ec9183221863631deba174f5b9b59c722699fbe29cb840bcd8b9f9e3893ec6de0844658d8df879ea20fad9b030e024ef1d2bcc0004d9f7e35c0c764a0f9d71c14ab8e469b6c26225f1abcd401518739e3683d2a04;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6b4bf836b79129c9c6644ead8c8723a3e85d2cb5d838459e464ac1a38c9b0f27fac351c5f7d4cadc06e695174c550209b7b2872cecaf9c89afaf6906e82f54df059025ba8d4b03dd62612a91c66650ecd5816d31d1942b1ee6be4b19f24a02fe3abcafd8b7c418be2805258f9310c56b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h609cb894b2aea1cdd85f6522825f9c87fd5821bca70c52df656e5a081d66a917b7d2bdf2f9f96cde33ba8b51c88386c9b9e4797b11ef5b5c4f33bf35bad99cf8f23d345f98dbbe19be965ea4ffabad177f501f9ae0a2e2dc93ac618006351840f3e4421a4aef158c1320ac01bf354b95e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc854fb588c09d4ab18e3ad7d987a2fe9cc8119490767eb931392553abeeee815758e2657ea57f7ebdba11612d2a7874ac93b0956b802a63293bb6c08f2aa2762f6678e086a174167e640584434a56479e8c9970531bc1b2c9cac15e2441e51566343ab1f079960f6d7fbc80ef97390434;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h805e5b8a469a847d37742e2a82e24df3d63f0b0ded313936b4cd17ce5fdcefc68a9ca7e2e22c34e13627777dc8333535ea281f72878d330934e46111466e8a6326bb8663fbec3bf230f578820fc83033a9304bd17ee77625d37697e8f6d47ae9bbe5a05386e247890b7df33ba92d1cef0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa91cbe3eaeca04dc995ed159199034d5a36e4f248b76fc2ca2cfa70ab8e88ca5daaecd1ca83c6f7ece385ad64f683f7fe8b0aecda97943dce20c1af5563f80611845605aa12624a330f5d14baec03b5695a5c42653041bbf59d456ffc8750c7176a131b601b140398fbd2cacf169dc79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa5851b5993ef6bf58cdc82d1827a18b73bacebfac4b0f30a05e6ac19a3883ed318b28aa7ff6a219b8461299c2d11793418b9ca7bfb71d339abf4a544be72c04d96bc88d320a24907d20b5f2e0d6b19842e71b23fc08e7a47554c5d3bc8d805aa87f5f385a37f01ee0685640862080f2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf383ecc19b4bb8e2ab5d7771e45826e018e172f60745682c5b85040578c0f0fe727f64010d9b1cf4ef59639e1d0ba47b3c87095c71858afce959f6e02861de57a71f6f15da2ed577cd15358c59b40266098c4b67e23e30e9d3949f270d45cd25b4731671dc288705d68835005056d369;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7b881add18fd0b2d00c72c8b51b731311240c74c6853ef2d401cae1b04b115d2866e55a33d71237c7a310c0c75df3291badf662b66c743e028a8b2a393f54dfd2bd275df94bb6ed0cb7cdee6362635e2927a72137026ef0eae8d932a30f46e84cb3ab5d2754b1c186645005b303cdd3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h437a61df252aef3b4dcebf450f304d6014a566a4078fca047cc43679f34df3c13080416d0a726f9b2c25e5ab892842dbf2df7d122ba4030c1859e4653d540872af91487bf0cd886e6e82d84420e9d71d39eb433fd6d8a2a4d25b19a4b8418259e68d91af0b0990771f8a31c3e412074df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56c56fe349b943bdaff1c463ab529eb16b860b6801e16d91c222a00b90cfb47fb8259096e3c3548f0b9570e57e6592f6fd0feda180108c7e78f5b3f7defe76828c697f1987bdeeb5cc17b60f4559c2c56df2a9f916b483f0c955864ceafe2c9e59522b0e3bc625d1e095ef6767cebc204;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbf5cdc0126d24c70172928cc03c9b940e99763539249c85f26baa837e9ebb69febcac7d2476e101466647a35ff1e5ceb09be9d99a2a252518231e370a0fc69a89558bde3da532e12f9fccd31ea7a6b2f185c073f8e3d81f5c60e46c4a7b1271c5c2f6e6b6aef54261b1761bd13cce4a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f7b7851d4029b9375389c452f6f31de5cc35a625bd3666882b3b9fb483537f131192e0aa79e6db93ece73632a9a7ff1229c8e8cba4b76402d436b75f40970b37caffeb7b99d44f96f90ce5587df85529912c72b3a0c18673c6f996fa3f240a5037572598e9dbe101c208002218d33e62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he77b7ff856bbe82dd86a3c70634a32c2c6c64eb7250faf2c0d9f8dfdf85a1706a97541d4433b8ae960556503ef83eae7e57d39395ab71e941d34ffba2277aab83f4c24a31e0da90f3d3645f0072c8d85769ef20809e95da07010f33d30e54a26f1d5766f5991651c2453238a42ff2fdbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2f3b4402dc073205c7892fec9d7c5c61fe38840694a0a54ccaf68e965eedc8f271b0c1d38c3501281102e2a2e5b6807e7f93c9344309c0435d087c3f43f6b035bd95ad649ed99f52992cb3015bb159ca7086f2caf007cd61d05d33af840c5539890d79c5a141fb644b2244b220a2a512;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73c275d8114f829c320bd2a0b071a6210b45edda3cbfb6bc220c4cf401fddb254311ef75bf3891b71c8b8810b8f1c7214c88450eedb5ff7981148dcb4e951ea75cfd67504219bbc71dd4852d9db46b294f4134c0bf7de53a1e0859a3c4dd28489dca4aa4b4c6a2e47a5d84f4d153ec6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcd0d5d8c39fca49b648683a45de4cc28d0e27a61a2d9fa3402e7ef20ca73a061a13ff6b35c12e790452e7d713e1650e34a6e27c6a02a41a367e9b67b72e5bf544cadef3c9ca62ea89fa0544653b852db4f973aa4049587184746c367026dcf1e5ec34ed84b28ca7026ce16b641f98233;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf89498d15fd1aecbe07109fc36283ae5c8a7c7d0dae6c2e41a4202afaf9310241ac8cb77672cbf36f6fbcb40d388396ecda136c5c3f710b57e81d0daceec919e4d5aa9bcca29ccc37a8a8dcf319b6833bb9751ae527186ff3c885bfa08e8cc4d6564cbbedb2c17af5620515a801f89eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac66e29535765376c71da9f921e5a55f1848e7706b86171f64d75925d6cbb86e53d1936c926e30d4fb6eec5d0e6a4587947b8d5aa0968d2e17b43560a5998d211921a52f0f4e4922b0e49211249221eb8975bef18849358954b9d48333560f54d6e703550147b4feeda096e185474f5e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h739cb8e54cf54abad9837e765f36363709bcb2ce3c5c99c9f4e281d85143407b64425b3c42163b215805b205c04640c9e5c913221a958848576486398cb75a8f664fa333b15da41400871613a9a0500e83c00ebbcd29921f2d4ad0dc4059bcfb8ac878c2cb4f7b609a0d38a4432493984;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h973f59171203241040375f5714f89f962ccf7b9d4e12e2dccd0edda341affa90e4a810f790c7f20b66c88ff11c1992a41ba0e4ecd36abab848fa3df48c78b392c5306beb6bbfa70aafabb1c7ab7affc1c384949921e1bcdb3d67b0df9af039116497376cbfab5c006da26a32956c18100;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffbed95ab2fecd94092027965eaed26e76ccd5ac9c7dc33f1ed660b743ef4fd436fc3ac750fa432796e5d09b2dcd8f9f9132656a604c2e598a8ef822731818f7971d7aa59efb82c89e73f74d496be0dd0c99704223a5705c7c736952719e33ed113f7a5e7945e232a0dbb330aca73f1fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe9da523d92ba97f5a67a27dfcd75947097f355c5e1520232a1bde6217ef9ac12a207fbb245de44ffe600ea5816d7c53e7250f35c72a98860fa2631878cdc3c4b7b9b62c3129362aaf69a82fe7f6d408eecdb7ab36d43e94ac033b1dcfdf3425c11edaf17cddf821b4d29765fe40138e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed1329d17a752f1d268c996ea1488dcb4004c43af48b142409a7cce7c8455f9790c733fe7c9839da54ae9c3f2489d150e02d33db9dc56b17b816bacc7972fc2168bae7464942cbd1cbb3f671a17108e84f4b48716296a621175c8d68bc816adfb9f42bebf3e57ae4e1d67ff4ef34ccce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d45a443f232a02ede31793b3e001ef868306c52c4eb697670373abb34f0b698ee4628284491dfef7d9b674eccac660d64d2c5f74afff09df6b8fe2e33d3f39858aa57e39a45a2dc8fc7014e346d2c740bbae5d7202b299389f099709b23ce75bd63af77b23a2274cfca18479b65658f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b0da26d580faa6c7c4c6142d63ff432b8717ecef97d24e5faea8b597e52a92000d3285ac96825691fb9ce2108a9b396cb12df36379c4b18838f411e17c0238706e427e49c013ff4484be01d8088ed87a3fb7cb9e702732197857212badb8949f4ebda33ed8436b91f6131f504aa78026;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8c35cdc501e13ba650f95790641d0becb6826062c2caa19a441dc212856a596e8504a57701c5cd88ca40c3b9c2624c84d1964e5651b5ef151051a2a0b88051522dd29325f0a17008262db906755dfbe0615a712d567d742527b352aec8901d003bdcffb24a9129722ec8111c0ac1d57a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8171ab067abc64a39336074f1224036f1e58ecf719582e29c28cdfd7aeabdbe5be3c6764741b0ed761222e469a21597744a616689f2f0ffe9aa27df92321236718edfaa6f2224dfb3f74db9ea9177fc48121818c4d2961d49e69314c6aeea9cacda66233e48d9ca0f07a262533dd6fd87;
        #1
        $finish();
    end
endmodule
