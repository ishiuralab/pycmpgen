module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [15:0] src17;
    reg [14:0] src18;
    reg [13:0] src19;
    reg [12:0] src20;
    reg [11:0] src21;
    reg [10:0] src22;
    reg [9:0] src23;
    reg [8:0] src24;
    reg [7:0] src25;
    reg [6:0] src26;
    reg [5:0] src27;
    reg [4:0] src28;
    reg [3:0] src29;
    reg [2:0] src30;
    reg [1:0] src31;
    reg [0:0] src32;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3])<<29) + ((src30[0] + src30[1] + src30[2])<<30) + ((src31[0] + src31[1])<<31) + ((src32[0])<<32);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c510c81fc298ebc0d22dae59eef5067630e013467ccb6fca351b2a42f0bd00010a78ebb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1273753b7ce008db89a0a15b0dbaca52825e74729c90ba86e1a50f94eb703288404a5623c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195785b46eaa81f394d194aa0e2effe8f1a24caadab3505616309b5ef0eee51d39639e7ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8199240110e2ebca0b4eb96990e07fb4476f9176b5abaa70b4e7fb805cab9c96225ce15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8ff909e69317480188f0e9a5b4aeb0bf0edcebe8dbf2bd59ab05d5e25d61f4f3439a800;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2126d14bdcc6d70fdb2e7b53bca7577ab0b51efcb3e3264346b36db375b4dd36897d4aa6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166207d44ab0d5cde5110f5d432ff5de74ab90d24e0783d5769a6ef4ca1573f74fe6f45ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18354bfb74143f58a18d4a9192b6b52e4b9a9f6a3bb16efa349819aacf43642f2ff602851;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdf38f1fa36d2adfc0015be2da26eeebba344eb2f994863e394bd767497a4516cefdcf3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbfe8ea23b1994845eb889e93ab9e3a70f5d0281e548b05f8f474484e4c2b0ba97e64e58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1625031c7e5e79e0a8c4c5ef0fa64878a7426fefba5938dfba24d98b54ac61c97667ba79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2000832c0c1c26131d1801c1d5f17826904f1e99a4e16a5d6b107534f30868eee0f5550;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5de315b410edc6d817e2653c5ff606e76f88d0dd2f0f5f2968a4e78bddb89d465ad98ee1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2055dc11ffb64995e32f7e6cebf760e5e515c5aeade4df43cd8fe00169c8dfca8eccb961;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a248ce373ee8fda0631fb03d08ac5b31f681fb9e723a212be460a451fe0187d0f0a6f6b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1beac23d37edf2ca50003a695cafe5d5c559d8ee4858d43ebdaaa9550962bff85f992d2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfac95353702ff64bf299a30f812d278fbc88a697f853e765ca9cd22e3c91aa44dd16fb58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2e54fe6a0f5ab9a4cdec9afcfc1686c59fd6e1b2e4d05fbee1b306853395f5377f3cc33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1393c851a1fec5d86c57c8268a36fd55616f86bf60d9557f9380e3afe3b0ee2b3022717c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10656e44c46f11c0c1b69477f894e29dfb3cb498d82c0bb10eee105e7b6e67abf7aa5b070;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f23de4242652dba93c4ff4dcdf40b45ead53dc5e1977e5183ddc253cb39f30694ee03d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a56b2056ee604aaf46a867865c6cb4fbdfbf015a8bdb5f0473308921040102cdd7359e2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb19f969fee06e9a8d95b47df925d70b46db421cb2084159ebb23f34dedcc746ede59a35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3d1f8e6a381853ba2531ed3d2f5be2671297931787269f9c5ed18db60d45cb67f522634;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159139abe0b85db815e044b5cb3c42ffd19dd5eae6dccd963cddd510443f25f608343354b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c037d2bf7aa2ee566843e7e24d67415e70ec820efbd6707614b0ba70933d9802d6ce0ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a892dd708acefac0814ffb5213f2db0b5c06468a68a558496ffbfa2cb3e015a142292239;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d72fc43da7b274a8df41d12b2a40fa401ea5e53e4b1c0332c042690e0ca8ec12dbafbe8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82d63ce96fc4687610d389ba019fca74395ea578fd378e802eb180253f7146ffc39f7d87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2dcef58bc6f8d10d259de1050ba4f8624db37a3d4c7bd56a720cef70c252b70ed157815;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b3cbb27495238ffc40e1ca4cdf80c1c7d2ce06be845645b3296043edd80b377e803a560;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b07c3db385c955abde6226785a71a9475f1c36e18a9460cc986618a5b516868fe1ec435;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185821c4c9c7e29d2525ab5a51cd2b752e84814777a4ef549fe1328e2cd8ca857ad64f99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h616bbbb4ad443e613e1c8b43259697e71bf1f1397d5ab4d6c7e36e251f1d0a7ec6e31a43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f838567a8aec00ab9b3c2c503a9f40a870e60242d25bb4e9efd10baac4d9d11ca9724ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114992b4ca00d184151083090fb39f45bbd202374c52afba8ce97f94086d17e718b46c38c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ff183a33242d15d95a3ce9346aca786747e17b8f03a740878df1f3c6b86c8f80173a067;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1301926139fe6f868f0255448b53bf7890ef793ea2772354af14d411521a05a0f613e0154;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83ae79b11ed9a0b522a510302d0e3192acce991eae8382e1aca7bb9da0ace47daf09a09f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38c96ef356f1cfc993659c59ba41692dd8d33a57f1769db8e943b8fb4cd330e7e0c6d1da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c8aad51ad06fdd0a51d84a17cf51f335dfc865d3a4d6420e05c759c095f532c56eec58e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158f5046c1c677ef86cee4da661760c923d3429105e672d7945f9de710b52cf2d8c01b022;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4f3072b43d51465575b62013b931164c25f3fbeefd858f3c2a990e8b5d14e6dd38ff966;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf753b7945ede51f215f6ac4035d79bbc7d0df8cea1640fbd4b08a4746d05b74179ed946;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67f60bd183f724a6c96198d156df816ac4e60262e76fea4715ccc8c530f7efba438b198b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23aa95873088e4918819ea0580a12b850d2e2196a3d97a39cb6fcffb1767185bf2d37eb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1314bed69176950359bb3856e1ed0f051c2bbba6e4e3616c056cc74b3ed4be4ff78159d45;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hddb2c21b6206e9f801f2cdc93dc302d4683b6671b5f036f457b84bd72c8f720dd6cb21de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156d45bc66973b694e76b782f520577a5eb9264101a8a2e27a00102c24579bc8228e020db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98cef82285834295ef084fe3946c8a5fb4f41ea71388587b44065e37af891e8d3d0fffd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1df048640da0538b20ffa86b0238fbef60e79ad51bd437578f5e9c7fa5e9e2adf1cce66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90dcc4c32cce147950d5d8212171173b90c4410e03aeae0e1ecafa525e9e7869d6471514;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18699c5c58d6bf0bc326fa4135dd5372db56aaa1f14db24b99bf3456c3d448010f57286d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147ae039ac7023d10dd0997d7680fabf75c8adfb254a2175a0d8c2315590af599471a7e7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17063891bc66d7496ca7331057abad1dc54489821686d4ef7803fdebb7882b31e8e67f5c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdec315ba36cc1fee35fe4f76bb263ff41a60053481d3f35e9d4df400475ed5ee0e9bf395;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc036db8295deb9def7bc43a3b0641f33d029a12312e7b0d3ee4b3c423ed00603a768a65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5f40910fce404a16664cab7148740386a2113ed95bc37492369562e18b227bb9d19a98d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f38809d2d5cb5573e5f9a4899f8cab4ae3b762e64d5e6dfebc1a4d0169588265b8de9692;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had2b227e6167942e750468f351917eabab654ee289a4eaf923d4731a9da260110c7d34e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d62113ce3de52a989ce23196b184648f495bdc01e1a4c5f39c207e56590206b54d67afa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104a9fee9b7e8c4379c0d88ccd971d0f503b7382c4c667bb554caf5ab1177998aae0352d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb201a37ec74f9414011320bde1efd1b74cf57b19ec9e2e6e644321d70a58fa2146939e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d3f507f3d12b1efff4be71118ef97fa65d641280314dd88f2d6b1db6e404a5be9ed890b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf85467389160c99dc8f732fe8c268bdd18e69c29a244c65ff92233828ebb25cd6ab2ce26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d1b9b5c026410c9d21429155f32096b784c04febd5727f74b0648cc5d60a9cc61e84dca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdaffe8d7887b15d5e7dbcfeae6c8822dbb58ec455c8d746dc21c290dee639c4f9b8245;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe15ec85e4e5b03966aa4e65c20c5f42b7b466281d7e6378cfba7ed73d35061305b672dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1d88477edc8cfdeda12fdfc09124324c88a0ed000d2c37bcf6d0b35616c781564798143;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h548d80f3bdc1c21f939764d072978cf2e2b08bed9986033ca2b19382c32e6aeaba2449a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b2905c5be6e7121ae1b06c5e0cf24782d9095c742f788a4e161766c7eac057990fe7d60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e53ffba12c4ea0f175eb9ada165535686ba18fc99df1ad063090b0ca7a67d0c4f2068e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143fdb6ff27271b26632f86232aba0c67a21065bff7234537fbf2b409fbe10fc7985ad31c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eda066e965b2caca188e7ec97e03a81108fe69580a88a8aae0262b3910b8e11bbd951698;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff80a7f842f7530cfe363393fa109446b791ad5cac0a9375087b2eecf495adaa5afb4c35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb90e809fd71935d893980269fb8e1187a77afa4a50e3ed681660b072287e4c7f1075486b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1248a9e971eb66a90573a88224a09f8122a8bc495320d02f60cc96532b0efdf34d0f6fa36;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80e340821af6e26bd37d0149ba0a99df7ecbcb405061991fd00241ea7fc3bf5f4a80f791;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1213de4bec26d3f31222611c98d4e6c41b0fd7551c2e7602d380f48dd87dc50ea83415f18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130dca396077703c92f0e6764d0dc7d4d2d7c820200364f7a14d22cbf5d532b151dd207c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16baf6ba44c5d9de05872dbcffdb800172b89d759db332a99c35b805fcf9367f9a86ba4ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f7af389458d60ce112620b33c0d8c2ea6e2a7fa8fb82082789e063e26ab02608af41b25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha12e38b36640e07e385a70bac752743179feeff9f466969d09592271c4e841f05972a3ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f6e036106ebab01829bf98c619b6cd8a468d117925469ee1da5de2b3d18340bfd17244;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1738ebbd79030cc58d24d7fa55113b43b8a0111e96a52bac9eca5eb821f6e7d9e47a35d91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1efb5ae6b165e7c224e167815af0eb95d86a444d3d84b9fc5d0d8550bdf599d725253ac5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce795d247a0f691f46f2be699a4223e1e7fc34125b001b4e04e33251b95804af693561fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1046dd97ebb62eace8b218934ac35329a222991a738ffd514e8ba3b7d1ed0a9d76486b79c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14108ec8a31b51b547600e0cdaf3ff09a73487806701fe27c78d00c22f7d572bbfff7247c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd04d13ec9e9fe614fd81c9bb98abcf40bb44f29b22dce09863a3ef36edb1e369c23d1e55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb03944101c68dc560fb480bc94c8b679380c98e7b5a978e35eefb5bd05f94b69b0d022f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b801bc398815fb76c29cb0062806905c046afbd7d731d468f2e5466a0e3a04639a275ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d64e1e4d243317eeba8d50baa398e18915976c990809fbdfdcbee1d9db0b47102f24a25f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184f0698a29439a9529ccfee48c9743ea3c434ba2f8761477369dce9175b04ccc1d0f4adb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d575fe4fa19b6d3d9378e0cf32691ae834cb8235990ffeb6eb445e740c0b874db206e2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7bdf764fa15baed58ec6399a2c0cadabbc7abbe5f1bfc47802e11b21250762afae25e0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44f3892ce043e24a73073b2559f2225f7274bd60fbd583c6b8f51d3bce9957d909344b3b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd16e8c402fed5b5f64b75cb34c770fac636d3a2f3101de5e46214a72fceaf9e5d589e58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a9ed83b984c78c8c23b7ad21be30523bcb8426a2d916c130cefe947976bb7b59c79d0f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0253300d4cf9c4faf7dd9cc2d8a1fd97d63ab8cd045ebe436348e27efefd2183b06c2bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17004982e5551c035b9f11853d82e3775f6a3179810dcb669f287deee1e929ce71aa57744;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf93f567426793a21a09d69734dc58ddaa1e505ed48ec6e50d8aefbaeb6bb79af45387fde;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h502e61e4d50868f66e047188044f31375ec539a290fe48226a8670b0bd079de70a5ccfe3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10957ae46335cd95a5fb71e4a7d9a1b9297ae4c2bc9c63aefddb621e98aa5f4ee791db0ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37a4510d96200fb93fc8cd4e953d794e9bb565d0e1abcbac8e1d2a1326f049089d933c54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a7b2cc0d598e29e972026d5e2d4ae7c37c7a1110061fa45267f1c90011d32bf0a5a4c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19bdf65872baccc8cf15ac7df0bc5088fcba3fdb55d5caf84bb3e4f1155e102000854db4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105d63dfa5a1e7c7a28c35b2d8eb6ce1ce36297de0236f8a7445336d9c3baeeeee2b93a61;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h335118e75f6f8758ef8b739a7ff54b5a6b5adc8a2e85c0dfc20be54b1868ad5d4d7fa0b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1baa1accdb0a1ea3e990033e13fcb2384dd42f9063bde7961916ea8ed194287beae95af65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab821d114779eade4fc613a4c0a7564b2f370b1a021f94cbb1e208fe0bbf86d2fc7f602d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b615dff9ad31b84fea20b93cbf59335326041d5254dd386a477100204493b92c117d96d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6fe5fc8f6177c8b635690daf8a6a949bc999f6a433575e3a7fcd81ea4f60134cef3aba2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1817002851254be7f1fe10cd9804e0261e0b8b31be625d059bfcbce1767bc44c5ed20518c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f496b1a2f5981318df80d271dbc352acdbd96253a5af1667dbf715b8d17eb102a29cf3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6fa88bde38b4283070350bcfbec35d5dc4072b2ad99fe4b470852c3a9018848585735ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1411fce2dbe6160e08bc68f1471a54ed938fa5a6a122da6c61aa50748a840c71253f358cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1911403035742a3d0082642474dd5c27234980cdb9a2d0a4ddb634a122980e98e002021ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bc12c639fa56a984f0452cebe6df851afab2da08a1dcce05842d059567f77c35a5c1029;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82d6f28d5087451d9ce4c7cbd022c000df4767db7b9705cb5b8ba486e73d692cccb8655;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155951785ca15440612a5e2955dd5965685d6ec3ca52d8a7b1cd0aa9f9700fe2d997ba0d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he97198362c96e5678970c079e8b5ec84795ba3b8b345e0c7236456db27f5140cd57a1943;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0e16e5389bb9a429b8608ee2b2fe7cfa33642375e0bd934e6b17866ffbaae902b462bbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195cb8a62de17419d1317a87bfca85734dc2a9078a084fe0b7dfcb8e7065fad99e0c70f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144b322ae130e9442d0b2290a7b5136c4b9485c0290ec59c5936d5837ba12c2277d98d6b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56432284504c5dccf11695c6af114256c84b967d76950f75c8034ff176175bbc1232d80a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81e7d00c3c978aeb7da13e96abf71c4c527577dc2ace6a84acbaf401b64b987ba25f2e97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f3259850eedacc482f3f2206d2469381e0edd62e0ef5712e4797f2008bde35d1dc612cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebba5702a1d8e71dfd1f0fe6b508a0d867af56aba21334db64e6d5f415b6ab3ffa2e2186;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42f4614fadd12d7442fb1607d44de1773083e133856b09064e6e2a700624f619b20cfa05;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1cfab08ed7e3edbac10200155817509df962c40db9ce09a9cdf5de8a1ef67b7c493b6a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf82d8694aab26cb1273b7f95e17cdd2f177a7c652b5d6907fddb826123dacb8bd7b972b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22ae1ba8edd4ee27723887da0240fe6c8938f8fc284f43dbf0b1003a60834e6e76758500;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e0934768ce3cf5a060c6266acdbe3bfc4883bd958fb75ef73450c5a7e604523a99da247;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2174988c2a9135ac8eeaf4fdb82f2e2f8ebe3910a40a84dd3f2c0ada06dad66ae244009f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12eb2d52a094c4c3b5b4a6e42435eb3733c659d6db9e60b72a00387d0f4fd70230b3aa90d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac4ba8d0b0608d1fe7bd54ef6b543a2e1eb4f43bdf230eecff8f2bdb14a789b704bd9c45;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177b8d303ef3b65382316d03543e66cbef6cfaeed9fcc92f7fb714a8e94791286bb653851;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a65feaa424d8ac5119db07bc5a17fbbecee79de594bb41a87b846f94aa71872b2ed8fd99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h513242989bc474f70c4d8b505bcdea2829959c6d323ef93a8a88df1f78314a79a23d7a9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c81bb37bc851230ab97435668195499f1b769a6e6fdd282365feab6fe486e56dc5ee4691;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd664d1e44ce501146b000491d2fc768e102c381c1812e3a4332e88613f40de0fcf15aac6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197df2d24f6d7076f5ae68483265408df7e0205e5b4670f1c846ac1e1af03217916821274;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1365b1308bb853e3e3ebf038c8a7da1e6896b831d70ff394e5e3696d6ee8e686ba45a39b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f9342ef36f84cb8f04ea81a78dff8cd98a21277c1ae62b02c8153ec7e46084828691b1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1280f00c4a973b549001f61a0fc8aa844cad0e91aecbcd5d302008c5997aff2a2d729b71c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habc2d915f3117c8ed727f2a06a52371ac7ebfe1f1678ecf8eb5b13ddd171837227b0db4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba56e1e86033f13b13df32b0ec8527aee314981e9c83bfc7ba2b6b58dd8d9c95caf67572;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133d11b0fdca039e79951a8d20b338f2e1c793811b4197b49327f785951aec43cf27097de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f8ce1581997fa858c0f7a0470dbbe16e2f3ad8e68cddcc9cd1d4d3632b37ca134e4f8bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166d73d349a997f864ceea9df110748506c8b24b03206b4ef51df53e34ea3a468ca7ef63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3352bf857c032d1d3122939900dc9a3b8d73a11dc10a7f6eac1b0c8b676dc388680be1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b41ff7d32636972457942376054fd0b156569c9a095cc4aaadf4033fcc524147ec56696;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c7d1c4553c0a01ece467d2462e5869d239283272075d0d02d15351f944d95b33b1f7f87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172ce10f4757d77cd98351d6c7289203b5e2394a22534b89e75097d177876e70ef4846b1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57fb8b0489cf61ac3d1a510d58e4c3921db362e8db855a3dbea0b53bf0c7a7f797ac4167;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f255ee31b3a98cce2b21391314cf1856c772eeb4d7bc1a9ac108c2a2e79589cff173894;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4a963285f0c0d901f79e4f395780b9bfcb8de24fbf40c69d512cac2de4ac4e5200dfc21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e84c689f2de6fe0b0d391adc3957d32e0a93ad85d5c135b00fc9fc8b39d29631f21f7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5e4104955137119af43101c01e054c06c66415004d250c1df2c31072aefb7338ffd0e35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h870ece5415da4031347783d7cfa911665d9361f8e9431584828fab72f0176c55d2d71f64;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b3e318325e4a3707aafb4679de51ff3a23917bb5afb2c1e19664eb7d9047d751e7a1b21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3fb9fc5435dbc809eb8857f3a7b93d9533f4adbcdfa33529fe712b0879123d5187cd8cdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f20a9072d3c310dbe7c033e0aa1b1a2706ff777c1e953b51fa4c68f413e369c3d6d2586;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc0da2a8b04393ec0463d9e7da0fc6a977eca2d8140ce1774742d5a86be2b63469534f4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcddb0ac41338a058817f89cec9ce7c6c35cac55c9bc9cb7f5d3e9b846c4c2d4688ede8d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4aa248140aec5fd8208b5a25fab11630e29ba3396b91c0a9ee8d7c80127597188d8dd8b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19bdb88a3cbc961d2455d8a2fc51c90eaac9bfbf4360f1092c98c0827b7e72abc2ce759d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6475241809726073e094c6b706c210992a684f8f1d2b2570c77fd8f4634d5b33bdb0e18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1170986a1e21c5e035115b8c06ef72d82be5d62b119440736c438547ce5640cc4cfdcf0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hceaf849fe614be7bd9e5db63d361b008c6091d6d71622d4110dae5bedc29762d2b6d1258;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16839d61f880822dcd955d105f66b18e779fc84dcbd76cefa145d0eed0f22343326a4f8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4fa20e4f2ef039dae636b39fdb9127be55f02c841378265467563eb5f1688ee0617179d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35986ea0a12316ef01f38a30072cc1d8cc42584a1f127f68b2ba7391ee5e6fe9846da25f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1e2ed44204517b28a934fe3cba23081c9eb5325dbc311f0e10f5b3004692d275e6b120b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc917cde0c26942f2eaf41339e205357783b95dc26de45042552b92414ff603b1c11b18f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86dc972e06bc1df33ddc1fbe6fd0c730df2691bc291c5cca58cab2a51c173e259de17a0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h225f7227b0f7f86717960965dac8b57182725d80937b9ce709219971a5e78b6966ca71eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13de136f0a5141cab37348ccb45d8f5effc00ee4c645724fcbc6a864eaa0eb36ae3482e88;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da8e7bcc191b52bc366ecf6744875f2c2a251e6e3d26142b89e55da16f044a75958827de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133b64fa33a2a340df35b83571ca24e7018cf15e79cae3e61394366eedd984c18879eb98d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff9786f2bb53875e75e46041d5719b36a1d574613292d32715e5a1f496735fa7fb9c2015;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1637d933881cc878b6d71874869db739ad581c7ba4c1057a8883c99c79ef8baa715e5f3f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dad3b5e89a81dffa8c8f14dc83a1c2447ed9ca5e28254e148aca554c695bd6fd12e51d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1ae8f7dce8545421dcf84857eeaadb6f1e89ba4e22637bf04ac38736c4175fa56862c8d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1c3c1c3d2f953d94f889dcd76413703debd2ef5010fde571e0633388b8088e5778a65dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff72b04a044ee4d4a7a9d200008823bde8e7339f19b4a5ca0be342fee5bcce97a2da3439;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b292e0989d80e3aa8be1547c49a99579644f7f98368d5b4009fdc78a7efd5094bc6935b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9588f2b929a8a32d8c45f9396972a0115a9476507535646b1ba9c895f039bd5dde05d8f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1925590da6eaadb74036376d388ed5c0cb703088a43d61bc1121e6e00d7a173a031535a95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152ce4b55f6d507b069780bb8f0e83b95dfbdb140b89e500e0d11c5de87a22ab2fe49f8dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41f0939ae2a04a7744a644b2f542101d75327bbaf3803c3486de904f27e24738caa721c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135a9e1a179254b94cb3cbde17d6b721b4b78d7cb2e83080df197e3984ff6aded0c62d09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd3959d723fb2d4d48ac9a07718eb885542a1645c93a7dd728f1b67923cd82187427c7e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b16250076e3d9c08f41e5744d000a9b4847da847a7d219d55f95f0da3eaebdf9b7e83bf8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7e0c5701ca013234bfd258c1949a45082b32ad75f2ffd3dc829eb13c46cb3d58d708ee8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5507a6d2519c65f8136e3f0052b6b4541a727015db77083c303b80a4497361c896a8c0da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h515364a77ffab9f18dca00bc22106005388307349e144335b1cd96f17c7831677864f4d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ab2210cd5b50e281fa5848fffae26866aa4fafdf31c610caf8514a957fd08f85e3f3fb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1499486f2f02bd415e8ac9103d2c53bfa37a03bf6f0e39343e185604ff272f80b5cf1ec7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f08d9541f7a4c23eaa53517666dde840962b7051d9951cfce56de4a687d329dbf85ec79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afe70b5a52cb156f6c0d9e476077daf2cd0f2e9373395866424147d86e06c932bb40e54d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0c4d721c12b4930d49fcb3148a5d794a4d3cebfc4e4c83e7387d02219572a7631a5781b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d7f969f2170a0604c60c54fc81eaacf2d2627c77b656834e947e8c0ce748adb6a47c500;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d69a26b152e0c5c5bd77df72cc5432c0fa6e2531ef5b777f4c1afbedee06e0cbcb2c1c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1a7e413d63a985d78add97dfe57d6d1771cd6dbe90590dd55b61f48cfb0d97bda170ddf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1177ce2b8fb713cfc9038d1a10d5f1bbcabd94cb64ee4922bbab6a158907f3b7e1b12ddca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1360fc6a4078a571a3889a142aa318aeceace2f4bb0b47a7a8a6dffba7e3d23da95788742;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h381b39450961e2072cad34d851cae4f6a0faf69ef0ca952d65d4d109780ad87f87ae8800;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h928be568447fb31416c05dab5e209d74b23c027b51a59e8a94c2a0bd3ae814e14cca392c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95331f5cc6cecefa43c3b1450aff281970a68228c84904cecad70399a73c6e91632a7cb7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137ac0963010b3e45e05b11be7cbdb8e6a2a8ec82a5db48dfd272ee4926ce31c129889a96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acea60bbc9d8f14aabe3ebc8b1d2e659a27666c0b070cfae06ae362bd2376181a0d18176;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194c41400888e21705117cd27f95b5acdce5f07df0c423be1877d52f56398a1fd087bd188;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1064615066d3854387d5235820d995e8e5b93ad159a1eee89fd481b07dad697363829ef37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4c950aec673a996c3606b40ea3e3313374e72ecc10670474e6434d001d67632f0617b43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132a67a5a3aba7a35ba97f7a37fd6140c1f5cfe8083ea5b0c9a7e3fa1c95f17b2733b8b24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1015a8194e5339293780174890e68cd0b794f070ff39a0634deab323ffe1aaa43b4893ac3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7161ee700b04213feeceabd45c6593cc96f3d32e70a259638649311aa4b7ed919c1d7268;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1244942209e07a805a91f19a0e9c06cb219570a1104de2e88ee1ac07acb9a470d35d0d4e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdcf539161622a1cae10dc3657e0129aeea2b3015d1dee162347ade0d1c0fedbd2f03e12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb625eb73a997e414c15517e32da3fe0882364680ce4223011f21e9853ac42cebf774e70e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15772c30b1dad6e72df2f928d8bd17a6b117ad1733019f889636faf82a0d5f429c8289061;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72b76f2d08c2d5ec748942a5d3ede19c822289653791633c7aa80c29d99017e4174ecf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fe74b84c197988b5edba5320ae60b340fdff312164d8a6098ea8cd7ed5a127f42122c0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c73f2c318e71d8aaf0b5a3f35e89c37f4da729c5821d44ed1ccf06916bc71194ffe5226b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e663058a080cb0567348176f4f7a77975df192b17367cc3ef9d639500260659cfcec788d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad28beacd3e553b58b15268492325e23f255acc874daf5dd2df9c8674e0399856bcfa97e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5a5222b98e0d1acf300122161baaf2d12d1a1e6cf15cec30ed957ac35ad2b545cb1f70e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97784ae9454f4c80196d0a1884fe45e6cfe389f1b5e21b79a91637f0d48a3003e383e8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d1efbee76bfdd9934192ae459319a97918733f93747aa8d3f3ef107340e85991c9545cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h425ec90d2b8d503570a381a1dc51106eb87bb4ea9c13b15dcac2f1f68bdf08ca0736eed1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0971360688fae623f1bcc74ce0dedddf5c9e33c712bccb1d3db2c6d29a4a02d0f243854;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1666069ebba70f1d6aae8ee42769135af6949a717754d9bd06b80795c015b0142c38b783;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h345894fad0d4f5f5a8b2c26ecdd7092382335e2780abd2ce4012bd427872065d1c98f223;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d93d107db77858ea9b696913673ce627660e2fb7827c37dcb9cc4cd930f2d31e3ee31d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2e54c086c163a8af5800b958fab4b83ef3820f1b85fa0473330dc461bcf0d576a821c7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h990ab662e436752bf26bfefbbee20797b5833fdbbc3d26014b6c1d541fbaf98b8a8650d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50a60ae63c2753246f8eb225c9aa435f16c865a026938e67685200233ddb98582fa1e6f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he44260afee9ea7b79723cd8a9e53583a0e2f1f5f8ce9337d21168babf75e7c84938c24e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17280f40f0aeb9457cbcf7338e8cc6d3b7d9734837cf81d781c474ccec20999571a0edb1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42e4f1588909f96cd1318298f0465225369c48e91d0d987246d1904f25d9983697c95b8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af9606dda8bb9d0154863b80014c5642140b82efb88c0f0e38738a9a685a856992c27ac9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a2bba3953ae0298e53690b5825503cffe85dd2e75f4c3d152a28f9988351061170b75fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e77968eb430ae2d55f79fc39caaa36ae602611267ba44a62e9317db22b280c45b8b38983;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f616203267993db5934e01431130b9c546442c2b62963f23f9e79252d558b004476a94b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c074adbcc3b61df1c7ad4c9ca59c7d8af3ac2529c7708b6296dab0014ef76d02c51146c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19940c89f0fb13bb7080aa2183525d7342efeeb5ad170d1c727916aa164580c3b34be4f7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57c900c431309b9079851ce343846dcafb0d680dfcfa419545eb05287f8ed9685dcfb939;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb93ce5e33d05829023ba6bb273ccef40e53d0ec6db13989d49a139aab20bbf210cb2fd58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14382eaa3660f012ee8deda051ce39ef6bcd6aad80914dd50e93bfd9849bf6875d1eeefa7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe50817b2706fdaa073298cd3e652877ca42101cbe15609ddcb1dba149522692fcac32a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c44dcaa3521847a6f6b93f92583e503a39630ff3f680ed29993e3a50bfadab2959b70441;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cc226eaef6280588ed878a265e66f0cd04adb5658ecd3df2d81d9a01b64a826975fb43a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11344d259cc1f3381adeb83904714708ae1b9352764d598fbbbd15a11999fda5e85f9bfca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb837fa5ad97f2e84c6180290f3ae177f7bd345c7a23f3e5ef28287b99f5f855172ffb551;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf7c2dc2abdb4513099a5526420b58b104796674264c254c0d5fc4eacf3a61eb37257bff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8465365089d826cd91fd951f50db592ddc2a70566874f00f8a92011305ce97d251d7c63e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a861a666df93e5aaa13e7e32ea9051a7ad0bf75b6bf3f729b7037633c0094a6eecd4678d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2469a9f375b0f92c6e3c2cd4a7245f10d0b8c819d6f6bbd1da112706e436a4a48c45d1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2a6d91e83d41e76a0ade62ce867a3a44afd7359748d9a3c1e07f9f24ce54f07f45aab5a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h649995f11f6a94d67363faf28380bff37381f3eec8d30307b1ce5075d9046353e8bc8533;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eca81967bc72b8bb9a4e246c783b8b14c419da883ac8eab8348394547c8150f978910b04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199faaa28057367e065a418a1dcf922af2f111b1f68359463596e2561fafb228830d32a12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125ae0b78e72e11b44ca2712c03d9984f24a0c44319b7831d57cdccf74e568a0fdf2e69ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1287f9346b9938a8709654ad72aa06169250d7b248722fa80e2a86666c0eaf209ab777525;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d591febf97afe4a8a5146ef00fd3e5a092a7d2c407aefa5ce7b36847defd9573c6e6cd0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24594f771a7a12eed9e060facd674c8c369fade49728e9a5d4c66e0ae9659a0b857c8c24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79cffdec47508df6115fc9062662af0162f4db66841b5ed24d5dd2511a6fa9cf06bb3e90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9159bc7240fd4332880a736a1426e25085cdf1c60a62c0dc051424cddf2d5f48dd9275a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafd7b009767d7a94eeb5d8845215ff0afc4007abe02dfc04ecfe51b0fcc91b7fe8a92288;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h265f3cb77cd4464449032eb02e4e1de7b599f4d399dd2e4535e657c66608859d38edf87a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da0f531955686ad1c410b63ab530554952e832090170b1d2be02f299dcdea26fbe8fcbf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he469d564cc04c40ce717ce3e0a4be3d853030884b1cf6f078d7005d526b54eb0d06da3c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bb5cc3a0d386cf67b0c471a37def1251a6fdbd8ed50b49c502c717b8485fad0d1776bc8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f96e0ee3734400f95972268051eddfc2eb9d6bb3a7e2530f15b7066e4c45cd651f803ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h940b712b0197e4d9747bfd3a25d32b731b6e1d310ddfeac043895a081360cc3894b422bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1955d73f8708ed8e91590a66264b7f33bad2ea3a1b60f60aaeef7f28a1beda9368d66a0f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f192af0004d8d02c641b170062bfc744a2a4778d263b2798921eb79f2f9224c2cad26f92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7dcaa066f31e91df12c82a2af3262820fb44a1505c8009fcc2c2b097b6af8b7863eb5252;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170355e9f152890a04fbf4e0d6971ca40cf62375693b80062ec98c27c4441237e9bc0bb79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc9cc224706e142bf18e276028b9689c7e60837259026bcc5b7861f9cc332b516bf32235;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd43aff826252128654caeb7d76d8f3627049c77d24cf60b3d6f802ecd6d21c6225092fba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10701ac619ac184a998987f17a97689ddc2aeeaebd11c7fe13093928861ad958c6a93e5ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h392609f12e5f73b76a24080ea4b062ff25f3100654d4b6c99fe78bbdcf835be4788c3811;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18188208094b167e5b30eacf82f29cc7b3615dd20cf4d443e70cadc3c4b9b0113df13d2ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13831e46444779b4893aa63441da0d7eaed4d100468f1295e33621ed4fad0a7667644f3c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba3c72414a72e3ea8ba011bfa8d09b44225d97096ceb2b24b66506db68b9721f9ccae414;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec382c7519043a301316562e8066c3160ce63878f0c3cb4dc3a4927f642dbb6c88aaee4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdac169e7053baed9f9b2642a30cd37d53d9a7bd30ac9b0f3b4ed4f6bfe473b812f8a294d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13835125a130f96cc8e81ab69a21f760de5d0d16ca101088e6561b33bf0cc1947b7aa3d2c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef7413ce4fe668ba4c511fa29eb5a36511e4dfe3856823a2fcde79e85b42fe5770752f3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha44764ea82a9c1b19cf9bee953acde9e08c5d1f691469cd8672604e181c7c23ae20427ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e761591692ca72f35de8b3bb514800ae2e864cde387ca8f45abeb06434ed79e45add7ffa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h574cb21faa577d504980a0ce513a44c952e72ddda85cb9953f015ac8f8966f9e0dd2c4da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a9bf8d2a973091e708af2726efa0c69e3f68b201b3dfe8a3443bb6f4e42ab8216522546;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ba336b202dd62be3a602d6c78ccf92e29546e21e3d9dc2eac8e08f18ca7db2afb89270;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d610d6e21f8b814e4ab78b04a212bbb9e830c0098f4678245adf36a2c4d9fad206c084;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8ffc0cb965655bd220d8be086e9867ca78ae8b3e620c6338810cb93bcbafa241254f23a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e1cb49b5fa0cd388efb5db8dce8853aac420b209597333de2652fae9b12bd14b707ea8f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h462fa785b6dae043660fcdfae1520f34214ab9da01ae3c673a02d5303462e74b974b20f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1163b2df3c12bea72148c20e6405366b6299822e2521779e1638b366c458a9c440684c503;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1baf7eed3deebf6cbf1547ed22fd0d57821d0ae40a0dcd6c3fc5b47f112a4e2320721e85;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5741b8f798dcef93cb928e80561b558dba61e6b482c5a828e2967f7500c584866d6fb35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc308ad29ece0427330abc4e7e478c2c92f52eef972c78670d6645fef84f8462123ea4677;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a104e37a6b50bdc21b463f434764bb6d92d29f9d055d229aa6622c725af394e27d4c482;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecc8f39e37b8ff0b34f118507af2bee08eb330c8791009366d86135d78cd50d7e43008af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52fc89ab812fc9d8be8fdd1adb7cd13c3d2d502a64bf0b1b3108f94ea101268941239c26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d28d3c61518f355f92d3c82a332bd87936b3c658e22c333d340086af22b4a1fa358b32e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17895cb050dbc801d957e62600f9c5cfbaaa5d84e05eaea53136a265bf2d5387cdd7133bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3a8c1a7701cc96f01ae78eba373c31befe9dd0225a0a3f542575c0eba949b04e2bf7925;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1249e7457bb936af8652c49adcdb3061069a1749ab1dc284486490b0856b18640f0f3637b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ca3d8d09fdf786ee98c088bf5ad9414fcc1b825e2d60a7720d4dfa609d4f7bb67492457;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc350726e3c6a35ee410667c13393c52d50839f550f0523284d45eaa671a7d9fd8fed824;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1627a568d6908ac2b2fa7c128fb8b5def02e4f0b9ac8f2b0e30e53bcae6368dcba6997a51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1caa61fe3eeb5af1677f6d0e235d7bcba38575627c16970d7d426222a1db36437de708a59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50278bb43dc723140681d7bd420339a53180a191585195cda1fbb80efdea60c22b72240d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e3ade226471987e58b9bf5b0a8917f3e9f9cf922f807319c1e2aea3a062598bb031c91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6ebb8b3bfd89d6504ac2962b61017c000a12ea0fff0bdb711c13b4e05884048cb3bb0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87e1c38369e6abf1a49e6510810f37cd196891711ae88cca95006eb8128f1b31f3cdeab1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfbab5a68f771894e664479d37544e933cd3e47a1025acde3624c2bde9b32c52b9887c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6816de9ee67489d3e4aa37eaf0c01d53a789ba660616bc926f9f81a3c92e65eacfc8323;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fa9202a9c54d914d222d91b99cdce9bb51ddd63af1551a787bd411be336b13acc549933;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcec770c55bd524ea5faf7c2d50a63c372fad21f1522922bb196447704317b8d46fccafad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d78f698d5b80f1624696ab03a4ad55cf4589ba6ba9fd49f0f9a015fe45a3fcdfcdad1435;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb4a965ff5bc93c776c33e979d37696858885ebdac5ead69b4316549d5fc9a4fc04282e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101c7c83eea4967a0ffb04f1aa5f9ff5c53dc60d711fddfc4b807d885a618653e74620693;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125e4316c6ac4836ec3abff18ec850f537aac566b354fbcd2c57eacb61f0d0714772dbbdc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha585811108772d11e1409161ebe6cf5182857b3a73a7785afec58ad449b64b1e27c1cd60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h844cb39e4b583be1f9182e867c161dc12113ed057efcd22ddd82c38c3e097af2d3a0c6fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101dc13f929a80f87ad18ce287cb67ebbc4b63bb1ab3805905e9bff1c6e87e262d85228e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1763d5bf641d61108fe3cca29d40f2f7d5d2372a914a9f886e9c0aa5855ebe888256b0740;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3c9e266f8e106b98927a902a3f9a5eb0051d6b72e35062762f013131e74fdd45f6e39ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14648efbae203b522fe998841748f6fceadba996e9da443a56d76f034b5f3c2efdcbd0f80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a9c9466d049dc433bdac0d50eb9c279ca93e567e09b2ff375bf6faa3ede6bb4bc664d9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d500a7908a3ecb849389971af99739b05b338c5b89d05dca879a5b93dedd361bea96ae2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178ba3810a62d8d904b62c3320f271b89f14f2adb9ecec87a54021f09bfc6074e6f3316f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f51b5f5c6b4b2dc020ed2cecd964ab6c291bf6751b4c88ac4244b91525b809adb6df38c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h514bab42632e5e6f7311a701f8453217219c1238e5f706732999ef80a0e8e8fb57b713c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43d0bbe23ac699adb127bf15e74d503ae5c5fb8aa02e6721bd1f48ba2d2045d38d8e892f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e21940c00ca397f561073d1b07e942501d6cc713bee20ef0ac932c60cac3ab17880717d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8b0bd2d41c0c82a791edea6397966d0e888f983f50c23a398ad3d4d22b3f53de2498d51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce88867540e1dfc296b8b25ae6fdf6106f25dc2e1ebee8f0b2665369ab082da3bea145f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11da21e90ffa546ed58a4416f691b0f4e98c326b5e59566088034a046984e5562d1655dd4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadec09ff2cca933809bbc2f1994fcaeef8f9557b7d95582fffbf39c79e88d58ca65a11b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h245e076bc933c8cbd20dcab2d82bc0ab986c879f88d8f1ea4be70c907a5f5b580b23c9ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e98e7df2917aec5579204c016d8f753c91cbef7fbe82a724c7814b20030003cb4734eea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9013415dc3bb6f008678eb34469654763d424ec533fe717f9f0cc605df8ab046a5dd1579;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e21dc2357ab8e81a0035467fabe39761b1298cb363234276672bb4ccb0931d319ce35f11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de4f9a04ba4f0ff98d2097b844cdb97d4d6fedc9364ecda164a0d33a0b249ec8f7ac2006;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23c17965724295895981e08df06f25b3f4d1b384281793b5cf17f22628b105516fc6384c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7efa5e46e8e1f45f4c219167bf9a5d95713b057ec2014508c18a59e1727a1568dad00ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a56d036682ea3849f0c4ae5e1cd26a011e82154f64fac7cf13e17c967fefa129af71ee0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7296b6bbfe4efe204c9d1b8aa7c6683ac866876fe4ed32eeaba82a417454db501f2a4b22;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78b370a825d5c700aa098e581858c665d7af016e9b3c1a68258f4dfbeb527ac6c4b2633;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc61cb15d6984e0b498c5dcc27981bf035a83c2b81eeba1b68d4f7b61c89070924c2ae88f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec7c2d2da3a0be0449caf3af314c2df19d70dd9ff4027308fd7ce353940a0d4acb9d2f96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1f431bc849fd74cfefedd3050ee54cb7a8db7f79569ba889993312a23e897c99fe0a46;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h474f1395b5f0ca8f0b724711af6b89c47b3afda9edcd8f8550fd27f106456826002eac3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1439a1910f371f414352bb95e0d83527bfdc780690ba083bdeaead8ac4797ffab44ffc3bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4d047afa572d46fc1a16fa031f2cc7954ee7de71b3646f1603b0c8c42d056d1f969bf9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14373be43d9c1cc678a1fe6dd4f877b661e49f8909b5c6410401d6810a62a864406407a0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hecadf41774aa350e33105eddd10963bccd8adddd9977c8f600344ee2b57f60369bb2ecb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a08aa4471cd6643c343b5e24e2a84483f2029f1c398139a2a1dec459c781f0018081bd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4f02c5a1a72018ea6c6e443c3fafe71828705440668a0996ad92d0cfc537d5aa7661126;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadfd1bf2d91a1ba252aad52ec80788537d8e8e3ae8408fa79d2491d52bccd43112cb637f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19537eee32a74c1580aa9b452cae1b917162cadff1f81f013e48efb14a5fb310ae5d8946;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdb8367a0d328e205aa7b5e318de25227ab09f0b8911f3190c6111cbc8944f8e6e52748a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164be5a55d26967f5a6853c7e1ce2971d8b0b29353e52c133139c4648a90822fd9729de03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd5494389fa218cc731d0c34deddb818af5f65bf14d904a95bc4024f88ae2824cbb00a79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d2e3ecbda8a97a9ab5a65ce352fe99a65c79752beb6bc9334a2cda3143de51dd41b85d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf26b939722f9f7d8a10c742576be65b1a5e1b77a555075e765dd3614ef6fcdb218cb7435;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0a48af0fc915ae7229246062b09c3f1bef6def1aa03ca6b1457661d7518f3218ca7ace0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5de8ef14813641751831bc47bcf93e196bfb9ccc9dcafe8af133b0e94d4f5a0154de5d4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2ca540475e946f4ce097d76edfb9b17f45e38b9fea1b977f8beb1cd62d66e3b1e1e2e72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ef0c7b76b501045a42c270ab78468765680ed74c670b4d241da3181258d3f1b82fd2c97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be4996c07500d3e9991fca5f45d2faabac33cfd568aa857490ba0ed13dd474de462ddcbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104b5c57cf4f34c973923aab4ccd744b699118ef650e8a43fe9f39e73eaeef699c72a99b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb524af468bbb67f14d74e862ba0190f3b481956317fda7b8d2568f893c13a8414966dd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16bda0457a0ba0ccbf8bdb37162da6676f61208f66255bf4f5cbf38badf11d84b786d7506;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc81a0b2492c8e16a3509b6b43362e224cf1b4853bdc7ec47090434be28091236f3445851;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70b677381efda923cb0be58f483480fc91cf00bb87f75af99a0188ae3d0a24f52d0dd4fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eebd40141f3139443c7ad8bcdb38e1e0e653fb4f1566698db15d860035c07d9e84f0ce19;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e09c732ce5e664c2df13a89572dfbb2f11f2a978223b4a9c92e490d4faf5cd5c05bf6e9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b658fa332c65e8fc9200a9b4fca0d39523d9c97595ba48550c997db3f6cd49395c670ea2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9dd9d9272ab7993021cc88f4c378b4a4a4dd6d3acd3c14bca4fe2edf00c46555b07aa604;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5c6e9b57b3571725578279e6a99ba229a67a04453a602c5892c555b3a7043168cdfa441;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b21c5e77af60d5f2c4c86f34da5eb8485643bfbe54565320637258df04207736419d55e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h521963ce69fdeeb0a65adb58f7864e3677128456413b7648f186b0928f7e786fe39897c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16deaacaeb6a9302c30eb9ab118a650ded959571f00c8012ef3767522f12f1d2435cbdf7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21843288c76a28c949f2961ad0a452619dc5f24cc43bed72e446b860f7195f3ece8b355f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb419238a1743f2e920686044408319b10c6ecff26499c8713f77823422dcfdfaf627396;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h297c688b74cdb7e3d5764ef4a4fda4eb414a618d617647c39d786d1bb26756a40bf0bf7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab741a8535eba410757f96b0cf535b023d6d8a3b309561cc3e10cf6256e8d0149d5829e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a438d95f27a44ed5afaa5a0ad0a681233a7d5ee6d5af7795a8e8cc547cce10936b45c22a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h682e356ad23d9b828a8693c563c2e8bdf12abf62b95d9fdf0939488f5b6a74b8622d7b65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16072f309b6f3d32711d6c61e449764f3ca5406548f492229f4ee31c48a38332052cbe7b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc15b6b0f3ffdd80f0f170de995ec9d4c7f97664e2a242f9794463af82b94fd910c3a33f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168a2c08b6c395bd644e99076814dbb35d9cc0080a80d1cc013232b27362d079bd40c002d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5a6d482b79a6f891a2456c4dde78b48806c716d1333163f8beaf0d275d0ff3f0c333ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12205f82f81d3b41148e50f1f3145dfc8a48b767b45929f1314ac81bd0e763bdf30edb680;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187229d83de778afe1231387455b9fce81226d1772cb9f0623385d2649c4db2e024344c6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123cde17bf1c3de13d87f893a70f54ce062814543b7309e81e5d83807e1f695ebe850d426;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bc6694a8f21195f1425e51a340a06aef9d2df8a4fc8e07b1d958c150c33e3ab0f5a146d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7b436a8667df562ce89f83c143e45cb2cb1897a6cacc92dcff1fa019cb8067aa8a3ab86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe008edab14931beefbe2a26e6aee949117a574e77fb8fc1a803d95f8b81bd0aa69aa806;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67d5fb888229c52d87c3c58a81d6445d1077c92a482080d7ad0574ac934dfca04e2453da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfea56d5de847150719e59b2d03576dcbefbe85a549d1a7f5666b1b6861fcb25ec90b31a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e0641e1889dd152991de64e170d9db788e419d2a3ffcd23549d423d53c6d4d2721489a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc6ab6d7e279ba9368cd474f8bade9922018a305325f8b7d92bef021be174ac5ef52fa48e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1b890ef4e146bce63138f02ec2a2bf2ec2f9b59ddf01772fa87dd66bed68b0e0acd9327;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fee352d534614de25c274d045a4531387d97e3df4ea0c9f2e0f35ab1fe49b8e89727cd4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d7bb70600736806214c7e97f602d3ae3b3a62acf178b671a1f2a0aa42d20ce8b56450b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f400d3c77642eb4c1cdfb3bf01256f4e2eda43446f29a39b760c24b7f4f510ebc3231d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b0f35a03543a557204074720ea7ceb74873590898ee78fa671a68f492d6261d3aba426a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bffe78ddb14b45f7dcd4f70a58b37f85d455c38ee6896f11c536c32385518ba8d91b7c5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc83149980dfab3642b8f37d621e009f1740902f04f7ca9f08a016bcf09462da49cbb3cf4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e5bce44a9340c279d4436ef990f53f947fa59107cfccaf7e116ebde5fa85ec8f7c4634e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3e78e6092586a6bcdfd0a932c5847c276faa99946b870507902e94c99a4f512890f9396;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bce64c5a2fc1eece644456d9639debbace375c94e25757ae7ada7c50d2666985a5fcd14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5b529c4295658b842022a014ed74930de9a100ada5f8127cc94845003fdd8826c70235a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13688127ac7154f191fd9abbc438679c357c5145d22d6e5a594f24c4b23be895328d8894f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abf62b1c080e531d2e820d3ad1c3b4edcde54ea2843f264ece81a8168e3a09de98b8b611;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfca4aae2f9cc648a3f777bbe89de02838113409375fe932029e684ef8d51dd81a4d7056e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3390debc7d8bbdf72ec07c411566d7cc224df284002027bea932789ea181a615cfc0b6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174ec49b1e4a60cb0a8d98a3556afed9cfd5dd8a3f3514afc1a3c98b530cbe1c50459a3ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefc2c6345558f329e258ec2496beee021e36d73b00c0bdc3adf1986dd2dd22b827112d61;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h213fc350b315738b1d8eb1bead57b59a1007c978abb4c1dfb760e0ed4df802c0e2b7bf77;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19af52e1cb1f9bab0fbd9bf179b2335c87f7e9bd618ff09efd81626b4d5786f1e60c3a31f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123f84bdd959f33c2efd5a8a26dcf99685b2f3a6ba0d501b4d00eff0ef715e2e02cc555c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bf1712cdde2eb1ca95b67cb535cddd3d93fb2be80c6fb45b6a1db65a614456aaf14dc28;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d76c4b9d73ddd1f4b61626ac5da47aa6996082f6a5d4e27eddedd04bba6c3ac98dd18c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fac51289db12e781f8b77c29890581e9e42b4c132aaf449193fa06fbe9890677e6628de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b05fdf6c1b5cd76b000583ceb90aa248e065ff74aab6fe3d9260c35fec9e832d8ab061ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28795482bc267f9a5fad6e317afdba3fcb2ea2b5a636690a1afb56d29f90ab263fc0bef8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1263513e101670ff345bcd34f9e3c5db947cb9d3d623a82c2fc8884d46121c0810f58672f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6718c2eb061ee979960b63f9d9dbf57b54b49066bb40b46bd745cd90a1b7aca68860a29a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6167e740e2223824ee4c4da5d2d0d4ff2547682bc4df0ea99e0d311a6d12f032ca8f1762;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab3367b0ba82c50f0128327b05017e9003cb90489b0cd02d682b7d3e344005fb3c429ea7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172a1070a162bc5ce3bb5f887e9bdb35e2ad572db554ec2df9be79d262de8c0840b7bd189;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11aa8db6611d7c1c12b6b29c4d736087e03645f81545afdfe006d8bf69d455dd953997ca4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb72aa01018ef357f6cce9732fb6adddaf8afa35acdae0df6c5315a52b88f51f6e25ae802;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8520f1b0a74be8010c5ed418c69bfef240e33c9ea3826749cc845e6ff227c44d9772d093;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb6d98278d748f3c12278ae3bc584ac8c42d1fba0fcdbb97fa3d580be401dce8d72740be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1daf1c7f2fce41501d9ee457ef4e40b3a1af11211917df28b0e34bd6896ed335aa7b201ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62379d378ff55d7214c88322cbfbdba358150bf083b8323f72be0f57fe304fd37f673130;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f29cc276af77814d848322edd2cdb52cc865589ae9f840cc1ba22756782a774bad950b14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f8cf96e8bc642f968a36a5d6d6c752e0ab42453174ad090201446a569fa990e9a910916;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156ec7f0866e2e9e23f1c4f5117abfc43a36db44ea01fcb55e4cd8f3c07c816c068dbb92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h272ceba3fec6229017ec6b3d6292d36ca6934e0c786f742885394f7827f7dedfa5c9eb7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebcbd779b8f3b6640dad6238dcba1b496d2bd5bd9fd966cbd7bb928d3fc508cd327b69e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e86de0707150786ddd51643bbe7fb757e627888af4aecf516b53802e7e2995c36c853fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1946d87702c8c0a912f303b731e441cde342fdcdf8d9cd44cb411866b18669a21b0e07740;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16445ac801c90802155eafabf37810da3f3409048aa57e45385489a551678aba86456ef08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf24dabf139496afb21003e1eb900b04479c84b9e71333d4c57d5722550d252495ebd130c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ff55397b11441449aa77fa056dd8c9584be437b900c2e2af7988616ea6644db98d2650;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12594d3ac1d44b00ca14f9cf2ef723d7b7178645e21913698c5952bdba55f7c0ae9600852;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16896f87590f887b07e42ec3f8c9065cf57639bba54cd8325c1e900b7349d7537d4a59a7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae90bdfd02b7f761114529c7f64a7b5eeb53fac626cc0d121fe4097bf22c3a06e3d07c1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cff455fb4b0ec1f51baefe2a597da73288007688808d220541abbd66e314d23c959aa2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a9b1274032101c87d36e977fd3b2e19d884206a6d125cff3fe7c9009f71064592ff9ccf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e41412f54563dc06540a2a244b43450a70b2f74690e396b110f3c149b5a2b4ee135c7f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1fe997fd2a5e33ce21aff6491c350cc1574b3471e9494bef0acf199a41cbb7d352edf65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h809688f7f4193f256910e28fa388c394064c76918be25ed91b043659ff293007596059d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e2ade13003d6ff75fc31fca098c7c7b2325586bb2d90f7d1bf3219e717169bbf829b3900;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ddb3438701a3ebb0da2e64368df03581c2bb0d5e751441437686079602b63bb4800a215;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he926a81f4eeb5167f2d4426cd93b317f95ff66f15bcd675b4a47ebf3a1b8f246c321f143;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145cd370bb53163aa976e7530d355124b0c8eb9678eefe3ed528999b3631dd9e162042fc2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18aa3761a3a965a52b0247d13257267dd88497ffe5d0892e49099b52ac1800a685203d02b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c075f81403b4c9efe1cc65d7d71759a8b0b4ba2f4ea4f9ffd5e82570850bf1d30c9027fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcebafa6678d7872e3805e0b337884e47c1623ea83b52b09cf37376072fcf2a46928c6e2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d73192d1041a66b375519cf679f436b28866c859dd88adcd935bd89c09b4164af5d981e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd60a913db65951d845a843e7b81e5999ceb56113a229de6a6b7e8e5f3e5f3e4cd1b9f4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14aa882f8fc7b26a75d7946f8f7ba24bbbb5e2469c3a2dfde3d9b4d2beaf4fe79a20c65dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfcd301cb6269dc843cba77d3495cf772f448e9652c7b649ab9911efe19957abc6f05b02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ceb3389f019c77d7ac5fdda6f1461bccbe65428e5e6ae7b220fa704c05733de307a8d429;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199a92c51f0def3e4d5850252e3d2f6cda92d920f3b3a5a568dad985e64218c37ecd227b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe65a4da190d60951ae5bed0ef23c7f2ac8c32aeb290ee818d726cb64b152a79201fa6e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190c3acad35cc39520cfb1c1538c33f8679ba81f6e61b8f8cb55828ba9d5e741c8f3041f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haaba509f20df2afec5b04f3afcfcf89d2f2cd7707ff4d20465e3024b2fb8be3b5d9d7244;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10854845c20ab71385e00ed04e186ed3c217c153f101d68ec1a4d9e9e66fcdb048a233240;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf962b3e61a0ab3eadf46b657e5bde63625647fddf181595244933c1f32d68f1a4f05253;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dd361003e0b6a95d504c3475e06085875266304fc8f6f70fb2e394f767a4b7b23b4ac3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd37815a1e8ffa61b7617202a7a31d6304d17df53d5b005a84d3feaecb37234212f1e657;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139c31e5ea2ab7f16abc59c440b6b9048cd4583503eb84987ee4174695c963774ecfa50eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h828bfa2df0934211754437d4ac135f07a1a6fc6d15b208a8e6e49d7eb9cc4dbf3b6d84f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6ebbd8059a088e1c3ee2a18ba2ce014e481bd45cc4b97710e355c05d4da2fe9ba354f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e49e6d798974aa7e05474e843c568929de6267500174061000ef6f1195945159d5544271;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4835181abbac5a78e0679a0a94d46181db6fe8cce5d9db056cc6b042c111c741e58f35de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156fe513caa7ebf887be41435318afccc4aae3a4304e0539d03eeb82823a87f4cffc58fc5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8e886afef5bd4730a5af44cd97bb44df8a725add7a3dd8468c5bba7d168a83f4cb332af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h548a8398eeadda69fdd31b463fd475ed7497098da07ccd965bdb793906ae8dc77fc05382;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha372d26421fd7913a2fc8c745448d9c73c8b2f026645b2fd135f207bc9399b0e544cd25e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6bcc688778bfd67129fc415992386413491e1c9fde2286af1dc2cba0448d97fa7fbe3ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e72520b9923b96a14974649693a303e225e450f07ecd13035ed47a036b99df961ecea1bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10511b3b1ef8e656e22751e8a90ea82a6c33ed4e698e0aa6f15abfac6e53e69def605ca12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4679068f381cdb3035dda4e6ab2eb109b26b75033ef08e91edd70a73859e84d8cfa11e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36322fb6f7f403dc96c55229a6031805d5cff4d6b6e7228279ddffe00435533e493f22fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc80adbff9e471a22cf124972dc9b1897668632374e4896770786776d3bd70c3327e77d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a9c007b5a0dd926c1ed8a52c9f2eaec8cf91612a8be3bc6922fffb4e6b3fcd723df4025;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19942984d0c37228d87c71f5f4a91afd39c1436a591108d895ae169a5c0326c29047fb6a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ab024dc6699204ecd808bc172e1813dec26eedad87b26059351a629ed8dcac90ae1129c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he24fd35ff73678fe7f1379ddbc09973cabe862e130935694fd5aef61f62d8fd2d312ef81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1396c1cdbb74821ed638dda64ef2790faebfe132e1392e1f983fb31d19efe6df78ecc7228;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1678e1bd577c1874b9fb6346e5d1435352bc126dae15d4c73016f86015bd4b6a246e88ee1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb03ee34743dda84d4e1a019f47022b7e7a8f721346c510be78dc89407a79cb386582ceb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1205962dd517bd1e08bca454ceb4648c1ecdee13dc3c102cab5e3d8dcaf5ac2b63ee808e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6a905d975c28141698b250f02ed91c5e83c7388a7639e6c7c48ab355a86091df6c3086a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45a6a39d65ee02cf7f3c5d6669b162cae4f383d06b5e3c40d6067773f1b4e9a3883efcaf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15246cc0ac649a745e15b08af50abf504d6ac2d78b46fd36bcace41057487766b43d23863;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acac8915db974f94e345c504696aeff46bda4887857594e26d45b66fff74c12429f25a10;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h551a4e761bd97a2f59fd57495952d44e5cf91a89ced0b23de2d4b67b68596ddcb8f09c74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb65dbb3b68b242206f7cad782d05531cab369b167f3da74c514db816a837c818fb96807b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af77b1b1f6e6525eeee7a8de62372d3fe13b867ee29c23b01d9193cbd628e43736006bd5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he026dcfabffffd60311b238bd5849a935014cef0c708b94a1106b1412b1213566d857469;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4073edcd1478b559e4aecd4fd61ca11d8c5e5a19ff9bbf5ad9493124d03234a4131153ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103f600c66678eb5396e92eb71c4d0e95a6bed0cd444b66078f6257ddd4e944ef9755ed3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1947a002f0b8f445f2f2ad211b8ab243c7275ecf28179ed5a87ebd25a4278725f5ccd6b2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117a7c24d61dbd5ed5a36aa05f8885ebd41bd1925e058f78523d0862cc0186279f0dbdcdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1305d18329c9e25c6af54e4977feb967889f8cc89b8019a992c6017da8bb079457053e6eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170747bc517c0a508ddeda80cac1b441229f82d2454d5a910c4a7dc0b110617a62a2cdc2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ed286b6af78b87010766ed44f2acc0699eabb9c046521baeeacac4c8ddbac3c17f7a74d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a3a1195b3953077a32cf5e00710c73475b815e4b58b3791d9c197b7616ebd0469f7a222;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c3d98029f02b25cfc63bbaa1183668df35548c12aa49219404f7a9197119985680467d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e92fd83a33f58b249b4436bc254a30987eddcef8f4587739d20c6a0ddab83adc8115615;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1190e268f55070e5bfdb0a0b310e0a570848a975881db74f0a694a776f22e9e7a7e53dd40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20c48bacef9f55868379710314121595a19f90772899619e94f8504191124c25ed81e6c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3d23a0b0190509e4fd25b77416d56dca951cbfaa0a1ceaa3413b132751f460b7fff44d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aaf1267d9d83f9faf6bd0fdd3024bfeefaa4541d3d74698f1eb3cddc1176f1c3bd02c7da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4b5a8da3d1b5451490e07a4bdea12169eb605a749ea32a74c5cfec3325bfbe349525e3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1896bbc8f0cc1a1a3f7474e9e594aa78b4f2d281defa2bba2bfc14ea2edcdc80dbaddef21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a8622ffea1d84076165fc638a283667b0d9fb0bb7308534377c808d3d6f5879d3dbf10b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdf1d917b79f7824d439fcc53b1a587d94b25ba8ae26322ec7a0e9d9565cee3a860140a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184cdf500fef65800845dc1f5b907c56c73699ae9c58c856408d007e777f2292b1435be1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9fe88e3e2ce64cefab1c1dbc607affb3d13dfc4178dd50ad55b1dec6a441c65e8f9dc0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e9e59ec85b33ac0583f43ea76f512e823da6fa6bb3dbddc1680b9997480a7c178758b06;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c6c53a51e684062de872836bcfd39da369496e35f61bcf3876ea7b92353bc17f5ea9fb2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b21390792bc97a0d00cb7f06fc4a98cc64e8cfb02989d10d76994cc378ad44d63abe4083;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9438bd2826ba720850058ec7d0ad26e63bbf7b14ddb834d2af5fec87f5949a7a2482c217;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haaf09bb8c3069d749a8f4d0212754371d914eaf7e003b355054c9c943f6c70ca57bed93e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h818f311365b7089bebf1af3bfe8dc5d84f72d376c8321b46377fece5c1363b1401b04c65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1547e73b236a0fd01494c26cad1077d6f293f212b02c86e799208db7e0079956a0e8a31af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bd837dfd08fc5251b4aac2155e9dff479cf8c8c5949749613791fce84f4abd807753404;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bb43eb9340f0720a1c491630f52271a1f4fe27c7b51ce0abf26b1662cea8098ec75531d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122308c9f192676426c5096e08f576a1072db821025fe5cd9645e6f65c03b8a3896c441f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f910dd4ff2d9a42ebec81a8ad8988b248918453a617bb1f0368041a9838e9a53993074d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4a88b1e2bdfa5e19a2610dd136b156758c44648a3e7d0d9096f3b27f2fd553bda8b638f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28b23cfc12c0d49da3930a5695ce722670bcdc0d6e3d84042bdddc9bb62da49a29b2730e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b024c110924dea34dc0d7dc45c2f9d1e5ebdfb2c166262060f612cd4522e28471ecaff80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88b00e2f4d2b567761f945a4145696633d9bc129fec3abf8dcc1fba80820d42a0304dc5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7639b727194d2c5c80f2ba7caf9f2845875e343af24a36c34a8e04d758bb42248d51851a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a7fd7bf3f10e7d0b37031fe53eda2f21bb0165d75c0380ba3fe27e757fbe96ac75bc856;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc184515b7ca1e129bbf44a57f8266419c35386b71e1096a01d61549404722159a838108;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5259158645f197b509f847c0464017fc5313cc6fed2a0900e096a55842a00897ba8cc79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145773926fb415a3342d9457938998ed686c69d82fa7c4b4e54cbe435ac30495493c5aa2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb109cf9deb8bdb5cba457c1d3f6774fd6ef58675437034b2d1b2b0fdef004b672924897b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd20afb65a49379f09de0d7868c29c9f75ff39a4d5e7866856401ceae8379605ee311f44a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48c25733662e67285079c896eb285b2e2e9e7d964781c1b6268c24c25e3abda70dad896e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba20373337b5ddb3588240943ff5ccaff55076f72d6f3bc67212a0722b430b1a95fd4949;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c78ed20915a94c5461fb262b55f2b03959acc9bf86682ba85909915a4075e3b75b7a5bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197270377dab5fc0e58b8c214c8778d8db8af5465dfbbfd035e87a0d0944b2757625470c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17830f600f7f82847661ca2010080cca0296ad1ea4695fd8a9161e81479d7136b7908e5dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd26efe740d61422b90b1ed009f2e4242481072b953a9f06637462c09dc06295891c76d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f13cc8c8b1d1a1d628a561b8f30fe0bafe418041b42ee287f41ced3618d34ff8210bcdf9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1506e91c149f567a38dc212a74d82e491a02c3aef485939f5eaac5fceb55f42d5716d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25bcfc286cbb6a2a7c45829ad510ed73c914cf7727839c1c6f1a42f9d8aa77130e242d40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6376709c21e63fad92c18d20e86d5848f28a69f6e0bcbfd98efeb646b002708adccccea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1178c5b2f7df66f6536758d91eeffe311ea84b563268abba172a7683b19390be055d010d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7a310239a9bf7e4682dd45a61bfbeecd2bf4fa4fbb40a46cd9eb30f1c4bb4c4c81ea300;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34f05bf48e18eb717bbc564369abace00b3883d74dd30aa24174609252b68f09d6c09b51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc37ecfe35bb87caf28d251cdfe11c9c9fbbd5df44dbc6c6145efb9809becad44f9766ac5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ac4f55997cc9cb4199cbe37bdc216ed119a4044416e63008fe8114a2aa2b917f5b799ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73e098e0b965321f515af9c0f7ecbca338fd6a6ab6c690736b6e2e14f8ac2950a50e0bbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f586b3d3e0d794c5f9cce6cdfb11d610c1c104f913f82f1685e98641073b504bb4239fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117fbea4ed53d812a854ad8713d01733cf722ba8efc3fb8da0bb9151207a6578ddbd9af43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a81bd77385fd433e4499706871c0495ce4bde9da782b711d47c4974624ef47890b475aa1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fc85f4141ee9491fc40421de6ebe9d37af977311ab87956df29a1ee5b964cf96b99839c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bbe1f9677b60c317e2997959307abfb7bd44d037d7f2759530a0e74973b37ca77921a7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161f9ad1e70fee07925d7aae4a623292c0cc7f0245977e864d06f21978d844a7f3f7fd91b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b8da58586934d235b297e19248a1a26856668fe5ff2e261f4f5ad3245c7884b01fd3e27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93a1c0c0d9c2ac8d745e516581499e7144f1ee5dcb2071cc7aab876e7c48e7380d1f0803;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b825c030717b4a56170b842c8b19a380f7e8e5d65d951b110ccfca7a4c78b92ea17951d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1bc7e2cd87d2c288519c2ee30071226071576108f65bb0e5b4006040182239bbb4ef9cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdca08f797096b0c1094beffea568f94aa8a93253e6838229a465e0925f3b5427da2900b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc9f2fe6278c1db4e316e72ef232d51b22d7598ce26d22caf8c7e5fc7c9664f995b1ef54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12442938e0d3b7cbe7cabfbf897b4796486f00772a4149d074579f65e60cbd9fae86afd54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181ed0266105c19301fc80f665c31e0c1de45799f4a29f4b5efc4d45b6118e87214a9ccb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f9b194a7977ec3e889d656ac67555a111cb045c5448041c236645696208a505867c4abb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77df58947fdefdee018487723ce27cb15411798cfec453eca75c9921819598e99d0c5766;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e8e6ba95a41d158543d58a8640fcc1b58291d517115a2b54c919aefaf66ce7f8bf34baf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3fddb44b6ee6a0def9cd2f348eeb5df80e4ac528d78dab99bbe7fe793733c7c5cd66721;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b902902a56b3ca79f4cfbb611b0e42830db7ace58de253e417653e00689738144e65dedc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3700ad374de5088921baacba15832c4f138c30e5f3a45e127524a1971a4d59bd2b6fda0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8ec06ea110424c07836dc3c79a5b44bc01777acc3c688b6b8bbfe84b722cf72e2021060;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1983e347c9e3b81141a50d03252cf1a84b5930b136f398ea92476ceac9cbdc16acaf04d82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87c335fa7da7d5e595f2ac4e811dc0472c7f974537d75e627d2109b8c8fd34ab63a528c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c14dae019c16e43d612622226fe1ea3f933bdee69be2baa2a2ae19d0c4eb99366abbe5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heaad43f07dcaf00712220909a20bd52e7f4fe29eeb144c6b7e79e80b3ce7c935649e8671;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141ce85b81469f5507d44a68ea37a094de6b2c13f278213cf3f612a8c06555dfd7f255794;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f33ff6619b9f89c31414fe35239967b8846bf62ea9414e408d064cebc39b02c1cd16fe3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e63adc3588e26a0dc74fc1f77c7e7b3e0b7ee9ca4f7214019dabe38426f0bd925fda050;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had0ba1870abf51af00e35cdbdfd737c2b63c5306e90a42bc9735522fc569e0d1220f446d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5cb48dff9b31cfb757963d5f06cb17a06aa5028c49b0b1bdbd4a0c97077de5ff8f00af7b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9419c54f7724203f014a436b7b9be56c2f22d4da09f4c655cfa894e821de09c7da852ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfabca9ca9f8298dbf968bacf9404dcc6742cff7e209b198e9fe0fd3fb0f7f1f110b1489f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67088709761c4a3c72d8421976c37d347c2e62ea4e626cfd709aaf6c70dda04b08e88a8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e799f53d3f0b3d502a44a4881340be0ebada54df86828180447f1fcbc3c797b2f15dc10f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1019947bd49a37be2445caa8233e56373d531da137260a8e89a09c2208d60e88fe502be9e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54af27868da34dd65d815109ad8ebcc5d19668c5aa7adc972e3c6f30b19111842c12a909;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123589017e8427858210ac160ac737cc556a218a55a79ea350b600eca805a881678288bfa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4feda295123c04e33933e265fce7a514238865986d7a78db38f104a6841137f3a9458cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heecbfac41a563a39c663f534ab2a053366d810d3afbb450ccf47c6edd78fcf548fe00001;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99390e75264ca6e7ba268fdcc89aba4c4a1a83aace58ed51efad03e209b95c42468d6774;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7958790f4a33276952d48c788591a4a4d5e3275fba31653d5c368cef139ac60b1760f687;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15feeccfddba1f3d193c1dfc1eadaed89c985e5167361a785f3e286a1d8f4b7751c7360c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1095c9fd4e3440dc328d907368d12708afe02bba423fb6920ccb3ad600f2fb082489c18d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a4c6fb6fb79c1c67f5111d2a713b23f5a8fe960b9b8f1330faf3be8f5941b8e0765371e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14dde58d56aa9c17d9448902f33822df28246d9ff250f55b80c3888ef36d67aca14645bcb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd948750e40bbda7bda0f8434d1c6c4a0510b9aa0175d035cc38bdd6c0efe3f7582da21c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf67ffcb3a39305dc6002408f03afeeea06d50d3be0021148843f2860626416aeb966027d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e788cb1fb022374ddae4acbb43dddeb5fdb49c142f6d2ac9220b48c6414382a32a1590;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103bcc8a3a43ed84e19aadad82fba065d43abcbd82cdf138278f0165d8f0506ecdcd1f4f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13604eeeaab258fb9b1d29dfb20c4293073bec2682493887d1270b30c7582e9a21c13096f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1984709d51c3991bdb0be37d8ddcd114662493624ca74bf70c5afcf189cdbae55f957e457;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc4ce48f94feb20b91e62677e8be5ba05b1bfd42f33b00d906f8c2ab45c2de6330f3ea537;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a4ea62670696c46bec0f90c24d5faa8fbb98e6afa4ecaf0e4fef484561008c14d17162b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f36f740cb617b6dda2355cbbf2494772e001271ed58517d791405caaf1ab87116d70cce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137c40ab3d647ca38e14bd253d66f3120ac1f9b1bd30bb2c51021ddb8b0bfb2994237c464;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190420c9e3c4279ffa4ff9f4a04ff0bdbde7df98a2936fae61dc8b092ac55a29fbd5ce388;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7887a6af5a90196fa49be440109b00bdcb88f6559f0a3d617e9ceb30fe3a3d94dc4420;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa4ffa6ec0f0dc8acc40d346af3c7eb5983c4be129adc48e0a96d2ee7c056654d93b1c58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ebcb9ad6d52b06dad2e8b71218d446a912d60aee181fe2a942e8be2158b4f5a7aba49a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h918baab6bc13a17804592c4794d93bdfdff0a7de85f2eb362c39ced520e67a9528c26c51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c4c6b3b921df4f851502a83fe444021e7f4b1ff09d684e77336bdad87b8cf32256bb734;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3d45265d135fec2bd9f98e4eea703747bb507b4406c5f1531beb1073119549b8aafebbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b4c9f9e9a564c0363095292c2d735fb71306df43c9e60cd3c783e70aa8374a3a70043b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e02873bce1dcebc67843c720549f1b12968ec01deb6dd7d52f38fa611e8aba1239ca297f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1e4349edb163014e4bb4d75e7e6cd4f4bf3b5ee554ad4ea3e94274d2669998944c383ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166b7b45880c77a1c1f2b6aa63882cac59bbeb51eaab79817b158f63a6565e2fd12b1ff9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cce027216225a68d87da559e80d092c3fa67ed6bed93ed258dbb145c645de968f91fcf44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e50ae0552a0f30a428f814ce514b02594e49cceb69b5e71eea60049d3422030c3302bf21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a60c435f5c7505480ca226fdd692628efad204369fc183c6c1cc2413fe7c4239f4ff39d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfb041bd04b032be70727dba2c8828b43a201127c7179020b0bd0b115fce44108054a64a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cae299e01aff2e0d672f1d3c7e394b99c7bf1fb8c206456385e2a6bb0a3b2c5117502b21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17da52dbbb47ac7ea415e387f2a4e6b879f1ff6b496ec574b59a61cd5d3ad1422325f5725;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2611ba7f1049125f14587f4d09f9ea22c0875f3b55b3c29690fc81d6cd7bedb85000007;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h892bcd67c5250736645e456d236b5a4cd53a77c95a30ed72224382adc6ab8761e367093c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6d417137a16d840980198a3d9768d64d0a1c308a5fa7eefaa1069fa80dff4b9462a4576;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188976e6c308c08ad473da6689e8615b414b980e73a157c3e91ece54e7f1481e637834cea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b8d30fd504428cc194ab5ca9cddf8fc2000eedb219283a5a7451c8561f30afc58de696e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0bd86fac1b3ab3554db71c7f49c6465378ec088d11985ed430715037ca2589cb9be2fbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181175a86d66e78423fcac892b3bd783ad981aa533b110e5272bd68880a16d2da016cbfdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da091d754a6d03ef7e6b102e8ff9305a04925fae7b3225358655d903b797b484e8bdd8f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69539cd9300c47ab16baa21bbb4a6a1e97cb5140c902cf4f2414a13b6584a520d603c117;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h434cb3aaad87975e687dbc1d24138b4ce4e88f3eeaafb6dfe24c2a5971f961b86ee30f30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e35f6348490c8e994bc3d410c590a42b8cf2a2e7a9bf17ae2b29641fc50f8801d4a8ba9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100d50f4fa8eed6ded0246e4ba712c31da70a5d84ebf4c34731e39a662c27270d1d4f612f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15cd0de616066590b27f5482c88af712413659d0ac14ac48961ae3ccb6ff36ea23f4380d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec50af197cd96dfd76b36114c929363a6194a3ffe641977862db81a01bfd550c999e52b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c733d7f1f320004c0711fad8625b8ebc45d32cbba21fb802b2d30f58ef1aa9e2cef84db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aae46775c0975ab6ef12ea8340d9d552fa58e645af461c46f7eb089f4f374e8f970b8543;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c8179c52ba811e887c15ae6ae3846ef0cc68b20e78273b9cd84911f417500d8d7f35c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3039d5b6820b6cf56c85a8638b66507912f2773518b75d312348a378aec92a406c1e7d7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbac2af173db93689e9861f68a678074b638a6d37b7b0ce2ce35d184070f001f6c662f206;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0c0797cd3a32a776f444a77712e12761f01991d4004474f9ca9e42b546f7c7be5208946;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7144db2fc573267aa4fc6456bb8434eca615e460e72cdda0ff938365cca1254f305bbc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98c7692f9660bb4c24154cf0a2f48bc264ebdd9bf3a90a365bc0c809682d4d2cbdd26e8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175de21d6dfa23c4ebf265fbcd55d65d43ca85c1e36618a34955e39345acc0e99d2277f50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad47dae67ea8c3979cb03d93a96895422a4b04ccdf4ac0b99e0a27b6fb7c71a140d4eece;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dc4943dc1c43e04e11fdcf3611fbb97c1025a9961f5fcdc3a6f7f2a08a27be088a6deeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4ff6739c4930c7dae127e1a4b7f04304a75ff2fab78720ca1fe1cc88a5fdbe4977a3554;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4a5b81c3ae47f9375659b54ef3e2aabbbf832947a88fe69f1088cd72f921de206e7cee9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2c629974b42097b35dcb52d768360128372af95baa7cde879e41ae2af8e14327e8b14b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79eaa608d5473f3390ffb617737f51ad4957b9a0c3a39054ebb7a08c1447696c269fc274;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd0774310f1ec75160416975c06ee4ddbdd7ed2302f33d370f25e662f98fb2c3cec3bf15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132ddb1be4a9e9009803fbb404d55e2b339f5c22efbd399a6bdcfb8120125726ca5a11fe4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h983c4e24c88d745c2ae7c54794b05824ad0bb9d2f5c8ac5152437ecef6bb30db44956fd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b06a879630c76122134a7872ebc14aab6536cc7705c9442f532c19479f64475be03ab5bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ca66c7f96b255ee4a001a4fe91c6cfb66dded52505a6ce7874d34333f2eb76542fbe530;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c73d97b2b580413f460ba6922a8f7790d8893c3514c54b3c1c9ac5bfcbe6a5c085c3298b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7d9a319fec85aecd9a7b566417501195a6c316fbf7bff7d6e64f7a79109cd3aa2b7a6a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h589bbe34334325fc225a063b0e12badce4fdf5f225f6f80afa3691a6ebcc17353e8a0c41;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2813672099a5ab2635547eac3a8833a16a98e03443fb1e84456c61326a4ea5184f1208f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3142e2537bc9f2a178d2d01fe4a71a24dd623bf0909cecb2022a877c57e0f2496d7d3868;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24a42f1b4a030230dad03d75d9e73bbdaecf260f170e8663e01f894204f3185784177bbc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1027df4921fa74e2e9aac7666ca71fe0725b648a10790fba71e35410f3fd7bd7b05d031ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1780f964401114332e67ff7ca55cafb860f916335d22382f9dd40eecefb5d38eb3cfa9b8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172bd037c15c80b9caf162de6097c00c6fb85b5e818478b9229c11924a1c754596bf6996;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef354a344a8efa287ef8aaa5e87a4766988dcc2f9336e95cfdb377f7a43ca7ad2f93adc2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14be22c3480948b46734425ec7b74e70236159d6861b1975f078cbbf05d7e04280228bf31;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ac404eaf89f71f1a468697eda98970b8802a88d3a96e6c51e399f42bdfd55d01c7befbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haad2ac75c177dd36fefb01691c50d920538b4b8214bdf215185aec91bff0d16b685d4e3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b47bc4ce804f2132a4115fcc789f075dc2c9bcc137649975c3d20428ba9703890524456e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175d8a02a8162f9088251d2765285af7b8e56a0fb4ea0690d268c681d6576ee54b6a5adba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18459dab79b8b743568ed4b3711d0a1df1b1adffd9947d88ccf79fa13d95bfe62aaa833d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb55c7572060aa11afc094cf670259f96ccac97c8fbc803611a821db46647f095160e3673;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87e574a295c0779420767256ac4dc085c6177c126d2c296f656cc00162774bcb3a87cea9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda08c2b0d8a294f54f40e4576dd2ae0f9d8815441ddbf3a89661506437bc80f14ef8c72b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf927d3ef1d8f7f65c655e1f427e08ae80babd101a643848a681681fad11aa265817c8d95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199a4efcfade125acd4387186f7fba6f660258c2ebf8f8e321c38ab4f899c01c1a078b2b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113c82041546c9d7c41a70841417f0435cc49dcec0ea29e5f724ed1a516daf9b9c39ecfc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbe82ba6990a3aca7d2665f02c1bdda817fa67d79aff9e1d57559f2045c7206e2808a25e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe96e0e3eb996ee5bcf4e264ca46f71bf027282c66e2369c5656c609017befed6fb6376e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he08e446ddb5de8418ad63080f587b83cd7f00cb5114ba9ba47ceaa48e594acc9886b8641;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105d262f71c3f64739b8a42cb3f45ba1574c8abbae3578dd24018753a0a446aabaaca00d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc739852ab66ba5ab51e15efbb9aeb3844cb4293bab92720902624609a1a04f3dff853970;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8525c07300636196e230c1191f63b602267ef1e31d57ba9666b48e53b2eb438f347f29f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149da9a40731b35b0877bc1972c457040a99f6f320dadf0a72dc2fecfd53bc00938410c9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b5f36192fc1bd77043e9fceba1df1667957d5f5cfda3fcb4b01bf6f0f1bf3eda795923c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f66746cfb919bb3c774a9b5d6bdf694ac6a2f55295ecac6578f5cc00862b3bf955fea750;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1802da560f47679a9a3dcc61b6aec4be3b86b60323a2e0cc2b977e65bc1453e62218b440;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147b56f0390513f08e7d428caf063e37e934008882131a7676660593f44da0255378195c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf51e94283aa3461a781d5d648c358e587731e363390719d597b403e1ed4f75e55b839a88;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d5082c5148b837e79f4b11987cafe92d8d6b345cb6c885e49611ba52b0407ef9d4588c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a42f46de571cc2b284b69e1357526ff81d41aa7a904f1e6b371358037877d7300e67648;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106f116eced7f913549e948b8bf576817bfa6c82ffc36a7857a4c40e9c30a2615e10e5e1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e67e497d83f9f9c2297c4be40301aea07f3301d9ed35a116138ff0e2757995ac3b1be4a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34a648429ca504dcb62c9f99f8419071c5515f356af9ac2d44da498b60e63ce933131911;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19bc7a23ac552913fd12782c0920019362bd52b21e0486e0cbb7abd80d25b532c9ef411b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18459a15e0f82df98fea0608fde14171e7ce5547b8d11bd8ac39855688cc4214f59c4b876;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13890b494d6e8c40d2ff31787d733691a713dcd19fc270211560bf0ca6afaabc883f9279f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13132a13440a4beed24492893155a4f33f5be29703af52c7208490a4830e26bce6318374;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ed21fe518ef01725817481f614dfc508665278a1c6cd1ca4feb119f070f906b0bab1978;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e60e636869af8e40d1585e2ff2147d5d784d4cbefcbaaca979d37ef824b0f1737114f5dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a191e241c9ff71991332128f932735f13b0841d6f1adf78c0ec075700dcfe88555e07318;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170455a7d5ef12326aa2eff6b3b0fa6f06697e4b56d4a8378d11097348db1cd0ecfb3e067;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1debe793a9df7c04203a8eb57808512c2f87728aca0b346afb6038f35dc3e3188c43d0cb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b0e81ca0a81c008b652838b361c20276ffc1f0cca0f77ccac32f2e12fd3675b5db15bc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63e5cb95ab390f56048fa60c389e1e75e26e068851ac33bce3085eaa7f17847fe775a04c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7cac502c6ffe8c890a9536c499072852974950f226cdd78d439e6ca1407890ccc46d3a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f1d156f0c811e23774d99fd6bb76b391f5f5e2f58855a1d194888ecfef0b3289e58c34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba3ceb38bfcae64abc17bb9ff3f507aafdd211ed9b41efff152d9b8ee9dbe2088aade408;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1cc90700258a16d5fb0508b23090b68fb132225b0b07a9c36611fc93444d4b53ba373b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51e71cc39c9976ee3dc7f8199bc8bbfee35b66eda89dcea82c10a1833701c33ad807594d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb153d64e36099200f6f468f56273202e5422f6da936eaf8478175ba5762143008a7fffc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ec5a3321a62bfa7b226f7d0e59df68ebcff65fa1a2923fb77421b10e56a889d27a1c5e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e84c1b2c4d877f7a4a88cf116b5c2325928528a6ea81e2f1afa865f054911ddcfcf826da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f694c4e6d3cbf5facb0b13fb3e52d2c3a87bed2aaa01d87a61e1789358fe5b57eada638b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125867f8915e3e8e8d5005bac9db2305ee5faad1f7481cad85700894e6aad5616729234b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d460c23da7b9279bc111c16b3be6eee2858ba51cc7ba84f9d584c78b9deda0da5f463f75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafc2b0d3c4b9bcbd2df5d46f3419f7f09c20a1edcd5d4f6c7a305a1bcfc52a549e4b3aff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h458cfead65f5142f4b389405db6e3bcff89689ab57d1533ce44e7d4d8e81df48ad3fcb55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d2859795a1c360565bec8659f8b3bfb177a85e6ffe0ac1ae8ec7e6b2fe1e4a01ca9182b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f07fc24cb9cbf27ea16674504b0a6500bb8fcaab0fac6dce2e407ff63af018bc13e59ffc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35f0caaec4d7ff59521b7663da3fdab7bf2090319f5b554c5beb7068c78c6f29895e6746;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171dc75b11762db8bbf67212ed940819e0c878eda79e47eb7842ea99df71ec52fe13e077;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1956d842ce6f318f8c4ed9d4613140b9a522d02b0ca2e199ee24680946f985d8c186c17f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac9a355fa21803c7117a3dd4f2f3f8070a089894a75d4686173ff7bb1a7dd859f083e3d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fcea712155d764c4075bb188d2dde7ce1c0cfe3ca992afdef32a1788941d46ba5b28c84;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82e633b974e151a5e45cf73ade7aa0c8e94a0aa22fcf67cac8e42ce0d3a0e39be5c3f05d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e9d5c8b831bcf829037bc236d6f613b013d1a90a616892b37c6bcd5a207808842663485;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169d8ad3a76eb0fc0fd7a9479725875bf81b4aee20183ac7ea6040cb06a8de553d4073b2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a8359d939b101fe961e47d08b415e27fd81667a49cee743eead7f37141b58d2d39b7de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da46fef14a38cc32f10a88bbaf8a073ac7685e44727a16d8fa1505a6ece36d46c72d574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1824cacf623b296a0c70869c518aade527f57b832ea24d6d9c6ec8d5f16182e186515d5c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f5d1dd12e8be7a6d72a4197580965bd684452c6700c80db80d859191ec7b557239e39f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18130f80a633767d08b4d8b2e57b5a36ad1933dfcb0157af89fb45afd39ed0acfc31c697e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec93a1729b5ad404da5f4c3e9a74f97e28b69219c381a98862de75bac77a32bdc9ae1092;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc98668034221ddb8686890887a8cc73a71b83bce65cfd464584a2812f067c17f3767de47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc54cfbf9b36bc4fae8656d75298eb41ae805bb9cf0d5ba2f54aec6733ccefaac85141261;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57088568dbc0753c8abad813557854d6ebe9a4295799c3c00799c24a2457eada81c8c4c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9517c2480446e0e9ed1a8c5d4d103f01d90d074157d4d2a983e16257ecb594ea08927d99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1caeaa89c99928648a849de2524c1c88aebcc235f3e0ab0c559cc9afe9d38169de3467ac9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114c7b0dfa379649df70448dac735551763f9bf266a59b1601200af81ff7e0a1b31e27143;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef40d5dca453e34f28139d31eef431992255ca74d42c55c2cf38f621dfe6ae48cff2be99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193090623278e911f78baa5512274b920845dce13ce66de53452674f86e478b8335e60c53;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h395c9e6c50402304077fa693ea612b0757b976aeb8e2e14e731a1625db6bd2cfc2e55450;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159867625bb61e4498eab97a9c3fd1b69d68aa817b8cb80eb7d5d4250a0b3ff35b9449cba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d597953a16a7a10fa1553dcd2de5687cb87d5e573e318ee3c8872a8bfcb750d1cca58e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde65a58c2810ca3e874514f5b017c23d4e2481a9097388fab14c68091b44b137280f6080;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c905c0d1b885a2a12ca7728ff44a6f83714800c50e30eeae75012d992cf5edf76b44f00e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f3cb6a0b21f985643dc5512ca402c698e8875c6bf006f9d1b5920a095037612dd67cb60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce2f56952a6e973c99e753fc410263f1552faa6ab69d72a720eb4eb4a2f1d85b7cee88a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef9bc948ab42f6bffc306c986927a90ccaa9590c0169aa6627b74ab7add5200be6c93c8f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bc3233ae2e0a867f391fe5ec276f5500b35fa725b59a6fbef00a2dc8a30122d228fa2e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57e5a8cdceca402ae0652e16c2ae285d51b4007fe94dd4ed8a7219844f6690532f4003e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e42582151587eda36207ba71e02e71cf6f358bca9b8ce1e51deec333c5a2956c2cabe61a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e8bb904d4a9afd5c82d67fa088b67195120fa8e735665a3decfd552246e260b5d94ce3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h798940c9ce420da8a2a651b4a072176af72453d32937cb71ae0298da7acbf33c53b55a6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7ce0943e68b8e5edb965d6eb77b8719ba6cd89d51e215112164e6375a9a35915257cc1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf34ee6603c9e8f34a79ea0e60881ca6f91fdd55b536a25a1f72f4581ab75b5b2dda00232;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95d6490e3fbd692dccafdcebcc768507428694f781fc86bfedc9e384fddb13eb13f4b9cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a60042301b039c2ac25c1b8a8e4915327dd8ed0a5b5753941fb7230bc827e98bd3cdc54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d4f71d43532ec32d6c68eb497d648dfb3fae4fddd15fb1f96416524fbc0d9d453956f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h711fc13e02f8201c885caf8f003987ff959bc5f6c01835fa7c51b3278d8cce1f1555fc04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17407138aa05b60a13d2869076c9b4361ce87aa3f567c14a3d52250a3c991c3fb56f01495;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1353173cbf6d430494040fe3edabe245a9101f8829a4a8548f17d1109068e426ae9853772;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee5e20b9f8cd8208c79342eb8f91e2d234db42969b0073764af7ba41c81bb8fd02f0b0e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44a9c3ff27e77e3be854010f36cb3513411805589e42106e43b9bd28908785a2abfdafbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d27074abf8b4446a8de68631b451347e9093719b4895f29805a5b279885d199ba1684737;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa0cc2905ba7a63d2a4f6726472d10d7bca67293301d371e044572fa662d473508cd2ad9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3aeeb59f01df15aeabcfea19f5e7cee112c47897af3a8a75d9d9693804cd30f9953dd369;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1363407928bfe70063bece555c1003eca278eec4f52710d4e75f0726cbd860861a061a942;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1979d0c9e0ba3c1cad22abb7df1c29538665e34e19824a774b48e02bb32a2b895050a9c6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14655f5485d3c600a92421fb0a50612f66dcd55dbe155fef14b43cd4d298bc80efd99be4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf2b13d523419c8a44d25aaec11cf3e5a207f2bc6912865b96411294c5d6c59b5e8d9aac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161b263457a2b1988e9f6631bc77f56d789c342c058726f35c0d98b7c3fd4095c962ad8ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc87658d40b5784ced907d7ce00c2ca242ede1337e054f094c3d8d422a5e4ba41345b9f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d4b137e5670e9a825f69595a09312eb1d92664118505c7cc95fe7aeaeaf1e9649602ffa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2353e10d8b3cc246133d9fc7a63f6a20e9f592e2bae2a8ad16e65a5acc789fdf1f44ac0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1939a04a46364de92620502524371483f92e05bf26cb57fca814eafa33b8bc7f5ad25870;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0984838c686b25ee2b79095d7910054656dfca408eab788ec21ada9cbe46a9fd057013b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1884ff2499ac67be6ec8f5130d7facef43c633387ef7f23f83ab4dd320ba47a82c2f30daa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h990756aaeaff5345df3446c6f81d9dd4104f5c27ed8cfee34ef0a63721d59e1a996a57dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158adeb95effc2c3dfb45ac1d1001afbef015cbddf00f68b24688d1065f26c48156af5afe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb20875b522e5aabc281791d169c85affff68ed5281632ff34a48192ea0bc7abae707811;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dfc6dc71e52f1c04ca7a42aabb9a332f29312137146b83daea268888e0b567b1e462570;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb90481d3430b93df73aa8af966fcb887588428e5cf10995fd60d40ff1b6bff9155f4868;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30a2132da92414543d396b9dbff194e988c19329598272dc486e4a8b38d5c95d0fb1f91b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb8c8fa0bf51e873e866d11880a9822c0dfc50c4668c9b9dedcf0b415ab0d1861fd292d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc58f58d4fb9882679e5d05299d39621d1f110a8c7fa72c74e17e8faf18ccca520b2b635e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heacb45148c62d2fc46630be076f97b15185f103524b204073fe9ec568f7e05c1609e338;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3a80b20af8c0bbb624251bc1e6f5dff898768d66172ab6cc292cc517434e020e26d3fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d329cfe0e9bf300dc29148ee7c10e4223b2fc3e9b25ea703d136ada9ef88ce1965f4a00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10191bc9522affe4fec72815549d05aad3c77faa94c7fae60e83e36c689051b141035e86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6379cc158d72b51222180352b47f67e78bfd67bc1c69ba326b1dbda7f27200316409d90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f45106f23754bdd60a81dc53588359c46743da4ce0a3933e645c4902fbf252aee9d36e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8959cb731f3a0938b75ca4af7bb699ac3024cd4a3b99794e485ecc3426200f70e80651d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c98345902fe862e8ec5ebbea2415e47dc2eefb4a3055c3888c6d309899022aa1316d2883;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b95ca929fa50141c66be171cd15a263abde5bfa049a1d1d90e03eb7365217003a47f75c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e511ccb6e56fa23eae654c1e6f65989b1d3b264a8661c9f1dfe085937ac98cc7480b5f25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57bbc724f28dcc5e8eb41a949c3335865d90a103f1d674c2f0271f8a83c64f3fc9f40a04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b4fca7f8a4c5871b98c10dabaad0130caf5ff478a741efd904824a56a0a8fc9000138b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13323cf8d1ddea5c29662c6a9463aba6c529838a2faac7ff8f618e87f9dd697c38996d5b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5319c0349a04ab805c562f282117751f7813905803ad9feb09f8b2343b5fdc0cc5b41d29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b76855fbeb6b0e471d448e2febbd72debad8c6db0840f0b45396d234009b28f3b2ab169;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110a85daf80883a9775f125021ecef442ddcb1c6c3e63f31a9261227b3e805aa5c3979a4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ac84b42fbd0533e6d1eecab6a60d66b9b0747ada87c61893b61104bc9f32d1fc3d9cf20;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecf602d6ff2bf68feffb630aac18f717ac96c43ab097a551fb5f98f6455b7d062b9680e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10426d6bd6bb56f41d6d21e46587269c7b0e89d9329c186fc08ce7716c005247cf78ce2aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb9c10deb2c4850e7f23bfa05051ffff3ec35f06bf8e7df43086d928fd9f121fe3dd65e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c2416eb070040a305c8682df8a2b134c5dd7b2b783e16f2d48c5128be6ecb60969f144f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd95534bd60512cf3f5c39c5bd09a5e006ec0160170f3c674a70d60ba307e612c47b12374;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6fba14025cbb254563423c71d028d6b1a2fbff223c72c620f1bf1c3b2b7eb0ae9515ddf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa05f4a113c5735adbf38b77c254497c6b3e5db9af08b4783a2d6bba13ca30746d4f828f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3db6f15268f8877e5d2a00c7f6654084be32a13c3f0d5dc33e77043d4df474540d5e3e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1347bee56702dd291e27f221674591cc66bd566770ba124c311e6a1659e441c97e16648c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f071026b1cafc4619d6569da6025a999dc04e823f327a4d09d452faaf8f96259753f6a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2d81030fac328d6844f2d7229965446698a6df74e8ac226438787002119eef5876ff41d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdaea6e519eaf252ff074e03d458bbcf9730b930a3bcc9e36511eb27162015d5c23eece37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5e872638c640b586bc89519bd80f28ebd4921389507ae2dce8fea276042c7b20c3995b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1c336c15a79c81f220c60411bf57780b843f0fb3c8a1e9f81a3f5c922819652ab324f3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1d8122e3ec8514c48385584e2aab74c02f10cb526b252cc27dd2730f1d13cf3c413552d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe119e5ee133f47825b2e8c9a82b40c05ba7f8ade5f5e970e132591f88645efd65dfc029;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9daec56c492589902c553b3c88cdafc32c7358c49df84afea65dd2cf4dc5b58121dba639;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3445eb1c118fb02fead1db6dcc435bd89d06737d9662a3c05818ef84840aa78a5927b96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa22d9a79d27d82005737ee1a4a7f2c98f11119b624837528d6062afca7033b333a696e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e56d04a46c513cdff4f9395b900b0b8a45f671765e4dd381a55f2cf2cd3bd970a6f427e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ab8e1dabc67d8e9f5a7cac99652ef9b3e25cde1369926cea8795fd91a7162b39c13bc24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe137035accee57bd3d1323696f91e9191d1438b907c898d179d63c05966bf6f25ff40f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9666cd579127557ae36efd6298f4b959ede1acd83d94870d64eb0933d021cfb0e045e788;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95fe495fb0673a407ca5224aa3137b125f996d9c0c88e2cdb0ef07faea814e636dc3c86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc10b7b89c0daff633c8152f943891d301730dd3ef9b7cc2e699a4b84bbdf5d2175dcaa2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1573b6ca7d481c8444503c67d6890ca6c1c4b7f9549419fde8574458052d74a87c5b6161d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac6d7a02483615bcb7d1dbf978f41b3e0c53c1e64e90d3a7af2a6b023e13433f4db96a37;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb63aa697d47663701815b90c42a3860e66e2e500125c88aa9036bd2f39222a6bae15e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c91070a90cedc494446c12173c29585b65d8fa4ef74a14557e285a12aa596c67856d90cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac5e5ad87c60973b65eaf10469dbd6bf5d1273580ab6c53a71a1b7123f0668364e920025;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef123bacb5f1439819c1463d742be253f45ff0c7c14382ef20a0eb3427b064d02c3a2542;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8f93bab942bee911447d208fbef7544813fc064d4a0c5233829ad4a8c06bf7b42b9032;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51ba2a257f978288f5020e390c4ff89f3cfcec9f26e3f9ce89701468927f2477629b8d90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd06171ff8a03962a6295010a7ac15a19fdc8ed08e38756ff98bd860fb6b243fd9691d163;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181c939e23c810f9453d79c9946552f665144cb9abf455b58b33c9a805e4ee4ba86783512;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc4fae125b5f20f80bf00c0be2c5fc894b72feacbfe576190babadc88621febcbb885623;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8e96b30a511d976400af6f89480090f55448c40f4cec7887eda2d01eca1fa70ce8128e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e443f3c0f2886315ddc52477c434c124b552b8ca0fa77aa5904a61f991a7ea32df160df7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e8b5e028abd5ad20030910204eba7b567f4bbf5c16df5995aa86bd07ba8bcafbe1b54f33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc874c26354e7cda4c5e68418eb8bfc1999777a5aba75e359a1da532b147c9719ba69a3fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177f65f34e245f24550d7b5a2dafcd1abf9da77f346f2adc80b53489cd81d118792f62c26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1caadf314ec85b6e54b6e67ac196c9b3bef33e396a95336588d25789ae8e4ddc7a9f70c62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1027de7413dfe563aa738c5045f0f29ba451feee92978dc0ff2261241ba3d027a54cc26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ffbc033230860be6362e4a8c6d263c3c4db77de0b25dd88c8d88d2510965ff211578acd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb37d26fd6233abf1f8161ab500092978cb89cfa26a339ef539501b4ec7c41b3bfc64b53c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h656c4929e6f6513f254f7e95d73ebd00afec3d158153934a226568b22c0109c3a736b53;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166a0ff7c53887d1540bfb71e4240399d1583cf52b6020bbe2067d0aaa43cf526d0e1dd7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42b23eba57e91d6534a7bbcd19828c40a251d7b92da918651885d9b3996ce53bafc9e19a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149ee1f3f485982681061f4062a9c4b307ca7dbedf054ae473ed5736c3cfdd7fadd941b8e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c1d74fc0048f660067c83331eaeef6f75959575b4e86713d542ede9d32e00c0fa689391;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he52ac06c6d4ee6173ce8ce8fc23dc175bd668c89fc19f62e9cb018cd37507a6a1ebbc6d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5d380efdb7bcd4e8c842bb67f47ff2baf717df5892cb77160a0014574c708d4a428331d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd34d9c5afda3deb0c8f658b6b2677c06020b5f7d567ed9c74d7a9a1c43d9cb8090cfff89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116b93478330df847e321ca7740bc21e9860594249e076f4a5559c7fa73ee2ea5510a17cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heeed567b89a8639629fd0c0669bdfec5839149e03cb5bf9dd0b371ad1e29ec6da511621b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85d6107c6b178054fb64c8ea406d82d22e79c051c9ab127d1e73ac0922e27b8bbefe3407;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190ce5d4474d82e5ca424bceeca2e759bc5c841177f8e4a2235c41ec92b9fbef1efcd313;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8497f94ffceeed1ec1202aa34b2369b1079742129075a143f840d10608950a2da5e3f4b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb4da9b80d191068920a68c0b7beeee1cf5e8629f2a31fcbe5dc1a899a2496af3c503a63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11db09b39e1f890a6c856b246385ce5dfaa7abf647d042e6143345b960e58daf926c97c16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1558fb3497d95bfd8b7b8a24552e5f31a01cc250530d253e3a9fda7a8db09fd4a855714;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac798ee12b42bbbc95cd65b45f1d65bbec4ccc0daa7eb407e718ae0b47ef6dc084fe2880;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b6d768572e968c01b06e30019d5d7dc8eeb5fb9644f57b17d625b3148dff7ed12830f5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11053315e2d81ec04731af4606e70ab61e58d68f5ebaf7791769b20b21adc52320857cab6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6796d306da8a2d292108396b4757fdafa720df492ebb8ae42333d8b11af255008286cc5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a8a64b5b1d6ffd57c2beb405f8ed8afe1ff4acc97e2ce22921aec0ee40221a5c95a1d98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107197a894a82f8df2c6943dc54b4857b36d3a9c73785dfba8ddf8881f4eac8c32401788f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0b7ef8bf78730168156a63c06047d9653cd6055b572c134ab988a29317de4ad12bb5fe4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fb8741e0db693b60c39cca9db4ddacf37d8842786e3dd2a39a54dc1cc5d2bf6fcf2abbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1700622bee4e40765a3ea9b4b5e0c031214a182af43b049b812590f8211c37b33c4378a93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6bbe268d179fd9eb482b57f5a920550feac00ffb87f5fbbb1df21a04d9ef7226af2bf2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdcabb527fff6f87dfc1c9eb299458cc233d261183a1e20e6501e9a058138035c499bd45b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19744df9389f745c7c195407f159f395953363476ba702cf7f9e3d38990b94090c11d6e20;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b20d6140bc389cc2fe9ae43d361d7cfa9f0b2ffc0d028c1f2e79c9d4db36d9ee0c39c40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83305fd4fd7afc79efa510eae5a65d537c3e5f3fedcb23e434aaa4d97b833bf1903ccf23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116fd174f25b877f6c7a248385a2849d812c9f0fd472ed94c0062d19cd9b1d1e5c9baa1b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc69ab368f4d394f5a9678e03f9f372a4da242172cd53ef9728036cbd17c698ae121957f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5984d7926f1ec4e3d072f43484ae07efebc8b603ebb754ccfc08ee7db3397f8e54970280;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b9ff93ea8beaf756687cb8308912cd8578371f3184b74837123be97f60e08dfc48c19f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e2eabd84f913078acb76fa27d57935537950eb58be94ff9d34674cc016f2ca6ad19d255;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18cec9855629de9e3c6367f70e42d093a580e842253c27cc080c73766dd3294f07167655;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd29f4f8dbc71869edc496dba9c769b5202e3372bf9bf039337b4c7bfb1d31bbd96c3b078;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14211fd7349ef11cccc46962963eb8bc971b97892fecb4931e173e11d1522d73e9437d3aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f4f9b4d4bf40ef8cb2f1bca321104e4f4f6549cc24f92ee94183b115918778a90157cc1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150529b0bbc875d108339d5b3ea8091d614ee6be3f0181f4a05cff7202e7e956c6fcb97a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h318748309f8fd254eee43335d46cddb07c44a18dbea1b53e36952f8bd68f12921f8772f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b99757e823d4ec784ea3faf04bb375d401f0761634bda8482bd9452993d56299e603c1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc04a19a93de303ae173caf5ad5987143b3f4f2732aad7086ec03309b39ce56749ea2bf5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184dfd151a6ab005e96d8cad31af0e2372397b27ae8842eb0accf60b21114aea5b0132d9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74df85339f727810cf0365e08c52e452bf6eef09c1ddc0e62cbee9c3d566913c026ba97a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8255494b6bdba6caf99b3e6a4a9d37848e07534a6bc8c950ad3eac71242edf8cb1209696;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbc58e7b822dc19a0fa39e37a5cacc68ce7e488ef07602ae9e2bc8ed6b6adf669efc26da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c338e11a108a1362071a3fdc000c1007abd8bd9e46438f59b799fb3f7196e646ab1ae726;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9a1dcb3e66419ac5145b977447a403efc816df1356f3e7781aa68bbce271001e5d06c6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ee5807a1e7416a851275b7885ea6c665c0a1c512fcde230294af56f20c2d0f6ef52eab4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e8b9136b2479fcc484b640f6bad839b2198b40a87e8b7f18ce27139d2523376564b6df16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b7b7af5db69262e4637205755f70fe142365d71e03d10fe18b8cd9da1ae0317e9f4c82f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189de630ae3b4fe06762c84772184c7da5aa067492f5fa096d81e04522448eaf15dfd4fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef8a388b102d39e45c4409086c0b740afdcb3946f159c6fc979230e129a39e5c32ce1c42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26ca0ebc64fd395e4a9d88421cd062829e8b8e4843a60afe2c8ccaf6457dd034962f4378;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96b4e352c74df4ce13c06dbb57a6035b85c63045dafa7c507f6edef7e9955c98a26d0d19;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cbf5ad889466fb572778dd82c2647d3919bc4cda7c41425b3a4050e09b93551478b2ba2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he203cb6cf04d35dc032f46f659ea60b7b5c6924aff390c62cf692f5e35e125070538b763;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ddd68c2859ea1ea9ccc03a73548436e67e371ed42958596addb958dbdcb090ccb44ad039;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9666cb85b06c8aaa03249d8638218985104ed6b04395dc2dcb670228b45cddef9ca8691;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8dd037ddc8b94a2e1765dfe79148570b50af43ecb8c63cb4b2c52accdc8d880c9a8a2394;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8835a42da892e397c36250140b21c3ba5bbac545acb1527136b9b23cbf07bcd3f82dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155cc93ac26f3c0a2aab5edcaa10c41e19583dcdff9fae6178a76911b3e1d57cf226eb523;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ced7efe2971e8dad956b2faa954fcc20c5f53d075b5cb59e2dc777fe879cba3b848d3c9e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a51a38d4cbe7a25576382e95c4d6f6f349a760282f7c352b897d8b40fa87daadb6cdf03e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1779a04916efb0f2652eebd816f7e2a7f50fcfeaf3b02b3bf74c42ad4d8ff2475e1c403e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc545ca986dd2c24cbd859f3e7219243274ca15cfe648218e8b533bb0d810365f30847be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9c4ec6216036a18c8c225a8ad87497e029bdb56b331ff6399f9553b81f1ee5a3e4e30be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48d6a7894f2407bef79abfce83ada115b64592478f943d753ba9bf2ec2d22cb621a2ee4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ceeffa0384cd21925d6c7704da4fda16bf543b37d6ba1452d2be12e55ebc95eb4d0f842;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c0ab9f4b5a60fdd0c1f468fc78f8ba6a021557cc0e584971a62320c86d1a0d0ced504ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ca70984f3297be551437b560e5d867aeb26d62583ee771df587758f38b15b13ec73905b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h274e1095ef6c968114c22c6a2d98119ab4a8f36a1b5740cd30993fc48d03feb6026b13e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha563f3a659b5fb95dedde9123e684841cdffcd5c1df0764a76a6a8bb41d2a5b4fcc1935e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e3784e673487b591e7bb059bea537e01fa83c47213a3e95a40ed0e2f8f4d468f2c24d50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2eb2e9b50de6f04028a06b73016271911610efa894f4ece4a25a3c3dd120e75a5d2c09c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9dcd3ef327de305c9f04c0df9442b1e5e189958e32f9fbc05d5f96d3b583ea054bacf01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4921dbba5f1f5ee01d546baa51e349c75c8164ece037c8fe0c46f6af5955923c385a343a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4c37677ea2eef1ebaa67a5340e24ae94c115eeae67547fcacb00186df38f3350b2defaf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc0a9d895974888983b5e14f6dd72cea2d1f3b0261a96982a2ee69f1127c654b10c8376b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25ca127c1be27025f581bf7c3f9824e21584586e7b17708e201723d7399ae1d490d0eefc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fd1720982a448f7d95190073b2a5e17ee180b7c203ec46a9fcf881562f3ed7ac9067ddd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195f973561f2f03f65279d065e866c784d626371eaf21fedc92d547831479b9fd174c8696;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189d8dbe7d94e8ffaffe6323250c7d13402b36b705c0aa12cf9f55b3c67b25a10c88ce95a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117b6d9244dec47e6d0dfd8e7536f27bca58ec85d0053847471627b88143acb9e663f653e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c0e1caa6b50c90165320c523fe30e429d1d222af7842291a56e54df2388c8e56da8e100;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e17d189c629477bc8c9303b5343aa3d747a0b2a04e3c32076ffa992fb6aa9cae4d81d93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fed7102f3ab9615784e69f08c4d265446825004f7b6b1dd0b814740ddd3bd7f9f515a8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b859ae9ee0add491c55825a05322835afebdfc3666366c285cf1f7fdf863a9267bc6ed2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66480c77876f829307550c7b01e5db447d38e9cd6276140e1944c8092a4cf8246da0778d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51a78ad28f4af69f5ebae6edf7d319b911c4778acc41b4187a96ff9db27d46d600c0c062;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f03d1dcc0bfcc5b000d3cfad419baeed589aae8c6a3cc8bb9c009064700743af2ec9874;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11abeef552661a7587a78ee4c01cf8c7349bc27bc4aa6d4041fc694dff04f9cbb9a0c5861;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177d141b19296be83cda3788e3f1c01a28bc732eaf0e9c764c9bd634f0978c9d154f7fe81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14048dc700258f1f49b17b1ce980f31bac4dc65ea688237c12e3356288f0a088e9cff9ef0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2c40da77ba71bdee69ac2afd116906b1781eedbe8cc39faad4e711b8d36d0c8dc847f5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cd49bbbfb4d8c03619d3227f0780e64bec7d64ab331133df88fbae487896b9ff6825ea9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b3d1e70fa36fb88287e267ce81d9fc15fda1d9881c7833265af351320d2a88113c262ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60c09d43a91c52cbccb3c3fb4da2bff6c5c7e8c4f9f80eacb943f1ece3960254eec18dda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b42b3db4f8c076cd08e89a56ac53160af69c32a4a352062f7f22e1f6a94b591a5810a2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab58b0572c4218d76a472e8e8cd7c3965ca1ff62d675ca4185fbb08b3df867c7c7cc9d65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51ad39461e693aef47f7e8e9dff91b606a295ed089d7cda92f08e039f7cefcae3426e328;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he074b1852b7498e16740f05a1023a5f9089c9b917f0ae5c77ecd9c7c6ff0c1c35115fdc8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6e89c343fbcbb855606bd20ee2b5061113dea2df95873859d8e600b0253ede53b521ae4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf8796638ee63d0b77bd99bd2798e84d8b573cef00265a5aafd69e3182b58ee5b796764a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2c6cc181eff28fe90b26f1c2cfcc5f1c499ad425777b6657a50b526338b2cfb3d4ab3d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117fb1bab1e25c395347cb16daef846e6526382614998faff6069b9e399fe88288fdf83c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d5ed6d202d24eb4f7e86484439ed037f4c8d177489eeb89f772832daaa099dd95fc4ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c9341f66ad89ef82b3120ceb0c343ae1c1ac6cf5b4f97e002455cdde95b3da81ecc0dc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124a9cd95140f799ec42a4612de83c87dd38dfcf805f25cb358011db676a21a58b48ebe3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0a87e427328fdea7acefb1b6c1a00b81eb4dbc6da747b5a801e6946dba81c0b94c9ae9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1994b2f821dc81e8c7aa0203f8da0b40b480b661e8874d2a1f57dfc52a1eb4344449b0733;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1badc6d1d603c63baa5c1b8ae843aa2df4ddf5bd3233b369860ff15626fb02f9269de6382;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10964baddbf889f9581bd8172e49902a4b6c696b9733594b41a8bc7b3c767380feb722584;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fa90511fe0f46259a19a3e488a9d4f15078a7d798a095b1d24cafa623d1fc10db0d74ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3a0d59afe4ddc422c5bdd338be28f647c7ce283c94f76fb64d118ef4d2bbaeb507234df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5fdc708ef99d0d8ae0b10e86a0f009d40e785b9da3622c4a03ab5f93be7e1128c97a337;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcba7a131476a3ba24b99af74a61e417324a845c8d6786ed31dab219c063591474e403008;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4a7fa43015fdc50bf77655d43708402e3176853ae4d271d7ef4a9a02cbd36bbc7c4232f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5d4201bad838c9a81b9e1ba4f716ee357c1d37743156f7c2631e78e4293fd80fd5cd5a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde256bc819be62b663b6066cddc547c4144ecddc35a0134d621de7866a89ba57d79100d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd92fc37e3f462ee51f0df7264893963c9f23c79231360cb0565fb495955418a6bcbdf3bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189f025394a9035c4b8f83d7aedfbe0157e48a75bf3b86c7ef1d5c24b27753764dbbdc94a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cc2797da71463571bd43918f23d00a30efa183b2737d81973e1c899a8bd91726e138693;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1debd189e5150a685647e2af7323f5565d92d85170bd97f3082d4ab1d51cff105b197fbb2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1192cc6be492e8ea09ab5ad9bd8694552f58d331ce2fac8bb21439c0abe7ba4d0bfb5c848;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1541eef0f4500e9f91b632bf9712295befc7433da97b8a5b2888c97b61f1021e6a6b39417;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e1c7e0934058e25acfaef337f9af1a82855ee90487a4161501cab5b4e413db7b386d517;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9aa10384789531472edfb96f79def7a33142289892011c1d62b0475282dbe31f696e284f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a36ace56147f79b29da1d7bb5b5498e1a76853ba4f0cda6e9f52e24860d0e08b0ba5810;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fa3505202f66f08aa963113f394c26c91465d5336561c7bd014949b4afc5260a86bf6cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb707fc053bf0c79d627acdba5b14ab9124baa25fdd5f98e229decf16bf16f759538a984;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10dad8e4653241018f8c03e7e60e4a2218418a156f8bb744673864ce4c18a5fdd5e3032ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef344e76f0a4833b3c29b163c39000405f83a53b2c26e10bd47e64e6ba065f947bb9bca7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6c93ec5d226720a7e9b01a342239ed549da39e1ccba5340add1062e202d409122bfb7f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ff021cc83288f7f6d6520d009b2fba5fe70d8a29b4a6eaa542a8f266fea03bad013b094;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2d25a838551dcabc920fbd6d050992ed9de7aa7325148ee343e9b9b37dea98e8ff5f04b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f32e765071526ad682bbbe9e90d15e3bf2fc78fd80e6e1555756737e6248135c86f2c29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175f955cbc5113f74637efcb16f131955280e22288d75f6f8c0de323ce484d8c19dd5b937;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdef873b60a4a7e798eb33d24683c9e84a2f69b0f6bd82a1aec379482e8c055b8dd6489a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ce40ac4528992344752f6a3621828dcbb6bb3916bc95499b5432e7bde20a3cfdc93f0cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61eb98adf5f744245e7a4a8261faea95ca79a47e6493cdbd969d4b19984c4b8ef0b7a163;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h767cd0aeee6b4b1f353d79f28d1677fb55167d625a8533faa9e919c1932a1becd6a577b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eba64fd3dc8e8d8f457bc5e46819adc1da02a6024ed67e0009c4a0cd247aef99364486ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2510047385a069fe3a2678959cd1b089fc262122db4ef786170d0da80ef7d48fd011869;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e7430226557c6f0c723a3af70a92b7324d4bef48501cd420ce3fba41b4be8b99bce6723;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7c8c9e5d17067d95a8c630335ba1719f65dfda6f57f3e8a0c5ca74fcde1d8c1b71d49db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac93416f208db1c223c8864ef9ecf3bffec989dcae469054e679b5464363ecf4fe25f22d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f1d9e1a730e638e1a04731428cf152496be91cc2030778757759082ae398d9216559c2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ad81b2b04adbe476789a23ffe90391a0915f3dd02d68eed8f383e77ed3d284042e30e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb5fcd31a0626616ed46320bf89daefdaaa40098ed3a1f9d2423ba11e5a10bf0459b1e7c;
        #1
        $finish();
    end
endmodule
