module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [28:0] src30;
    reg [27:0] src31;
    reg [26:0] src32;
    reg [25:0] src33;
    reg [24:0] src34;
    reg [23:0] src35;
    reg [22:0] src36;
    reg [21:0] src37;
    reg [20:0] src38;
    reg [19:0] src39;
    reg [18:0] src40;
    reg [17:0] src41;
    reg [16:0] src42;
    reg [15:0] src43;
    reg [14:0] src44;
    reg [13:0] src45;
    reg [12:0] src46;
    reg [11:0] src47;
    reg [10:0] src48;
    reg [9:0] src49;
    reg [8:0] src50;
    reg [7:0] src51;
    reg [6:0] src52;
    reg [5:0] src53;
    reg [4:0] src54;
    reg [3:0] src55;
    reg [2:0] src56;
    reg [1:0] src57;
    reg [0:0] src58;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [59:0] srcsum;
    wire [59:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3])<<55) + ((src56[0] + src56[1] + src56[2])<<56) + ((src57[0] + src57[1])<<57) + ((src58[0])<<58);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f437820fe2cea0215b3eff3b3f0309013b7dcf4dfb88e1f9439a29d6ee642e2234967488c1d7af0fee3c2ec06142c679a175c6f1b90f6a1a977ab1d24e56d508f8cb38857dcb558f5c73219f3c09c7a29d6c8c1fd0940242619fde91d37164a7058f9eeb367fe40a0911a5e0975c5a90;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51c59e05b3b48bef4e4e76a363e3d2d41cd7af85a99a378254a64bba49b5937aafddbcdfdd482047e148e27d0e37af4f3001c025a1cb72b83bcde22817e15c6f46d7ce7bb1360a12f2350f7f52ccd8a94015953a84d98de371bbfe29aba57e9398e387a8881890effe2db1dad0341bfba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23ce35952bac4518a143d671a33e424b118da5184f56016db995fa6e0474fd9f6a09c2c3873080dd0ac18ed33893433af2de451fa7e1760f2d2ed0fcf5a6bb362a12c28d7613b787991923dc4b015b5f5954e16c5543fd8a2a3f46f087452232b84d50a5a19d1681f9c55178ea097e176;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc435ba3b74697f1790ed21885788ac1215de17cdc54c96ff03150a8a9e87a6f40702498b68e6d6fe0468a43038b957c319561182c9f3ec0bac405b5282c97687e612c64f8316bef7885780939f0710763ec2555a3e641317ba5af76ca7c59d04faadc7813e7ea792c6d78271088ab4424;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8b9d991f2aaaf579e154780fe8381cf4251f72a91a99881671d756d432360b1264de87ef1f8c00cf32bfc2139404425a23bd22b094dc959f326de13481ab982290787c8643b697dd96188ec84d609675607dec1a841ece7447bc5bfd26ac022f4e46d5d583e9fda58dd947869f604333;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hace40c55d425380abfdf397a90e682a3e6077410aaa198aeddfda1935cd53454ecf08d09acbe67483eefa124fa37586746384274575b51cde51e6c34fef40ea678a85beec9aaef073972a39a6d2e116d0d41c4facb3da895003cd83e0a377e2fdb4595065fee5a15814bfffd24f34a97f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23c0ef3ac6417f5762b2549f06fe68f48ec746f9361a9b4b4ae73cb95092420801573bf042a766b4c05d1f8d28088dbde706413a2f9a68152cc75e7d3ef5a14885e53981a2efc9e97f5a428ed1230f1729efcd5c7fd06ed75197594b81355b3ae23307fd09b394f58a968d37b5b06fb30;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32bcd83c1582dc55db077a1e20cc213f0b2e8558c43a4d99044bc62a0472db5d37fcf7d50166383aa7904581911b513e065d9c7d208cfc3c3f5e43bf9f312495833c38108f5128cb6fe098ab2bc52e3631b2d428220d86f2007564af81266785bfddf1874569bff6bcbddf213a7dd5454;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79ab9ed8d8c0b925fccf31f8c66f227023adb84c8a5266e721d15d93a39ee339ff706985af396238b97d52668f3c1db45db119e3279c4707dd2a4ca4e1c12292ec4a13aaa754cbded40de8907952dfc2426e920266ee8fbf9bac9de8374c5c56d30b86fabd1e371d4c503513426126052;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea621c2e084c85c29ff4b1b735bf818a920f60a4c1c9310c10cf9da4c2731910ade64f28646650da35405bec1385d60b871a93a58edce5230629ea380ff2048f59097696a85c74ae6debcb124805b41f5a8b022794f615af7726674b2118437f0c77c7e26d8358fe83bd3740ff466e2bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b14c8523386e1c86d0aa2bc915da6ef975304ef87c9aec2de3db4507ce1f4602532b982476ad1d2dd8571649831dc18449a7e1a07e7b6c54ca7f7e7b53ca94bc00bf93141ce1ff2b870071c7aaad6208f05f6a2c2693707d3fbe3c59703acc3bfdc6682719f31333dfeec26bb34acce6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74b0b8337ee2111d27e021d2b0a1e150070e1ec637da7e151f6ad833619372b9334713a7c237a99833ca9c680be828fe3e8ae6610a526a118fe194740effebf620a86d010273ae69f8639facc04dc40cf454cbec8065274725b34aa0393fd78d4aa0283375a370abb9ad9ef70c0b30a1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haacde43162156ff8a0dc9fcfbbd586acf79845ae674ddcbcba418a0436c66670c531b2dc5e21e33d20f90fd9633cc6f9b5b70f5dbaacf50098e067a9bb01ea9cf5663e175d850b4c781e7a7f5bd59759a6b534cd623ac4b9045e158d9a3fc9229756c61404f6bdd3023b551cc832218b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h406b3a7468d1e8aa7ad151afd417f242ab23348c29da498861051cb4a5072718243361ba3f3252dde215a4750b0347c03195cfe19963bc1aeebe30dc84eb1207436778613e2e00161780c7db4e020381cb7f9e82eccafc5d02fc2349bccfbfab0753b78b325a2b3aba7d32f03c02c8067;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76dc1b84f5f42fc80bf3fbfbcf2dd1df34155875a03d4a7a7f49e440b75915acf99240d91c6485ea3298b7090d23177b89a0dd1e30435bc871311a85d9b6c7d0b139fbb930a1601d66de34f407f60ac2a76f116f3df93d7ab71345f377533ca2454d6397bb47ff51c0a4efb63dbbba52c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fd5687641f9f65fd6e4e01bfb7aa23f2e8063e1b8fdbfa17698652d7f85b109f431fb5957ab78efa49525073950ee90dda1c0ad221031f2887b6039e3eeb6adb7b727f7db695c450f5345765ae2592374fc868d975540e056cdfa392ea5a51204eed86dddc5f8598a9956f1ebe49f222;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb31782bab4a1fb0a7ce54fa7a36bfa57c47e843e61c8319933f3c0cebdf4a2b70c8612e8dacedc7e3867981b323420dcc46b43a2dc15239d2fb3a16ad2daa70fae5e6f7e5d859f47821ff8fb53cb148cb04ed71ce5436f180393e47dd6474951e3696645e10e95ef52686fc50bbe7eeea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf4afab8100270c1bdcae193d8e6175f04522a5dac5b4ad2bc51ebc0f69e0992e9b207f9e19a513787addedee48cb7a28ace0511acca70d40dfe3ef3c2f809931142daad5383994d5783feba0078e3cf67eca56cb79257315d45cd54c3e775058e6cebba9294dce27d82f736cad0b1279;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cb96051b4312b37aec114fa4732bdccca0b2b7ff84bbcfe1a95341a6e030faa818ed2d87dfaef44a729aea8eac43dbb9f3946a2622e404373ee934ba2bf4fa9406e8b46b242a306e02a34c1341803b5260521670de78bbb133025fddeabc7cb4b790c704a72aa4a2d6171c6aa6336035;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he266ba70eb78359d5f760d8695e00e623acd88d5e0ef27df10ac34d1aa85c3cb5239812677d1c2f1e8013e0e3ba01920f9ee3034b55a805c5ba1a2f022619e97fb7e32b4fc11514856fe39fc1e7e5104d1e60811621ebb99fa22fc05a6b2bb9ce363505d20efc388e911f37e9f583ced8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd7178c94cbedfca105d70fc7099f9e2f4aeee7578b37bb2b037cf6d490649021caf1db5e09bd497b1b397320eb87100b7d46d30ff6413a999fe7c5e1502535106c296ec920c902c9c74dc7f550da83cc5496914b34db9b0e2aaa6c5d6389ea559264b79b6734a6b2ceb018cd78d64b4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f5367f29026fbf44cb2351720c0afd3a562191e95d252010a3de5f8a95982ef6793db5301c5233ab54a2cf43ddbf972d0272ea3da47ea573c96cd829f4e49c18c2d817d5f90af729a09a1badf9f1c7efc5686eaaa2c5b937a25ee4717a8aac89740ccdad09e57c9ac1860f6f8587a2fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77fb84afb11958fa456d35316dca97abbb330f5ba9c6e1eb5ad1b192c3a395bd32240b24577a1672bc031979102d25dbabad92b1c83667bfbb2e29c53d4a474b1b11055161a0bd11455708cd0571a06f313d4f304b84741e0efca0101c18588e08416cfb3db6d907d3e760cdc3d36b66b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3518ebb0c109bf9f92f263c22fd0dd2f549c0172764a4ca2663da23dd10da5fac388a97ead2575c5ab3209dcf00e675cd8ef013b81c80ae97d74fe7eb8abba62d63ca564a38eb9f70c66f0936e9798f937cbd5d9aadbe8d4a43c9771befeef331cf69984c806981039f0b73409489cff1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e5145d1f4cde564d8398d3df063b1dcbc89ea8d58539b61cb5f89722ab11ddafe66f239ab83af986ee80d773a8fe94ca8a053968d692605bb7db207979e1e89cbc887996f609067833e7d39ef5af9201e086ada4f36d7e59a1bbc8856bd902d63a316e7520cc5716aa63a481d08365e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29b925324eaf17ab889d06b1292d5da7550e380e06a326088cac0c64df86f934821228ef780fe588aead42954a99eccabf33334442682a630d1da90a4b51366ec7a0dbebdeea8f9ff0e9d8040bfed43a51a77b1a0e381e3b0b554cd080e29e59a16ec4059062941e3879ae55e5cfd9c1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heaa04f8f8c49343ca63dba7d4d541b2f9c5374f7c96baf58ead8abc7b685b26e38168f0f2a25aec4ea7c8621bca8ecedd20497232b28e2a4b0363de294ecc310cc468b82618a2b1900e554f8760b722a2b1fbbe3f8f5923ba0e503865786b0b3b300effe7a6fd686429b16d1dbe732824;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h975336fdc8e73a26d65df7c7fb4ee254bb8db05d07291b49356e70b3a6fd6adf767675353ef0a7504918971d8a22f7e507f4aa0be0e0ad1fd6d9e0e648b042db46e52b537465b6aac34945d6ae5148a5829e4fe92fcce1da4768a496179d5dec1194c20a547b6f0229a7ee49b1a9e4ffb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had584463457a5f27ced2927fc29f3f9967cc7bc8ab087eb3587e9f11b834b384e82719d687699b69fad28b43a0e3d926641376db5de329902f780ed1bb9044fd90d40ea464e0f6ac6a5da2ec27d2b0cdba4a0a466aa020abfed34cebbfdab12e3c4f3f7a0e1d349588c2819a516f6b907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff30f266734cb8851cabd4387c06505ce1154ed78265a812e3c577b4368482e7dbb5eff92169610b5697e6284dea961116d563d6f5eaef4fda1ed9ec8a9fb7d4dac2a04441b6cddfe05f0c36285deb97bb7ce03259616e804b0d18943346d0cfaf79699ed1f32eb775c5835d60d2ae1c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e3013c11177e0595f55bf22e45811396b9bd767a3aae2311eece703cc8d8819bc3b8fdf9ee65198e04f3a32afee15b95f6b17ab877fc94eb05f23dd19a6e2368c062e118b8b6d804abcfb3bc6ff82f77265fc811d80d5ea056816642f1fd73e17f1e74beffb5242d89b86d5695283ae9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a5a168d513f2d49d69be4d393f996f653bbd9966cbb0bd2c95512a338d585e14ed9c28ab2141e449d33cdc3a4cff0068c84da47d225540e76b104e184600a4dfd32b1eedc98e3ec2216da94bd5e66e728451af1d4b26a1eae03c4078ce94e0f588ed12e9f09da1e88b692395b3e8f7ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78d381ded1780499956b6734845f546146fcd5a7f682af8c137b5dc1b8632c470c73184d0af36c16ed6935a5546d1061c2eb8f0136e1374fc690b2abd740150bff1f600ca82d483f74dda44673195ba33d12f98b6fc1dd5b4f1b8b9b86fc8ec064317e3425b8f67b2f1b465ddf3903e8d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1aee31dc1ad32e321c21e20aa85f127243c25c53a22205be2f08e40202a8f37f4646b6d751ff90c03e34b65d16dc24e427203325e05db3fef466752de55896fc0babbfc9e46e7c477497b2911c6b6a25eb315b2683721f5d30325ef59b15b8177626ffcf03b0a10ed885e6eb822e5651a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36cfd7f018ba4d82e16ff1371f8390392b8e6ab8f476ccfac8f93f28f9da5d84fb82c5155dbc87dcc2dd047d5078d3c1c82b7cafdae7cee2d1bf0c28d4c59f9012bcb272e545975cfb705bced86fb2429aa51d6bc69f344fdee2a436b7301d503139e268d3160deca03eed7f51b8773b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h902f24f09640c0adc3845394f1d9a4e3c7913c1b04eda7435a348b6a324d01caf1b1cdaa5619edc38c583efbcdb8f25e38f2ce35f19d6eca5ad7eb90a618c6602d3d744a6e3f8e9b66888f35e540126abc5342e88fc6e2cbb72f723778f39090be4f8b4ca0e0d31e3d416c5393b40c09d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92597f9f524a45ab3efb1babcd7c03037abc6a3eed237ccdf9cecef711447376d61ef80438201fbe836cfd7efeed0ccf851df5bd5caefcb1daf8646bba3f009c129631d22ca147e0e5dd1f21d14fa63c0a3f39e5da9dfd51f58233869f2409c83218763d3285f5e673f966e4273740f1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d450d2948b1977c837b3d6bb9a89b595e5e0b6b05cee3f2b0f989aea82127365224b3786e9ad3682f626e2783f190fc9cb24d4c399c41cb49bdd110ae20eb7f95d0210484b62b7954bcee60c8adc19fa8cb3f757bd6e6d1ad1ad9d4fcc8490a99be4b7119920c5fdfee17209ffff9d9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cb93161eefa2289edf5c38b8214f756a0e8a928b83a3b7dabb4f4560b612d1c12dc42c05b3d8d9411ec902d2602185198c698b40627c23677562e7fd906d20f36ea2820bc2cad6543c7e176252d3097211129ca549784a7be9ffa5ea95f170d9ad76101f6068e4720c901c5f27cc1f88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ff54d69fd21f7aa229049827843a0998a71a13297c9adc00f1a2576833af29784c80be823e102c15d2438334f1a4ceb174338b30c6646aede1660cb30d3e0e0c020830990940864202ebb6d28904cb0f2579c1bc77acfa0b874877bdf41df0cf82fa2fdc0318d167c83b7995eda45fd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1b54312af874e0ec8b92c3e9dcbd391300acf44df26d1eb677cdffe8289b180cec3a9e63289b42b8e31af270a5319f52eed124d206c49dd0100fb5eabbd10b184a0b5115f1870bfdc05018c4cb19cf2a96335ce4af6c291e10ff67b5c1975fbae31f025d0418c78e8ef63288ce93bf8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2627bd243201a877fb9e661ddb9e0f187858f68cd7815fc234d50a31bd2e66e5d1a8a539275bde2018bbeaba2881efd52793fbf871473b7d46ef9691128aba764f0ec23b76913e457b1406dfc9b97ad6dc05b0e80ae1f4b301a79832202b1aa25d07f1467828fd57fc614edcc841b8f62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23671ff007153df45a57f8e859330e83ffe051c99a9882f27730a8e390e067ce53d73de25c50ce7c41d03a8b6babbd4005c76bc527ef5b3d90cd1d974219c3dba1d772263aac6ba1f73000421670e71ebc66bd912203e7fe6d2732d7050a6a91dc49cf1cea566de0c7fa123b4176a9776;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haafb7bec91bf3679089c67afd70ad3fb22c928aa7074d36faa12dbb9e040a15cdd406209117b64267f175f6a4ac74e6171345e61928cda38e62178b06eeb52df211c6721fcf1fd81a0b4fef1d8ea1b35fb2cdcab0e3bfdc94ca068f810cd2755f88fbdf4e81c000d5c50e4d7d7403cbee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6de1640088d8ba9e9ae4b15bac98d530313d8fc5dac5ccad2d19edde96fbd491417715d1124f7907b572d39383a4fbf004930e03ab58a90782532e1fa5c6b8cecb8a387a98301f8c4757d2a60cc34ef7ac6ac3ff7d86edc8055479f7d888f0b4685235e8698a5e4455e30ed2e85b0cb91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcafd1a29601ce9aa23d02a22641af8c7675109b6ad95c311084c3e452354e25fae8c69a0659793f026f30119fb951c6562287d4577faaf027c76b8267af7abfa59f81ea29e97839e33b4b39c5a60438e79dc91edbb6f9806b65571bfe473cbd597e68634d105940256b53db1b012b5f82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2225c729e1d9d585a5be7d4e3961ad75067b1e757acbc0e4032b7bd3c0eb4b758cbe566156fd25fa0d7341dde491ee99e48cd6b152253d56dc63425ae7f1aa6a925c9f2d1ab99c321213dcb6c61963825f107b5586aba9cd12f9d01243a9b14db0e41f87a53f2e8ee456e8175f5a6c0df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdff03fd227c381fd770a46601b556e7c5337e0b61fe181c041001fa431c26b2ad6bbe847ea867401da5fde3f9adce1f780448b0808fef82f740929c59de9e0e062df0ed4c113f4e5e8e4258f0b0e2284ff8b290c46ba2492dbbdc5132cc4a7eced35d300d1e833dbdd012bcf6fccd786;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf294935c90ad73f51945a42c179cc1e06eb5e93199fba76645922cdc68cf133f9862786f70c11df1cff2e65d4296ee6b40bc1f355b3de2928709726d9066e2e67dc5cef5e126cc2f3783628420f7d112d212f54aec9bccd70af669461e52b375cbd33df3490f7005c95045b834da11201;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8ab2b4e9387ddd4aa4839a1f1b31aa7a7dc07f2ccd1ad0bd3643d68388e60efc13d07f678cd4e83e8c4dc3b9429ab9fb68a87d0dc916629a88785bfa0157db17a5d92c41d5d1bf65851f31e8837219ded47a732f3fa6f76c41ee76e49b052a551b06ae945e4dc9ecda2c5b4aa47e834;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6b08e8d385ef2377f3619660a2b57e87bbc4190e285e048384d28a189b0a4ecfb73060940cbbb266f32d8241bb587db981a86d19cd747cbd995d6bd517d9a4f76ecffa214234480effe227e6ad1c004e74f1348d57ec6a33fc78ee0d4d695ad486f917d08ae9de1a92931f1914073571;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32b4c2eeb58d69ce3b5767d45cdb96725e864a458d74825206be6fa6f6d73bae6ca57997c3802fbf487572a3449f4cd86d6cd3f2d0dcf270864175a5b3e9ed79a33adccce1802e4bd44fcfef9e110e130986167e49018b642a4d601c99ce48282d2a467975f6bab25901ab8935f0d68ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf46395dd042e6b7de79563322175b947e5cabe0427b890d2cad749f4596b60a30d80efa44deb880048d3fb6da3e6e029c5e8c30522e6a45b6b0227a0c3570de1d13dc8cfdf00770267a07f21af1e679db9c86ef4fc0175e80833daaa8370de772ef4b602907bb47329d950bef5164ffeb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17c0cd9886c98eb6ac72a8fdfd587fe2cb7205fd78b8fffc4e010412805e7021cc9c232885159a229a6512c0df6d6da805bce5696c38af580651d63ada5b92e24d98443bf88f450ecf2595c45069a7eb433e5f146c5674f8a2357737c4d3dd9f2e4e92bb28ba5c009a9e786d7652559ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31c90623ec58423823fdbf6def8ea9ef9f9efea99e04c9b0243e5dc90f5ee93ab8b290cb72a15aa9dd68eaf4a39984ff324c42a19ff1c7f8331b563fc6ecadcfe46429b51e6f117fb7f8491b8917d4291f5196fb2543ca60f56b05cc2eb112a3b418318c5eaccacdf4a347fdf0ff9c134;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb58d83a3e693ea2ab98af594150f162421668a3bc97ce69eb8509939a1cf17f4028e82df369e1ab258dec1a2c20c44ee49c563f617cde7fef7fb9636a1babf67cbb2d7cbb733ecf81d85cfd4e92731104b3b0508b8d0b4a75a86a14a8349daca7fe668bcf4e4361732a3f802cbddddda;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18c258c6090e7b08795847675d4a6a5ed031d77541d889e3fa0cba7786ae140a36355ef746525645db9c8909403f56caa0267e15572c88c5f96f31f92ca703a5aa1f7f014447a126747de200c7d00f188374da60dc823488d11feb4a1e99c24528a549122153bb48e865f6b7b2cb91c73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54b75b21a421de0f436208686e9a1fcdc47515b524f016f1fd620b157350369f3956332cd3143cb1ca2f5d038f5ddb65c8f7d9765a42bd81684ddff0933f54265a52116f41acb92218d9950309cc98118e1d276395986922c82c920fe5df975da994f5cb470d6dc94017b016c005beeaa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1444fe3df3fd5bed7cc47a54498423a902c2d119bdfc47fa6208613f34e6431225779bdad408cb8326e7ef1a67af8f0741a2ffcdd9ae93b97b0eb2982619dbb5ea61898f6266363f1ce918858484cc8378f4863ddbd7649e19c53f5ef701d1ab94057b2f723df1893eee5a9637343f95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5507719962a183330d9ce00ae7296f78c1b84804af4de4709c676430c62bce2f6a41f2a5c054faa2f1649416b4f2dfd03a41eb89fe5d3f03e2df9fe21b404e873b45d04a313aeb9705179a7434dbf332d1b50e4c9678e89a4ffd04c6451f8feb5dee6980d308d996409074a0b5f44473;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ab3eaa1bf021101ddcac57f2684debe26c365d8e56c8cfde58ed576b477dae181749b52d1136d3fe73bcbb74fbf85268eae830542f6f7b290a84ec5350391e169ccee85a14d7b35b993e9de29d270e4083f5775bd0119c8fd29ab3876730620bbc83a4ebd04e3a04ef7e405c7477d2d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4119d5c5d354307eb6a332b28a94030f4e87186ef396ff8ef263e904a0bc5e61d4154db0c9668715e26d7366f19b8ba52e523c4539400f052039ce744734d73115ccf6bd67199c65d5c2cc5aacfe68b7693ec9c1d17df6a8d30dfd970f0aeb2711983c95cf433fa54cf81606bcdb92c95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c62e2a3ef2194064b17300b09aa51950b825fafbd45f4bad8e846cbdeea3aad96ade57c5b6ba04ff75552f887baca4943e07d89fe9614090731bec784f96e4acfb6e281d931e816d542ba7389fa673641651be6e80b782ee7d6248a67708f52dfc9103891e6da5ffab43f18a8a5ff3de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b3494a3915c3b0c2c53b38650deda8fa65d8d2342ff1b6ccb3138b918f430987ce74b1c22774e4cf31c65cb3df8e1c5d8728f706221d68b6fe36a2300020e5c74cd15c67d654a30cdb07d4001642b38ca7dc0a241cf63a9a5fddb1a416b736e5ea5402bf05d9fa72a5f5e838c5dc807c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a5fa84afcdcce4bbc6c4de714ce6e75819fcbc34033e9e4a9a714689fd87ce4d2763d83705d48903f70e9471651f3a5d7e8be3b38cdf9ee4265cb9514fcc89e0567ab21a8417432fec51392d5e6198554f1be4f0fb0d0589685f1225c4fffd599d971b2470fa4ffde5f9d4e67bbe635e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96d8478768f168c7a86651afe09fa336cc838b9e4ec067c67d6c9de341ce9640865c96ae9ac795e7c313b57dd24fbe87c6b2cfed7a90a0e9bf9607dbfcabcc23bcb4ea8e7539c43cc5cfe5d331d035d96e21eb1b096e9dee1211d7c0c519cc20c2ad9d7d5f1f832722dddef0ed2180f97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8e0fa5302e735c2f83622057f2e841e69b431b0e862fb7c7f7b46cf78f33bb1f3797a1a15c285471898f48acfaf1dc5268d963598864e2547d21d06287a10a00442f470583f80ff87a31c11d94b1894e4ac4315eabacd5538358b1e578e33a036ffd2bf101c557c1f366dc4bf6bb1b5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h725f4c64feaf4a3315e2a46073bf5372bcdbfb1eef7072bcc952aab8dc7418704a97c7148bda3b6e9ff2104c4bd73a33669c75a807b00bedd20b1dbd68fadb932895a414140ceb3b13ff6e32ff06a2a8f0ac463a84771f56fa9fd3c2349dc7a9768f7c51c84506ee443375065e347d518;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9a511e7beda6f8c4c5a66dfdc4a58d728d176f2e7a7703eca840b0829678bf10fb3f86dcc2461dfea424fe0d3d47ad4272bbb24de61bf9df18ff2efbbd38de25ae0f4859693de33c1a66e76b5fd4a527c2fccc5bc5b6d969c27c439f2e67ceecffdb80782b8d588ba0312f8b771b0b02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0a56e3e55099c503cfff86583c1a6c1b5f28ab1e3d37cb7bd55391e16168f72fc3d0798abb740ed17d571100ab4f68f8b79139092f3d9ec164f98f1c65bee3f81e9678fb36f32c1205b8ee2dee4d7aa92c383e0cfac150e032060d702ec1059aaa1ccdd11c4d408bb0f557015e53896a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcae4482d170c10c0bc4d0270b4b669612d28c292849ca82ba5fbcba8adf94d7bd87d703f9c19ab8e90913ec0707a68bb35680db4c3fe83863ef201fa633e155f6329c7991f1fe46811652fa3823499047569a9c437fbaefb68c3a1cce0fb096103a7fb1df7ed29f0cdf6e3ee17f165034;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he55f23684d4b1a47ae22f21fddc2e5cfdaac390c0ebdf92c89d045fa190b914b504cbda1722a030ddaf087431e4d4838468bfc5d9769f8f255bce17a93162c2823efbba8bf9321084b3aa2ab3b9e6e3f56e73498178642f934f02d45747383bb2adb19b5542704fd7b2a272355568b21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ca61b3b564199c3a2a2f040b1e57adc9d0575642127b29152ce12c6d0b65ae76e02f750672e364f97fc42f6f370dfdafdebac15c3045ed996fce8b5527eee73765167c9f0efd506771d150d35ff7ff24625a6461d46605adda964d1b3fe9d33f847db34ddc1ad61d049f3a232ade5052;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52c00dda371dd204fdac20d48e7cdcf979b179977325306cc617534385fdc357afc9e54b073bf015875017f0b2727a45f3f161518dc31d21f493e3f144e5e4ba12c47a729a981ac750da4247c73de60095875f208dd9580a5c13dcb19731ad6db3ec04b87dd62b9e1700e64881a206832;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b3c0e6a6f3b26205f3729572998bcf04ed941b8909eb6acce62f34d09c93d182b7dc20af3f955852ad00036bc2ae0e18c31cc5fd1fed1fb9c4460eea7a60f2739d48b6ecff772398183b73e70c339fce9862e45d35a9ed16b78ce68b06a59a7bf9ccff5d57cba44ea5f90c2b2cd9eebe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee85f61567ff6bb07e303b5d86aef6ec21c5258464e771c0770b96ff58c0ca2485328d5783c79347c255e7fb65dda2dc598fabe3635d8be75e06951388750a0aa60357173715fd8e610c36a0b3bfbc39052da3a036f3feb03d1e5336df36ea65fad9abff5f5f5ea87b9e5d0e2d9ca6e23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11dd10420d0c0ca86753d2b01404e7dc8066b0283cd7ccf3da207d9954cc24247982ef08a37706883b92564c296a728e3c7b34bdbf6738bdd5cb08c44734892d1dd7be2d14f6ce9526ce7e35ffa57d550cd32ac03bfe8a9e32c98ae320337b70d67a50b140fd90b5fcbde51edd63b8f3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3a9629e89f083458060e322262ecff7fd55fef09584d088cb4f11d4a09cf43bc9626822f5558eca285a121c40fc37da9073cd8ee7d0108c7f02a349730ff53305b6c4d2e5c7c5b2c11e63aad1642a49c910f9b612e9a2f3e229628bc15fdf712910a8bc7049687d8861ce0287ed73283;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45a24948c10eb60423a06548ce094dd78936611203c0cab60d6f7495e33d053abc0fd9e1130f19e0803d13128718afb3ce8dd235c8cdb106310582ced546ef9c215c5f6968a6d5cd028230cb610cfb19a5a3b73b4dd4a8faa916d39e383e8cfa72fd405a6a3e61ce95d1fd2fd6983c1a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4467195b78e15c53811e94674b7c6b8da94b8a0051721c34359b56a482e4120434c1c4c77cfc994b32e5e6855bbd8418fcecf8d6c41286d70396ab8a33625c14925d34e56d16ae9e48f55fce0091d07ecebea08219b98941fc7848b2e52e1705fc0caed5f385dd33ff0a6613986fcf6ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb0b66b175583b8e9c61368d5d65d80d08c57e6953006482439c2ce74f1b43acc787c4e5f63e861100bce5eb4f4e5bee283d917df6d7a46a3b56e62bc1acbe6241ec5850178fd81a8a879ccfea2c9a2c71171b94d18913e4439e1e80bdf1a634a043fd2739662a7c7772d009fc3f94142;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90167a1dcda093f689217cb499241fbb24b91e0c2426ab5dd0cb7c9ac21be0c3541155de22bc8754dbb2c6cab584785808cc9f3b6d37b1da05a888bababb210ccdd5bd861ea4ea8ba31dac24d06dc66e092cde62247ba360c7773e0cf4e0fb94902e80d6491e087e2f8ce7efa316a9f53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd3f7d5820eea00cb4c613ade50df569527eac4c5f138d270f3715d2a84ca289ee42f343492cd640dad25ee4a07a013b69363dc5f1359e20e993eb4ed4820f7c2690acdf3ab64968490c740e34d15e5a89c595fd0be4a711fcbff92b7366b52248c4c78252bb940ac2b68163f14cc16d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3391146b5de6d1cf00f919dcffba5b81768b900c650a4ae1f8d4a8b9843632f1d614ee4385c0800081407d40faeb4fa8b12b4409abc6f2c651ac8105d2a32446dab43364ace3b20077d7a05404e19742d4cdf7fbf43e1584d7e773b14e112b6b0bcc0311f53f3d2c1073b7c0a46a9cda7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45d2000c32f9752a5dacee640561120174b39052bd8c3c99a58f75959eaec6d9539a0f8ccfe556311cd37b7dae6df000d2d5e50375916926be2d89e7ad6a42ea685bfb72469177756a140634dff7b1cda4193a95b45af216cb082abb435214c9838fba7050c4608ad9cc15c5d2eb6c2f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he74c8e0ffdc8c48a0182d04a5c39dbf69781722662c2962c90e1e829799de7a1e2cc01ede63529e89f257d38998c124394b50574625214ecf0616b0853008c768b9701b4170c8e99431f9eb79861c6f29166edd1c9f3354e6605f693be480f0d0454ddd2c34e0895a8b11d287082deaeb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3568fd40ffb6e2acc6c050bd8a98f5683fec1e8bb98104bd6be166a6f19b52bbec0fcd30ec06cbc2ddf0f0309ced9c535cb9fad37d0e028b95d27b91f105f1ac3bb7be0fe92fdef8c1b6c6bf2e4953b3b2bba6c5785ab578e2c540616dd1a49dcf8b146aeacdd4e9466f1f5d0dfc82bcc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e3dcd3168e58be6d24c271818c0c5076bb5f030bbe2ae9f957316475312a4e0c0a12123a568f47479ae30e52d423fc25e2583a27b4605b393e7986ad761519a9302f8b0c0506c7fe02a35cabfafbe51c4e70790cb24bc4420d309d23da3fe99043958419cd3baa9d656274a9b451bed6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2219d5d4dc814f1cfe31b7fddff1acdc9497670bfd15b9fabd9ccc9abca56365a9be78313ca48c5dbd7e54cb2d471886b9ec4261f7f5c723f455f3cdb99f6bd70e6065874e6674ff93286a6f68f8160784cdd6ec4400a015c36fdfa2a25a9bf622b29e1d6dae3c5cd6d2daaff3d3d9ce0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf937607c8a41fa72ba08d7ef9faae7cc145c25f9d090870de3fd5fd8940e92bc6c78390747ad78a7b53446d99b39e5be1948f1384f23143447ff005def0db7fd5df8403900ee0c9ea8ed2869812ffdaee8f617369a975dc3fbf6b6c2d40fa70ed205d2b4fa1371c2e2a419372c5dc087;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7fc17556899603c09dabf9010047c6ff83d94fb53f20086b965cbbb9e761804474fc772679b8113bc9246c2ee3c7a4e027d2961528e2ce3b421d1e8f4be3f9962ec1c6d267af80495a41983ba680830e3e0a99407077bd0d9e9728c1b7dfac5b4b84a5a95ed523bf8871aa5becdd8e54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a5d1c3bb1c9b4b3eeb1cba6eaa683353dccf9356e64bd50db077578b9bd06754751bae5f2e7a029ae6bae0c26ada2bb332bb2f9e9c2d11e49eaa9169af4ff5cc05ce09eebaa5c4b73ff331284c9c426d1a9ffbf6cfa26a9a22bb02b47bebd522b1498dac4b75350500dee86608fcc593;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb119ead1b0c141afb7ce1b67818bc03e821512ef9d16d308caf38a1e46f147175ea7be0a7e2bd96f8564a9ef123046e55c7090047ff39169442856a2a124dbb2756c8befcf30afba6a841f3982bf60829b689c8087d734e26ebf7ec8d4b6b4ab8d777e0829019d9955c2afe673815bde5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd46f28830b811da57f3acfbbe8f4af7e5bf6983421f1c1f9deca4d38a93ba63bbf36ab3fc2081cd2bc70424cec459637c884670c3c1753b80aa72ae203c243c7d72f969c06841aa516db9701f781d4b90b4484eb5d8c33f3b01dde00825b4647d1e6c85a38f40863905deb8530f2be5ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b541d8a0521a00fe338097e7ce54ddb737477064595a9ec6ac4e521c923dd4e28987f1e256946df0dd5150eca24dd65539fea0d155a20e810f2085485e890d0e76b97dca0f521ad340b8733c3bacf0701c27cf041297f98e3bbc81e0a22f9c7a4f1bcb77fe8c90510347f90008f2c41a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7749a71933950b0697820b64bdf87dfc11949a11e61243c9bf7f958912f095ffc34a2b7f19fd2feeb2e4c934a53476b308521b0cc518914c1864bfdd65b02afcf9ffd27c7809224f948067e3f7afe6ad347e3c8e5222d0e8d129105aa27f5779c3a291aa831a9866746025090e7c01b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc31872499b5c2e10dec5abd0e7d81a0925c052e279e72c89852ade9ec7e85f382fe2bd5c052ecb17fbe57ae1e697cdc5e8f2c73d427205eb7011602fa58ec75b20c0ee52ec5797357d14124a2b3852d83e7c58c8fd26ba982c6e85b3cdba748192b4c489e57ed9fb625cd10ee5b002021;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57e881eb6713546bbfe9b559686bb029000ef1621b30c1b92cbb38477ea954e385a6bf93e48870caa01914383e99ff091c61ccd5653ff4ab0149cfb40b7681e0fa03fe86957a35828ec5bc78ba2430803430808a007b6b73d3882faf62868981e1c79028e82cde4562b7217977156a2e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf0a95fe4abb457212c7be2d7acc98b9d229e0df004fa80164b01f1da54350c0041837aa4bd78cd79feb94c61ee30442d6eee11541ddf2b2b6dfeaba3d3267cd79eee73355f0ec4f383379d6333f92c8f95700e98101260e8b2a8f6907fa10f8d55b89d9b0eb3792f0fe75f962878c358;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h922ff44879656417c4951986a0e3e93244b3e5d3dcda80e04a4eb8d49278366712bb6a705a139ef88c480f19fa73b8f4e66ee3e7b214eb82adc78dc6babe142431adf1114b4aa674cde1d527b2f9f18ca9a64f3b3920a373a5c0b1d38c32d9312289c07ba27f074f4132867e9554470e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed177e80f7e112c327111535f882a4eb954ef212d5e3936a25b32c8e4c65d4cf5d6bdca0bbf817b0379f7685fafe51fca89bae25be28e693635e626cfecd414cb99b1f09a40cf4beec9a49142b4972333db4596aa1371f98d2893fdec5d065ca90108a349a92b53f6767f86d8d8b04d98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h558c776f3d632464eb77b59f9173445559a42a64a2932a002e58ddcb9d84a45b9e30c0182ce6076e8312613c334a3338423e4f9296f9d805d630d12397710d5f9ce5e7e54c58d1863c8840398dae3b9db1edebe973d5b17c97a4d127df8eb8c6fa9d6b408856a69770e904a1298b6da6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5e43a639bc282c60705b502d9615928894dd9f2a251c434402fc6fceef558cb76f1218a0cc2c3722d0c2d027ece8e5178b3d6eea6694a76e6f9fd36258c975acdfa935c7f1f27e673fd3d505b64d26dd52c6ff862d7133d4122c806c3a6ab41df381366691ea882875b3f646abf3292d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c4ea66e701c768a31360a7a2305b16f5ae8eeb97f1bdbf9fe3d02f3651afc3435c9027f0f862730b6638d680f46e664acec6599646bdd6c83da5acc590c268fff9a6c0a22fdd320097d78a06498b5de20c197347c1c3f639c792940373f0c5edd411f068e8e56f184db7da87c424aa72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89a9dce0d47f477c77137860424025772edec63b03ce13b252dbfe56eefc114bea53aed21f0da376176598d87a36d6b445dddedc75fc1b0cedbceb91bd74fc89ec30eca2befeb2d69b479a53a76e6ed6ee93b0b103a80c9260c71c8cd2a60f10c52f3707619f5acb353c90caf44c00821;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a3264a838e4ce85228b4e520aacf13d0b3099002c689650a1aa13a76d881637353ec7612b02518626e642eb8f848b488c2f44ee0308141d856521289ce280fb51f727dab2673300d4be1616e03d7c7ac23320be405fa0ebafb4d5d329884d9048c1650ea7ed84873cae26c1e4b64c27a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11e9fe3d706a6ab6e77313d2fcc04686d24f9acf268fde3265a7fbb0ba3c91dddcef60f192a150c896939acefaec0170b609267a4608f972d76d92565194531d0c69d7156b0a285ac01f580c1d498b18faa9dab8c7f3948dda0129250db819700163c1d03335dc2981228a63f1a55be9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe86828e095eec4477ae8eb48d7e0c968495a7a68efbd61e984a1b88b398263d9c8bbb4b9b1b25e40de8e66199f7c805b85b08673d8d5aa89694919b9e98c660e02cdd01f95b998a526367ca7f4f18cdb3fc8d49d560f321e7f4cd5235166d0a0131be31ead9dd01a0934ba5772513a99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h806459df0ed86392edb4b2d0738dfb84082dd7c672c3000ac3abbadf50a4c328dd5d5942a1d236d3ec06a7fa94e5bb96b656eb2a5505619ccebc1ad365ce16b3b47ebfae8233f2dfe9142f2cc9dced265ef99e06bddd53e058239b791dfa52946f085f22cf396ec03f64488c773f93a32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h128b177382bbe22445112406f32d8f9e92ce82362fbd3b01986694db9a831e52aef03c9ae979c6e1ced72eacbecf1fec6ee972334a78f46c1d02d6016decd6b656a714357e4327a387fb3392cebd8651699ce8274929ce8b2091c54b78ce01ee50457e233465298a9f06ca4af5043df9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55b49b9843980948c44a71311cbf2b979b79d790a467c32159e1d2dbe406c4537c8d491f48d8302eb6881a8403c491db7cd75cd22db0ef2ba12fd7f44ecd818446b74413b8e2f8ee2302a60ecd6c1518fc90544abf9a51e59acdee3e970e998a72eeb23522e8eaa80732a453e5c399fe6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97c167c1a5e1478554e46a5756c21c56acd01fc528e7366a4683817cfa8e1806b1eb6a590cc7306d67edea1bdf893765940d114a70bccd4be998f6af20867f9bffc7867e7317763dd890afe6ba230701e5784dbf2424c2ec69351bfdec07f6bc174b3ebe1dcd581c5659518f1ef8392f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b94c188d35b69a46036fda6eb7ef499f03785ad202a9b267bfe37a45ca175a9aaa9da0db35b0df340a4847125f77f9894185d9f274896cb1ff10ae09ecd8329508347260f7c76ccefb32db63d702cbe635ad48ce9daf1fc66e57117c4c9f32d920f87e959a488078cbca73af8151c1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha74bf5858ba14b801f6bcdeb76fb8523de1fb621b2bdeb023c32d45493c5b885963d0e6980aa1f771aae21fe31313aa3765204a1be267fb8a92102e08514c8019dfa5ab266eeb5cbfb82b2ea7ffeb46e09a097f95b79eea9d58670355a2b356def7499d2f7b42ed1c5854491f9c89fe80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e765d2b5680b73d35d8125aff977dd7281b0b22b632223c939ebda48d128559cd3d5b60b5de6846b2c8716db92c627da712719d1f0a8c5b7ee40fdb31788c8f89ab0520cd79143c70aa624bebaa82eedbf460a1a15bacc2e7e911d0649d6905c9d19416d4d0bafb1aed8399c3294f2c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4613157ec415111be8f279ae5cfa74624589089feb94ddd1e52904e20cab707d4da4f0841ccbc477434c95210194d9af90eb48e0629dbbb2fc334ee0beda4d6929a2a8c1b3f8d509f88c0e9eb60b5db64f0a572af405b2b8f2d49512f8e16caf1915fbf5fe9c1dfc9d1828551b2e99d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8ebbe60af2ef910afa5d6f308282da32e8728bb857891bacab79fd85cd79732d388cb04e6d8bf23d4cab8544a18191540d0c42837c6076094772c399d0b42128d3bf9e8dbd7cf2547b7c459b150a028010698b751541ce496cd4a7fc0919fdd4ca6c0807a4f70b34309196dc9f662568;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38fa3587eefe0b0953bf91e57de23030ed0a612d0cffb3c9df1b5d7f541fbe966c481e59084b406f135fb9aecef774df12b42d18571993f8d91f018ba3c493699669d2e101aabcd3797a26efff560bb16b2bebf34907ae3c9f1847d7672861df5851b23b2e53c9cf3f26202a47b6433a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe8636365b3ed048fdec1c171a19ff90d1214d97ee1ea2d68f3410a169a96a12818cb1086504f2599b9ad5d08fd4dbf51c33f82eb66f02276b179f0c4e2d435328fd83b2defacf6de10c07b7480108e02aa197e84abe40b7f6183cd3cd99685b6030c9424bb19b61569e228628fa372d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed913a869d023c858e579e6bcdde2555be45731c887c39ee6a313802b0e2be7cba640468e4b002bf231bc65cb9a0a724e624bf48073e42c418680830abd12b3f8619c7ae4709db6f301f1ff5e063728734dcb89cb6d4e5d07e1ffb0df37675b538a4b3b24f12533f216e5076dd3f893ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a34d0ac8e1e1e7bcce99150cabed51f13ef9fd720ac726db6571168fbba31e6694ab77e18cbcba284c84924740d410be201aec58bd50292dd5f0a571c9fb03e6004174b10e9c6f6da47eb020694cc38526244b6a0bfcdec3f31ae8b94c4b33669cadb2097e7eb090dceb8599af09f022;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0ee86321ef615773fbd3582999ea485128f7b2c6b642abd3530b471f719b1cbe2bc7ab9c63d64aa678d1945a8c20e2370a15c5c1d55773bdaa5e3cd761af5edc81ca3bdcfe8637bda54d9acc2782af5f1635fbdfdd464b97d983d6b5515717148c8227448e79498b6084398f07473e5f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dfdf6b1ce4cda261fa3bf8008fd0e199e0940d980b78be41ddd1c4e1dbda12331dd540d03f8e9c9640a0df23396983f14bff52a0400779b71f8d7214a74405449c24cf2ae68c6b3b571436122562c13388a9e69210dbee2f01d9d8f601977aadac4e186a305e3ea0eb3e977dfaad572e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha503d5b902e5e6d4b0f32c1b609c02ec983f891381373bb66f731ba91399b278a555f6c524ce7f041e2de6f5a1c94bbc70056c2c8f86205338233438df09a3ba0c34f6cbec136396ea2cfb499d224764309f9abfdb01db523e928bd11071ae55eff1e2cfaee9d8d90ccef705a4f1b6c5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba2f2755a5213a5cc736ad051a141cf0a68f794bef50430d8db052bc61be2287c44ef1ef8682f5960e69aa2965354b0ec9f9080fef24728dc879a6833f6d53dd50df0401f06a88786a8a50ea8ba99c8ebd1c93e3f35e0fa30f70565ab990f166b2885399280a13d4e2f3a4e8caf81ac5f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde45521d5b15a53e203d26f84ed71b455bc1e96f171063a120fec0569d5f50f83d8a5356a63a78192b2bc37c272f94c61e55ff3a9a8df50e8f0e333c8c5d44c345bd593bdde21138d2abfedd6bf2b6f49f294392be54246b02b0e2ef837ba0da6214c74960773a4824186ef6bd4c31b41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d45edd58470e5e2c58b50ead7c217f74b76144ba7245a4d0a1192478b5c30a17dc7789e856c749586223ea8b5405f164a561d9416e73efc379b41b5878faf797049f5054d2d52b52b5ff6e7597556f84f94c2adef00c7e67b8fa88c2bd219a88d76643a21d6b7ffdeb95ad6dd3d2afb6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78da20464b4aec1abe463254e872a874e65ef7677e9d36d0daca30a00cf72ef9662a6dcd33347c159afe12fc4ec0a743f470d524bc849f679751ab0f94429d6020536d87c86343a768d29513426e247ca68f69768ad5aa584f578fa494974c77876194c641b53425a5a6dd006c6f751f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h628934347bd6b02b45c39ff8bc213e5ed0d27ebc02c10f0ca98c3fc46e173a0525029bd74c73524072192e8fa11e6a83a5dbcc897f467ea8b9be5b67ba2f8d83afb130f72590df4104330b566a3e665db3a2a3070c55684e2c8afad252c66072e9a55503a9f3b13fa5e68fcb711090b8c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79458a379313d75148bad0bfa839e7b5177cd63028b582ac88d58d69a9a049a699142971883e1298ef96ccffe633657ba3d5e44a9c3fdee8ca1d9e8d88763dd8e897b3fbba21e9b6f1aeb95d610f3795c33073ebdb797b2cc9c2f519a184e0cef3b2e249f500fa8fd7f2f9f62b7d7cf62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha296a47626cbf046f155769f4a58d27199a50cd1426b2089ca56da7a81910fda776db44d37e32fd2b6c009753d67227f6f18caf6e45b689720993bc1bc602c7345ff47aa22286c6d1804c6479e577db1cc45c43fefb4ec543ef1f26a67d2ffa1b578aa7f6284d0aa667554e7912c4725f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21a8acdab88eb194ec9244ac6d83f5b610887943026c0438202fefaedf03983c3ed6c466c15a2c574a61e20181ba43d21461a9d4a571f099e3d5b9225cb83fb1cdf59585b66532bf7084860942006a2d6765783476a68a5ba1a0eaf4eb14b8f0f6c1d34e09220342824831407d096f405;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0e042da53c51303d73162a578e7a3fd9fc23670b45713379bc1a2f1e5bf3984556b8212b047997126d2043e7b1a24e31918b5ace74cc82911a88e27b9dd97d3d1dc945ebefbd7f8eb5a4d0ade3bd387983f147f99c43f6d506bd5667bec26898525efeb036c42ddd0ec26449f020409a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a86d92dd281990a9c6e96b89135adf5f3997168883ae5978115dd637e2b4fe51ed7e78f1f0dca2db651b550d580f7228ffde4fa3b469c26eb0b93077bc3722a795f58f89366645de762fd6d852bbf9ca3702165bd5c4d2c53c961757f2180501b5fcae8702c81d30c5364418e28dbae3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29195e90a89828d946b5fc6afbc2a1598be894f6f4f3f0df0fd61d6c4ba2ff1d14e3f50b0512fcef2e457e2f44dd8767f4a06500822e10f24cf2e150d4d7b500628d59c68cbdb0423a1f0cf7a049044e5295b05b199795ff4a7dabcf834822b575ca6b2fa01ed07db276944b684324a20;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc927bb174592a885440fb99a45f422fcd9267f62b5fcaa126d9c130da559d1b1ced3b4b7299a715331f99eefe0818f6167d378829e6fb75cdd3dc95b84d79544e6b36cc93b91d7237cb34b4c8afbebcdf4c98b4ffa5115d6273cd79709da78bde181e9ad4a73d1cf64f6102e4351dee39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd08c82be186eb1a4b7e6386ad48d2f9c5039df77b8e6836aa7dc825262adc75531547ee9330bf830762c3716b4aadb8db4aeeae8d7a02a889bc287a381d8407873789c0d8f71b0d4d09da55e6b384825fd2fb0c577640f06f44c7eb91dce4eda3697c62ec1e0dfbf09a7277b2defe95a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eb076ee8e753880d3fda27b7151ff60bf34291b40a42b8f885fb8e0fd2befb08329a4b7ebfd3a2a05bb309406f6b7e7953088a4c509ccb99915b05c6bb25f45cfb03d43d3aec16923d8fe2a56a3939d6eaeaf734d218995c5168b330bd3105a995fd29d52b8db937e9d595ec26114941;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef7f6b69f7f9a83efc83c388eddac3a4c963bb2fa5d4f3af95c90bd28bf4c8c7c365327623f3d9832e93dd833be3e8c17fcf031882b98139ffcf86553864c59feef6b8a137f8bbb1b6393e07bbf1fee4f73a82132b8b6c342c7b21cca01859c0dbf566d662b38cbb1c1703c190b296312;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha106b5b64d47399be6abf4c9b056a85097e254743561ad8f7021a64a1dc97973bdbdf4ab75781ea6b45313e4a0d596b3a03f3e81763eb1bce57f00caeccc24a86bcf3705207573af149fef3326f3656b35cfe6906c36ab852112db24827884ddd1d67265dddfe9c2e62a572b46851a3db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2a561d10c75964fc4136e013496f3737a27393d69a97ffc348d199ad8274c15480e98f124ac0fad63cb24298f9164f752c8b2eb72b30583c91aac05bfed7522016b0ca3a1580b80af9604bf19d7373f8f41b794fa7d3a18d9ed920fdc9ccfad7646e89a3b4855dfa8671a235b38ab6ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8db59f52d0ee52bfb1087f81a5f3b0070dd9abbc24c55f435e953c784b7c3f17d2909c9ff5d31560f4bcec7b7260620690dcb25eefec969a95aff762dcfa1165cf932c1d874da1233da22519303e390d973f1f678457821575a184927d597d1e7a63fe19daf7758d5465eac73098d61d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb9a2d9e03dc3e65513e671d6d0730fe388636650ac30e1909919a44464a9588e457145e05335e8e9aae8fcb121ad99552f0d4c8e64240d59219600b0331a495ced1359c153ea420140fc5dff594dcf88ff170aeb60039cd7941aee5a2387e917dafe0352a58025b00f0c4fb73345475d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h700fbce6584156f4a38066dec860290485e8e4480f0625b1f2aa08d40cb11ae71988e0de2a4152c9281c4708dbf25782f8a3679b1359fb8862a7f5611475d59a7c8ec83b179fdd324486b7a946acac4826ce95f361531a373e708df475d0ee4f8c41700afac6cfb14193be3d3e34f48fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85b24a12f1a3b3e4dc7361b95b59a5fb9201e6c0274e4994db12714e3af74d9430923e8cb0d6767b7f50548af7c8a2913af73ee3bf553b632a60f14c094992690cb48ea0e06b903a4b730a2b2104c10e64ef7db4223cc5928325c913d5950e2d60c236da5e4fa66a1457d54d4af3d0fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27db287eb63b781c8297efd8f7dc07869866a4b31d836d7b900ca871f208ef06d8063390f95912518bb9163dde270635b25705e5f4807001d161053a76f469883bb43f24f6f5e00bacfb8e49fe7e94adc37086d2f7ca69538b54af022aa2c36ff812f592e86f1a0cb6b06644b2f1a100a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdc370ed936afe669dc8cfe98226acffbc8b61ffac880bedcba3e03f724bf614b2e20b9a5c25c7d311c8488bf1b4165d75a98c14e699efb5d21a82fa1a2b82f34618915d19994e4f2fbc4e4fdd38653963590de96b1eddb6eb0fad45715661db2a47af2eb4986dfe86441c6771475f1b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd922da339a55b1530d393f4a03823f9a620ac6f3aa3074decae2c7fd16c48ce2103c07bacf113bab51500b55b287c1776f81b9634e4489e2c9646da81365fedde1ff1c5ff2e46b8d82bf7692876a6a00d710c3253e7ecfbff4a078a9e5b0d5503b373ab5dac22a9742f6d49af0a16c17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha012f7539ac57ca46ef6aa9e5c12475d41068482b2fe3c68d45885970dd4d255d523a7373bf531d4070591b6c86a47372234537e5fce6764e8f9244483985852b386be4a44d43ae8cff7f3c120cc5fa5f1fbbd57a82dfc3b1e8cba7481ca5746c24358a9caf5f041495fc67e52b9f6667;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd8f4a4f923eff40a9bba5732fee094d9606527c7035f6699b3a4b98be42f8c80ca24fa736f2a6e6c6409916bf52493eeb975a9acbc465e729fa9b91a3124180f3a331b9f18db721568dbef8146d2f65b7c09b4fdce58d2b80e80b468c82bb053d1786c4e718abdb26e6eccad4c1306ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42310e2424fe7e1d82311470087fa7eb773ffa7f766b65d71cb3b658d2f6e0586bc8d7d808278690c233de384bca571ae7057e6ff2d9104517541c84f60c404725b7ad0588c1fe270c16b8c4a246afd7c5ccac23d8368d3e6137057a641058a13054a5bb77d859d3857e6f7bc3efa88a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45ebbd470049a3628d05cd041af9ff24f10e833f5ba22e382285df9de86c6d916cb4ddf90311464912cfe125b90ac6b30e3ba228b9a4c2e21d0b337d54ad74822515404c4897e08a026c543eb544b7acf53e2d0ed9496e3287c57a0ae428d5258643ff478f5b5e63b5de4dda3d5d5b819;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c8d33ab4ea8be6eb79eb5eab7faaa01656c5d417433a7fe70147d0baf8f92f0f37bec1f06c785d74189b3c28d4d46cdd4c6bc694378d979860fa3ad4f1bad1502dfbcd300f4b074b100de8997d14dc5183c6c00d02acea119642a72b2bc2f2ed3c6f2e8d265cfc3cbcc94224e38391d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha650488df6b2056072ad8c2e0933dc75f5fa4825ed1e85f135ddf51862847f38f0a51c4ab2a261f16504c8b1dd0aa10ad7d4c7a9318c6b6c846da25c45f212ffff6055a089c1c0786e03a66c14b0fe431608acafcfbcf811596eb19a73218ab33433438382bf854b1f3ed9b14cffad82f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h634f364255fdd92f746d54368115bbc8b0d16ec0f420cdab749a3e117795f5b9f1dc33ede40aaa95cd0032cdad87bc9969809156664c8f530a2c6380bcc24b6df3c37b5352a5a20c8e3fa56f794da0f3cf1e8ae1beb122e9cfa55cf7c98e37ee99478e8667bfada94ec651ef032f92390;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9495eb7649fd330949eebda06d2c169fb9c7dd8b780075986179b258c0995b61823fed71949ed19c675653e09710bce859f1b0c388907f6d0eb2cca2d155c0d61f0116b329518c8d395b541293cc617461adb51b63171f0a63a100ea259062a0722afdc5d3da9fcff21753208552a440;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h952c09026740ed37cc57264542f529376f59a55aac2368449759d789ed2359d93a026f9217c2a4ccee7f4976662d2e33e9226c2d2e1678280803ee60c9cd5054d5ce095797d5b0dcd0e5b03b9d7eaf0a8c34f1907c0f3c1b9e3efd1ae9b5c9c051cbfcd7a3575afac41ce4dada1c24c8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9b7df4a006b9a38250d8afa772d4ce27e3a852e08ace806457e8fd10639f9094d4e1dd5252f33ad49c1df13bfc8d2ef1acf99fe64a53991d0a4c52e059cb9e75c9feed68ec75b3857b3f8c35039b0cfd973b3b33919875796e907e3fb1719bcfd84c1c34e890334c68a1281a57d12569;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h237c483aca5455f3fd5500fedbd6664fc80d2ae6b69ffbb527f4755618281c9f91f75a48306b0c8a9d1d924d3ca34a33dbec67817ddaeb9a0fe9c46487c86c8a8e24166e18ab6ca47e2336a1715836fd7882dd8101e7bcf893be1e4d545bc35b48c826766f40c5f5d05801347990f756f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h605df15ed73a07120dcdb1028cc592f6102598427ba7df31bff0784cfaa97fdc491a980af0a622a2cafda383371f5bc3a667be645407b1234e6ce8a72803d125856716e8809163c5dba458b61e168c87268bc99426fbb18ac238e143fd10f36fa3427ce941b9357e0b959a2436c8849d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d6b3c5f966da9b08c40be1b169dca5d88e347c83aaeee48abdf49a38baf978f530f60f18ebf42d5fb0eca8c91fb19fcd798832e2c23be2f8ef776b75e01aaf1c53015f157b3d18f53a1e01daddc6f86c0abf79e41757a62f33cdf1f8c66cf049993e2b3ebfc764be6c80097290de75de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d52c1e738c0f375f7bcb9ca8a6c2c7be5c77cc12e594d98e901419d8bbe941145d0f9a9be8f55916dc14456eb81038101af7670d21a31ff38e54250fc6d50081dadd3978a1a1d21bd53e6f929c6cb5c43a0b097f8c46cefbce088a87337c10b4c8103278c7cb8d53cb5fb876969b342a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbaef9dcfc41e2f6c83b02529e8cdcd76a703e609a3d1fcfe450737a4b0ac731736bf669c5b8fa26aac6fd29c9a7a42885d5f629f2edcaadfcdd0b002138d9c0561e4332668270e6c6fc809d0e8878e21b7d85cd001569bc98837fff348fddadf85f0a4fb3529203d7cb5f2fb6b98608d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1241a11e018e32ab29837652afb2c24b232e1b93fdb0417360827932d6b3c4b399eaf2e3b5bde659532361cb772051400a4d5e38d9d9be340db816edd39adf2576895f0b7e6891ea5e7e55343a51ba4e765cb77d9db53608da6d44857e0074afc49e8e0035f180169d073780ee0065bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8ea90a06181faf6a03a216ef1134550bc156b85bdd16d55b3fc0df6347bde4b023244516013319486c50479015c823bb8f82fe1a9b80f3488896e7716439cb378f889b70a1dcaf8df5b2074a8f3d73541fdb486171f13ad88e2ae9347272c7662d2d957ceafee08b51dc878b5a8970ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf64aa2306a6d7b59cef22f6b115a3c76259e65e0de78266b7b12fc8d8e44cec663164d2f2a5ce8ed8af0e305abd898e696a3b0c0b49cfa94464e0cf3be8caed4f9e0f190f8487bf5cc11285c2299aa626db43124beaa3549393ada90a69306e762e303d7fe40fc36bd77c62ad9c00bc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e86a60f780d777a703a16f3593ce8af8946de74f0679d2a72a96ccee28827ce28fc022a7b54fba50c9f0a3fcee77a246a02399cbd534e106785253a44c3e6806c0186b3f77f0c940531efbd5faab62e403de2133515ae5a33b80812df4f27edbdef5f8df2381b589cc23bf16fcf3224b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc725f92dc39982d56459ec9579a289324e072779eef17ab42d85b220766093e1c4d19ca1c7d50982497406d0fdbfbdada7e831e36165b9a299b170a283a61725580c2df833b1bbe9d56e7635b01c31c7304be00522ca051ca064d05e0b06c0ca5d591e9145d1e3b2cb0a9c568ceba6f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5aa08d5c9d2f76a0fda3902acf815d02a01fa87a348ced74427e34246b6dac5827245552878edba7c196356912506f91db85b479446623a01712abc4370a813ea381e4fff1a61659d6e1d6976873e359bd2a5b66f4e755197bcc8cd22a964e825f37650503f62d6e3e5173bde9cba5d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa64eb4bb7987a1a2721ac1d4aeca875217994fb765ddecb77136bad5df5a154f4beab9e6981d9fd343996388f7d9b7058b2e1e449a00b1af4541b006f71373607fd58178079cd109be55f4d0dd13ecad5fb40d44d06dd1a2cdb23500332bcffc0eafe4a1ed3c624b42c453e0db1d949d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb74783f07a2a4abb3c768bbe1e5156707d52c89a063e6c36a56176d47d4c3bf133d2a0c0b42c94ef9677c01bd2dd647481649823bee1b794234fe83ecd5503037870b55a36e863f8f7ac93fb903589301a8669a1509966710d6c7c7bd7325554a196f31d9d19286b842ff1244bb1acd6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d3e18c342139e93663c9a24333e16369b1c656018641f8b374f940d43812e09d00e13f457b2439092f8840d8aa8a13e6464a9f13d6d8b40abbcd733bc18d9ba24baa3f0bb2b2ad72818a7469eead8efa20a8de5d897ea70ee7da557f8c3c03025a6203cebcf1d6fb5d649e9afa2f0787;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf8184c92ed712043df6d36c9a71e60d3264fbde2b5638af7d0851b2f1a1b0877122f13b07435f00b2715e812c29b98f2865ce828a30b8f6620bea59d5c30e927475fec04c74a80c4c41a47c6e3d512dc4f15ad951c0767055914af004e84398afbd34adc901326e6938c83a1abd13e5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb782761f9208dcb839d74cc5c8f103d2eb3ddb34e618629267581d14afe8e62f369d34f388eda17ad5f3781a9bc4a8ed0eebfdc4ce4af101aeddd72a8bf9da838462e471f7cad4a3d4455cf784d62151a31299cac53f68a7da99ff7e207ce751bc93e7274d66ca26f2ccbfa6f58ef77f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f3c40a33cb85a2b462000673dd3b406fd5cf179684ac0d8be0160c40f2304e026ceaa74518fdd7d62ed1b77c1a971e34a0fd56efcf36b1df46bf27bc466722e2f1c5c6bc3d2e7cd250c40a3d08019c3b09116f5fd0dc1da4b02bd7a56f8872f7b8e894b00212e9004de369009f0f242d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f2ffc243754a280061f1ad92571da2a1945e39d6630b83ee538d1af175091b969614fa63b38b541a2f0bfebf804d1ca4094c36bf8efc12092a60a589d19a329ba281331f78ef8f607005781ed9158e8a7f04d3f752f6d6efa2a13677e061d7ecadfde88bf3c2a95a47f60ac35c57628d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84d50c48e4cecd1f5f412919f7ec8a4d0da7800db6effa7f1e968c18ffc9accbf06d9c8ab7c3c8eccae4676cdbdb3f48364e7dd35a77d9dd9d038be088c8ca330cf6957e876a3586cc1c14f2521191884687a97d382bcc624618480548bcef1584048cefb8716137d029cea9184e3294b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d3342b4f784a78fff8ae336388e1a83750c2b28299b65b5558811182e5d415e7dfce2fe91b7476965d89fbd6ab886a4a3e90198a83eb2bab1df74c6554e60b3351e9c7e8781ee95005768b6da489d1ae829bb9899c5ded27745c0f46a9768967b80cc891b323b227654ba9153a73a366;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h426b3b88bae4992ff6703f8418314c30d5c26031a75ec185c4ddeb908f0f2e03871e6947796f3f303868281faea5fdda23d0ba0b4d1ba9accf72f9cf4d33c3df059bef0f473b123c94da91e134ce08035c30cc2f1f629b230c13a21d7cd37ae708afa3d40d0079f89b5dd39d4bea21349;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h611f8b0351369e8e42505f80b2e763737f0b78eaad07d7f853b20ef5f82512c24eb0758e66ac1538ef10690be7678fbfc293518d493698d7686158a06bbadaa0c393fba621c17a8cda9f05be6d8c2211b1aba64cdcf44ca209126f195dc341eb6fa3c161d121cd5c89e8d96db108cb88c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c6b8e36a1feb883201dba48f165eb4b3fb07d02a62a2a30414589c033445a1c459043618f5f5c7b371283bcc46edc192b2f182c0bd1f1054a61bd2abca7f7d3cb60de67c1ebaae00de2e95ee3a8b5e6f1018dc649ea5528a7cfad4cf2fd0aef896975a81ac547cb81cd841b2dd7f0dfa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2ec9ef0275647834d7e575e6a734e9fc190589b1badbc6e2e7f4246f0e18df1beee4e4c9dc9825a8d1dcff29e1b43622428de1729411ca83b6066fae3f3481f326243ec4239c8f030bf739278f57752a44542339dfa92604f670bd55e14fcb0f1e74c9741adf7fb6c2f43cc367716350;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4337b4840b73377a8d283bee0635cc335996f67b800572f795fc9d937639ba795345d7cd03343cafeb179d14a9ec7f70d0898d1f29637a5be436a627fa6f0bde3c5cbd79b408ac56efaf23e7916a369d68763ee9534ff6a431a9f0d12d69d78e6d9e744f11ca52fcf9cc9d5da55fda455;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3245df0dad58ee2ef7149649b450441a45274db8c1c64d2d1429a560aa3e1ffa465e62b32b6b38eefa47ff77fa1d50ceb8a1d6e6a009154b78344eade4b916566c0c31211ae2ace5a3bd3a57608f3786f59b70769ec5362cae8040897aaa520bb875e9d5a8ab8d6d9fd7d19a474c2bc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf1d41c52896ff7651b031fcdcfb4bae3f0ec7390612c46e95afc96b439c416ce64e667b132b407f63bc8b9e289e25aef31f16be4b790fbb5157b62589600cdf9e6504f85256df6e2c9de8f6f27923038a7758ba65a3baeb5e342c595d0ea3423ea7e2fddd52103516daae1119f6f117f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3980fe91434e8d0cd36126aaaf9f181ad61931da1063553cfc070e638a2f9feceedbe33b73360c6bf6d29ac71231376b52c88836200d8a7886ce6c699cee45b40c81271721ad7b55e269d2e174e43a93c1a9e1c1ff78ac4072683c2f0a155bfdd042e1620132b38737010788f1e2c35f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h228ec2b721bcbbf8b0667e2a081cfa60f349752a678635909c14e7cdc5fafafb3251fa739702a0fa749839cefc2397fe9371c77f43d9085019d2b216281859b1235b96ce3237a4d2101d2a3e40b29fe2fb7aa45200fa401c5b384496977631a8078d78d20fe2a4c68a475cd0dbc9ddec6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0afdeb801ff20207e73e56caaeb242e73ca93663a1d9876efda82fd51814a9324dc914d0ad7b5c36e16edc3a8fddf0f6b5acf7f13a7dbbdbc90d172e6c28cddb48ebe713e90861fb6ceea4413eb1412c8d085de5ff134326c2ccf9cd00fc04f43de4a0a02d2c14ecd684b7a7ac1f6358;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he80a280005f835e3aac15b16d29a3ecd81646589afc5afcf538a48f35bacfc5bc628c976760b973ec41243de5d2a50c00fdd3baf772c579951c4e3e4ca424817435d52505aba9cab67f9ecc87e85e7773f49c1af925f357c7b4b4ef185402fc9f64c438cc9dc9fea792aefdeeeb1ff1cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h945b46b879dd9d14a3d4d77ebe27828015d31163d107ed3c181cd8c410af5a8f8c2beba9666612c2e1c9e14434f44b2c93e37a6d413215086917d0c57ad3ae37c4132dcd4bb8a318b0a99b153e67b0b9d5534d0172826102623a69c579e48c564bb16018aa46a23eb910b6ac1ac690938;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcb42da1382f650be2cf3f32e929d34a50797d6e189f82e790d4088965da31704f986871847d7f7c7ea1ffab028fb3ffa67a7454f4fe89723b6d3503d0566f79a939652d087f1a039ccb5cfbcc2fb5e8fb9717e6a49dbe8d6ded90a0acd86907aea7a5e48f58b03ac6d9534871c54e5d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d44a0e1dfce1cf8e5c42f8601f9972ee049085e5f810a66bf22224098aeac69b0024bfcd20c9917eb124488319cafd2243e2aae2450b2b2e0047018d9007c06b01fab48613eed6ed19c66f88beb9f1052242a7e70274541b99f31c92150feb495a1e037da079de228e779f49f332d448;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29971fbd043eb6918c45a0973fb4a2c85243ca7549ed75888ffc6d31ef47a74390013da36efbfb2a4452aab606677f3a0d6adf412344d6fd25fbe62d7097ca83cea38635c63a79d0303bea5f3139e10c05384722ac122ee1a7f9a5cc32e56e49f4c91619e871fbd93fc15a4e0a062238e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53fe302cb946330d3c1c1bdaedb9c1783e2c71326377e4fc60782b9804debd5bb8e80a47ff8de04b0657b40fcd262e65c2fe7d80bee5fe2fea0f99796481a93c9cbc2501d552aa860de2ae9d2226bee40c9410d2b03e7d444da49894f24048a6ea96d6e28c2dd9ebb60ae6d2ca57288d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b395438ad882f110be1e652657cdc68945f1a408f939dd5673325b0eb92bce9f7fdf522101e72c242dc294930173fcb016a1c733bea97ad25df4cbc4036de79a4a5fbe7431caf088d0acf1771b5e8d98ad47e9e87d5fc63220f548a7198258e5832fb5b009b96bd8f0c7de8fda7a7e2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h837647dbdaa54bb446161bba6e43b89d26becfff573344e2c3b2713823da110c5f3049362bd718fd18a783599ab3158482cd9aeea04220c9e94985dc0da4ddd5e53264f0e14e3ce6aafdaeff6c29b69c6a4e228603dd75246ff0724c1c7025b9cc7599dab897e62106b60de3c6549a5a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cf1910adbf435e0ceed56936383fccaeeaf3c3951189ee6719ba8382a0ffe31e1b1459f5b06c97ff1c306e78947f6742483a7c7bbff2f8a49314b24b1ff6d9ef681feb15dfceb6ba932782b6fdb7dd7bdb4ba86a35fb949d004b228ba04860080163e0e59c116eb6fc5321752d72f272;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h651810d400c8719da5a9112911d5627fd4e2745194778b03d13b0079395002e0ff08872d5ba98f4697ea4889ab48d99a46bd0de3a782bdebd04dd0405d90bedc07c58873dc0368f6e9a9558769a2942d4d0843367f940c9f4a22918d67c5357d53713750dbe5bacf39499760348599ce4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e38f9a1e4406451c381a14d4a32aa24f130533a4edefd3542fea2f10447ddd4f59dcfc3231787ec600cde087ed50efcc97008596741fc13e79c1d2504fa4eceec6bfb8f67d36400ada7468929bdac00759d036fdbd03a424e324d956bb5bf47c54eadee3a3daf981a1002f56e33d698c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd36d610ca1e68badc4452a2af0399295801e2f3bc301de3cb93e57b276df1185c5e003bff000b24cadf474e1963ab8ee87a3c2b416cfb6fb53eab7031a0bd961aee9eedc3c0907548c5905c77ef8957d56e201e0f82704e7203201888adbe836ec80652d599f1373165c4894533699be2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h612d7700ce7e5cd9bde4c6bbeda2db851fbfa7dfa276a4585bde860cd195fd3f7b1706143f0d6bc758d05fad5cdd32c63b24d952c0f8e77c45d2412a896384e364a69c567d9c2aac80fb78b20026695ca99adf02b5ea26e6303e9fd5e3eab2c08ac5335038eeaf060f88692b9d853d107;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5dffbd0de8085b1075480ac919a4d2bc2c780d2fa77b30e04dc0bb0132bb6d1e93b811a5378e108f626983db7f00082dd5456e326875cbc07026115ee4ed7e027be3e83c9b4571152f42d753d34a7a299703335042934734ce56e1f0e05e05f578aa96c2488f13de8098c1e25911193cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc767c3388f9290588a461487297a8cd6b352c47002bab2659b1441bacd7712d27fc30ac76e285be7abf2fef1d2f2d1d7a4f4ed5c7c16d55d705222be79354ad6fd4c302fbbbee9d2d0c169e88046259ff01876ef281ee6a7113a63e30a8d27f06730c768e4e35e60e1245698735552870;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61c6e3b6cd67a94f522067732e47a15c3134b8dbc4c858471c1e03d9e6c81a7c756d8a1e582666ca6df5114507c8008e7993f4a614953ec0c364dd00a8ac63910965031a9c9facc902cb260fe389a6e2ffdfb507129b54b6f4eb382de87d4af2739d67b07bb5e9c85258b65a9a3b9e9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc48ab26460a6478ed5c6d9253771595e2bc2ced9fc809bf83b270818faad4a498dcf8e52bae8d3b6d5e4291b027158aaab5ea0a0fd9ad6a52ed34d04b8168435e0cc8449a6732eafbd5660ef0fa1fd285aaa717ffe8b245f5baca3145336fff5427e07555056867d5c26cbc290b0d7030;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35b45009933aaa51fbbbee6b242fde8bbe6bcbb680c29274ac62a5397db7d202623c33f1abf32ed073c63405ae94f16c75df856e618829aede67d7110d88a37e743c13ec55750fd4ec91e3cfe343677759f9fb21b07829b730b8c67046873cda3033a2b5818c7705e56ef110c2dfb28df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h473453043ee67a7ade869e8ed63ad38d0fc57c31f9a0341e3290f0f9b92d3f4399b21681c2442dd9788812c6e308ad477cf8bbda7c5bf08c9101700072f53dfff0c898521baa38fe1675cf9af6908ccdd529acec5b0ba7d6059b6946c9974801158684aa526fe3a5a35a0b748967c0d1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfeba410a25885ae16ba7114f3bbc07d44a082e1ed23c3b61ea4380b762db6ecc743eed477eada08720af1aafbf3a09d438c84dbb355ca89fab5e5a0511eb249681ba9967043e64785e1cc0997b6b1609e88a38d05f4dd4dd75fb5b95e5b85cf0c84e9cd1462ebb87edbba712be2b0d67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673fbf70ede9a7816f06a88514cd849ab9a821837d45bd14b923d8d14e08a0e64948fa69f5f739a03761b2bc4b6338cb151e487e74cc98351669d16dbc9c1cc334179d8c3ac7e6da28b822122a27c2308580e6e89fb2cc1ed4cf38b0dff9cd3028ea7b9e60ab2e21fb7b530f6839a821f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde99a12a5a97f0740bdd02b5c50c1e0d25b9e9ed58259cc2550e8fbd6673d36948cdd1f866e05d363270db6f4ce01c69280c69070d65e1cf754151bfd92bdcc9deb150f143c435ab0a9f7e11ab6ca895e519d0c6031f3e07c6c51e8cc03b6a3ccc9ac9ba89229428c24e100ec474a1da4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e28e0f2492a104d24d70c88eed3aa6f5774e6ece52ab82493138553723d493f938621b2c4da7ffff08e054f7940735a2e41eaf81a96069a43884835466432129d0c8cc89089ec9fe5b7b3a53cf59c01ff19e213d46b2a195376da8003f1e4658d3ec706bc026ef2435b3ff33fc6a20d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2907f92638880f05b9ed001fe99831cc0f95479f555503ff3891d81b0eecbeff10a9b25386a48583fb30adfd6851e89540e04d2fca18997e2777780eb92e374a7456e724b7bc5dfaade5fb4622650e83a9b844baa51713b2c22c79f206a0e1301be0d539f3033d6a84ce06b21ba94b1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h328ca7444311d0dea12f90b5385f6b2e1dfac38405b923fbc052e4a9f1143c8a5881d4bc1d73efaaef3d4611743fdaf8242fa9961036333be14bbd0db83daf16f9c721e53fbab3a4f646255f4c06a1c49db4491e5a971af6d6b10b3a28b34fcb2e597d8ea5878bb25746401d9446bdf17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3101810e924d06aac6a5dd9a46482230cd1c9a4e3492073f5b3a07240a68a8902542a2da0c8fd352f7e6e87271aab417f16ab74895f13f458860d2e27f653d40dbed0e6ceb403163fe8f54abd933cdb65c267bc206ef4745eff66c6a796b6598acce20334319c03b5a1f30ad8179dc79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1936d5661410573ee1033d552de6dbd222c33095446c4315e887bc12b4ef14271655a3df20f87e796df0dc1cde9b0d2d6d0b0ecb6e50e7ac5d767abde9bff752885317c819823b4552857d3983758bb955bf5de2ace7ec5335544a5cde1d56fc0f4404296e6e607fbc861c66e27f013c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1058832fcabff4cf8996e18e75708cb89c36bb06147caa9afbc8dd0dab448de072eca56f5f63fe933ac67a87f3bca3a42f73720722e3fb67ed3cdb997991cbd96527865cd44c66e5dda0be2b4b74f8ff1023f0adc8694513ded060cc7d4c8253d820318cbaa72e9b0e0dc97cafdf3543a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98a708bff505760d39aa18a6e1020bfe9b40e9129847f3efc23a7e863dcb5bc704770f918916019bb8d1aa09d5228a1b57bfba3c731072819d5b86e4237da5977e520b9431f3ade2cba62682d58a2fdb19579dd3be6b22c00a6ceb7f7c887290fe236b9fef870792cf510f8ec70eaafa4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5197ae0bd267a7b82ce7722b0a20cb46dbebce38b8694f40be0c4bee679572abcd10b5f3b5a02cd60ebd571b4863d0fd23107d18c871b420eae5447a39628f3d795ca080d3dbed3a9a0185d8482ca8617de0947c596bed907039dc910f7863120ac3103969d8c2d37e737a7acc5a72da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b94e3604a921526494eeee21abb69acc054ceec20846a8c3ff915b77387be8bfa2593237011fd3079771619c897fdf9960b01d2854b81533e4992f2571eff96f58f79d52ca3bf0a39fd288b47a8926604114b6f96b3abc41deab0084d74185ba54d08e77cf94aeec06ec4c613c164540;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b14ae9dcf7713aa9d6816983e424c38e48140fd34c42254171f42596e79473ebcbcfd64b8a55d3918f489920fe757329aca7470efa6c5e0c8047d8de9922dae35b4b236ba374a04753d7c3a28c88cf0991c2abdef62bd8f6fba7c55960a084cae9ea06d09dd5782268d5cb9b09e126e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1282901afd1b7e88db21cedd4abbcd1bb6ec165d2095d16359ba491db12d6ccd58b97edb6cfb77f1f9d4e66cbf923f977cc3e1ecb33b0cb64ab96ee6a436ed16e811a282540cf77d3b8537b1dd80c59ebaf455e9d4dd23643c064bc7efa86981839dee4dfa2cd2f9adcd04be62f9d94aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4a8c4d7379630830247249d9fbbe1d5796340d35fa9b18e1f66ace5cde462d99a78c2b4c4ecfbe42b0ab1b707a22d16a2682795afa606c86a1a41d582306e04affbaf742ecfb27e03a40228e1308354e41f5c92a19c5d42cfabad4e1bae0dd90de408c3ee20166733fa9a30b0d1325d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf691790886a04019c7fa6ea6677e2798c7902b75a23b0707025e8b59542ee9f0a5e64c0495552daecc016af4130c1220488037ae5406d79ee03794dc5a7e2fd5c76cec2cc780b76a5df537ea29ee6d13e11d62df0e7f37d3e602317e25c35f762d2ff65d6aa121ef2c57f22d12cd925b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20d8ccb0136222ebbc7a749b26033fe4e3f1ec688a8bfcbfab3f45b00526f7aad9ea471fa1a17eca69a632e9ddf3a4804e833890521d7adfb617b594f49f893a9936acd6bb0a6dd5fb0bc05729b957888e82cac8db4b1c04b7f951cb2db6118fe86ca3a1df47718c8bb53caf166117e9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e402afa3e9a12b9befd9b625eb688fb97585caea0f98fed162d1e265359a5a313af1438f8c585739adfa571edf08d338aa41cee16fe0b9ae89903d75f7c5ec80625ba3d6034768b0d1d71dcdc797db7912cca372a70bbca8589e7f0d662aeb3de9f1a879cf00214d8fe9dc0019403321;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd78a32c5dc3a0e7bd1134736494eae1701312e645706d59a321d1ac39d4609058b6dd2056685706a42e0d12cd2e9af3587677f28bf00787bb54974122f65ff6a49b4350dfd9ad5b615b1dec0849ebfa86d72802735ec3f250755db2ca46bf648184b3b8879a7dc8e09774cd37775643fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc99a73f20557833a7dbd64446e250e298f6854db4998312b610be28da9aa3bf3616d4e4944d6284042803dfc841d8a42c05103b3fabf34e0fe16d86be43e722f3b6cf5ccea728cca809d813bc2d1ed11d0cf944de1b132c120ef0bc6210f5b4d0ccee73d13cf14c34d480450b7f2376b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16be846cda4915c901055a8c82a84bc1e7020842dcbe8031c0dc45730f656b6cc104d2aed9ec7407a7a85739d90fee5161a1379b642946d04313bbd61858945bfde7a905975e067fe35e421cf7c05064efa4c8718e15a5e439ad0b7dea1732625ae0ee43f753e9042b3f30e0ab52dd93b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f105b07bb0b881f1b275823323a0bc5e09ca2307d2668079a5cdbfe3d2398c2a77aab846df0e382d22aa2f1daaede2667ec983635d3e101bc04ca28c8c6c3f891f3ddf6d6decbfbd748840780899bf37698814087322e594e9852c20e65824c353455b6170484c5c7a72bbb94991ca79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee172d4d1e0dd487966fe8f7b13632cb62b96a79aa759a59bbb5abf0ad5cba7288aee9673b223fa57d53997ddc166da390dbfe5ce3d97b6154f0e5285e5f15b8b6c4e6eb5e76890d3e257abb2c85928c87072b3241584867fe1139ec7bf436cb028709eef102702b63e429cb216c89f01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaa42a2004d9ff63f6b43a06a82aea52e7efd7387cd3f5d01a90a2a230e0c13db7e2a807a9f82770715984b664049a25eb32d9e45e11df94d5dc484fc551d8585ad1cafe241c0d50c8d1c240833282053cba7573857ef1832fd75796503d1ac5c7aa04d94eff3fb54ede8f43a08c72899;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34cbe1c3251db175bbd091588890732896a0fdc48a28d4403970d09881994def2c3bf657dfa18aaf6f4f59b19bde38417144b21057911a5e98a402c0638fa210c1d7661ba52ce861fd0a08f73f35323d2ebbc0b56d9c5aa7bffe4435f9258a82a98e499dfdffb4907ba042b0311371d0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cd12c9719d7363fddd6d3b5cf7440afb338905a104554ee4c3e39b28c709902c0582c6d30fd3753f6eb5d12b4acc1ef744104f4cfbb98db39d594307592822cda44c54269aa4d42e23c9ff5e8c2c6354854f2d8b59d2fa7aadabe10c7bb82c9b6de45c256ac4fe03925a752db043480f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcef5757f893f0083d08ad6d8bf338a6184bb5c66c17b48a8f56d3ea4f21f5d5105c31a81b59177e541a760ac9221182096f4d51ed04ebfb3f878e077c7c65e445f52653a161abeae6a7a703fd8c627285e6938a899938b94a240ad3fb596d516f81d24d3f0c1678b1cd296aa053f7d12b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f6d45c15ca4143b7a19b823f5815f6355e21affb824c6dec274cb715894141cf70144995a4851c2f199d824e3810ac48064231c65c983d279f12c97f8e9e40d9839684b17205ca24db58662a3d3d7e792cea9a17f51cf385fd4c774f8f401edcdbc5ab7fa77a550dd6a596c28c9d85cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5a468c1489ab5babb18d13d72669dbf2c03b48c5145966091234ab1abe367e08315746c0103fdbddc0d66a5a0629486ea40972640ea4b3bb76ffe6cbf1b5a73734feca3b4a2588f3055a738254fd94e47eee70d3dff78b7bc6d8d5225f8def678d3653d70e98e058d963dd3e812d100d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha14b61ba86c7fa2e7c2a2cd53af21be90a19041a44d9699238262456419ffb7e9a626114df677271378c82d094703dc36e2158eec3cc7a604cbb7186d7e7e036b444f1061c1b80fb5c6dc1fc78a192957135aced612891ded00adeaf0d496a75137c322ed112d4ef8ba0aa3d4b8206443;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a0ba1235c2746ccedece08db5face6cf0688365996e8572945f076ecd2959b2adba363acef84ef5fae6a98238a8668c6a8b70d6fd64049753d83053d362791d48594770be8361dd695899f25881877d080a493882b28d93c5d17c1a6a4e1d0a87b90768224028327358a6dd9bdbc2e79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5236ed1de483e2dd61ce6c72d7995a872f986446288c74d0888e1af61c51787d957aa106acb9a176b99d35463d8e7fcc70201473879f379a6a17fec0eb8944ea43510117d7aefe6cdba3bbca75d72da5e1d54af86aa157451692c158e1d096ab2820d473471b685ffbec188af3ff98c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddda3e82199759cf37e6a5f8052bce194c5a8f686ef93e224ee1864d606ff2ae0ab18c5cb10f546e047d3ff2ca613842cc439b738976075014ab9257894e2610509a3b370dcf3fb37a7b50d6fff8b3e1d49762c86b67f1103ca2605b6073b45daded5c2cb618a07ebb480595f0fe21233;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0755968093a09262b0e4cea5db73d409dc114227422cf4d3d2ae4f5995c6f460b2091047a9607d80d7b2801e7067bca6e143a6dcfe1743f7424368be69a2cb1fd3f2964de649b335b2ec3d73c65cc86f2f4309ddc940c2db9a3cbd96ed2d9a0cbd382ca01b60ba22f9bd94a78be743d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fb947dc43154c3367662a7a89b538b50571dc401d2d2191776efbdb4bfce4432088f64fb8d8a785e6bc11404093b7dc23260a90623c77f15a9da767c8526311c941586f0f2c04c36806787d5ea7c6027a54cce0bc27dc2e4b886b9b29674477ecb5cf0817bc6ffbaaf73b0d75d06101;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2730ad4369c1ef63082dd09b2703cb53c8718b925b8d51e23475d395e181be10ea807b68b0552e74c00451bd60a1ec03784ffca817fde20ce7017194bcb23322fc3f9f28c3f63e6d5cd245efd1ff34482f09955ff61a454170dd7c2151e69b9fcaa8069e318e43a81a2c363041080025c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb52aef2b12de31ae858dd13c22d3c5cef1fb96be84b475338308876ed919a6eb50d5db777e821eff821a0b7e9950d8f4588156d9794eab48d362831cd3b225ff6355c7bd8985cf1bca55447c30cdd0d7274aea95bdee6854714e08c00dcc4005887da816eb2614d3fd13568ef666375fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37caecb8f8fc4485cd47176574404da90278d969974985ddbd09068082a6c953b9e7271e3398a7dc0001b9088e1998074dde33862cab162c56f211a72d1204aa253c52f5a60e819660eea66e1072bd6f1e69bfae1d5285e24f14d5f0c8a31e8b4e8dded0958f52e61f08a44f49aef6c81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h354bb92f2155659222bc0c2c734625cd6d6ba29bbc6f35274066f43be46c18e1746308684e77c224a667275cfe441138fd3ab8ea00a739606236c9a79d410f6d6458ad8690655337ff070d5ad74e1fa6cd5b8b3ce9c1ac3f19fa9b02e404ac5751f3e044f0f6dbc4cb6103d0c8ad082b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d740d847a9767adae4ad35b5ac93cf4a7405389b78728b3526d9749697aa41a876042657bcd2adae69034694b72de16238418490b28e197bfffdba5559439a7568569b8580c32b71f6486e377c27b0f654b591171c0beb805e35b78c61a6663ea9e847dd5a50723ee63e72f2ec4b7cec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha581a162459423b9392648ff0728074374499ba98cbafbb7b42fbae3d1d6204d78f55ddaca0d56d94cc3dca9d99cbd7cd53515fef2dd01e5d5b32dcd2c40772160377133e148c0ff14ee8d09b9c71c2abdfddb926ee93427c3a21c6c3ee95cd9063f08085c6f06778fc85337924a410ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha91b4461395eafb1597f6545bf2c2e8ee2a76a5a41013e6ff23f47c6d39caf6e092a347ec7e5f27ab94ae4345c0ff36205fe79b48090fa386695314648a08d101cafda150e8e48771f271895668585fbddc4bb2633c96bee864f6a714af48e54e6a0c8fafa7915c2ab0d143380720a98a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha21012f8a62ddd15c4ceda862aa54f1a00b7fb3ec037fcbb19b443f86081f733b638c7e070656b17aa286c89f9fe371d72598534299a9dbbac21643c6627c535accaffe8ce0f3c052b00de2c65ec352ea4597ee6563516c8143c2ace7cf427be94174bee8e3ab8ef0df66c7cc3ae85bd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48932759be797d367f21c2d0a7d21ee79d5b08ec784452cef6c0456e6e88e33265739b7b14353414056ff8e8d17952b1397f086c6b9abfc69a9e850c648626afe5e055fd4175162cc3928cf0558d8f23af808a87f98289c85b21d856b5b67205b4e1a766e39ba367bd2ae1c3ba0c42c5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h724643923d05273cb9d1877053d2b4f980366f8e317cd7ddd4d70c706cd8a7f8ffe7a548503426ba769e21a224c27923e6f669b182eb4fdfc822e6dbd23d3de822b8e4b545f07eb62f3145fa6e3a2c33a1c1fa7902a8f9739a9b0d4f6e105ceb3f8f416daf7e4826a3181822d3e98ceca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8828b39b910b4d6bbcb6318cb16c8cd558d1a212fb2d65459f69583a3df30528f6454fcb9467947b8752a1691d4ca59a9d6f13672b4c634cf943d068b6f55267e0954f94e1e69399720c22473354b0293e37d8a83e226cceecc4f6795ba2ceeb761339b90e6feabe8acae83327bb7b62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59e47cbc1f2bfbb296c79b411221bdff71ec6500a6fe78bd6a6553a3040750544ece13b16900672acc2294ebfe0260910bb4d86e67902a36845b1cb48d7758b6de03817b5e911eecb2f07ccf3aef9619056f1a5e666371943b440dd7b85ac18630e36a7b33f8d5c44a4eebc77e11dfdd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b1e39afa7961470b8cd0aeed983f268c7a1d8079882f369e7b6fa8a8bcf20afcc6df9caf52ae38174841c42c89848ec7621a4fe909bdd69c46b701522c951eacabda98631ef95acda82b742a8a89cd91891a4ba777cc4d437e826b80cb59cfa7a590b0af66a9a9b6fa5b62af7612c731;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8df74bcdb93d77aae74ef88a8f9ba75f2544a9fc10f578b134a9862f2f79d4c0d9a8b418126878739f8ce834f631e722f2f32b42e46940bb8295880cbc934ffa9250a6a1ca595be34e553fb9d8f256a45fb30861329267618ea2868d6f3dce0d5f4d2f4b0bac9c28ac8f866faca5d12dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34bcee65e3299e8ddce142d850b635ea43b5a8231a52dac79a89cec85139bb2f77d5bd27a496783acd3ae981538df240dcd0b468c3f12709ebb69a98179c991d3a6b4753fcaecae4da3c52e24d068e94e518815675ec895c4961dc0c944424fba73d10cea829419bec97978d9cb7545eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8065b3cba4696c4096586db618cfaa8edd848269ef0488e718894f396dbe62a13ea6fdd1fad263e44260ffa494152c7588e56f9e2129d61b6df92cdfe3dc2746fe89c40dc7df9fa502a7742a39f806d92b045674625da35b8b4bfdd9699cf67c59ce6a1256c8ac63f03c4bb242182e38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda113d0d7eaccff0dc77bc189bfdb13b7678e8c44a692b093eabe24adf4cc34bb7fc36365cea40e07ca13c5b092d314f64e7b2b3d2aa85aa8b4ebcc18a1acc1469099455d3b4d2a791616c32b61ff2f26ba3f2cf65e1c2428324b0a9239e73d5aa2c3e7fe63a3e6c266cb424a512c72bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93d6133dc6a1728044bbf51c28b8b21d791c2e3ed15e221d492b6ab7c6607a00a8b9f522a029c89e401e397ffb12230c8d1ecabc5969a5dc455157cb7cfc48ef8136dee7a6402e3ae585f708c1f2b73e3c9e507134e3719c3ace9429a3e48e84f64a485dc9aacbe36f2db2e3ea9856dca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97d8568b75b42d91a3aca376d97932676982d02416099a78c7f22328d78888f47ac2d29a0eb2c5b8f81880c7703d1cc9a9e2a8ce3d81a2c71738a02d8f1c117cf560d313fca45b9ab4261ad0666e82a71df06eadd011982d3369cded3f383b219c12d193c85ec703e86603987f49164d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cc3cc2d773dd571ef6542d6414fbaf511b2c2059027176d5ff2aaac73333f2783f21de0cf229a0cbcb98ae9c72bf4f90458d95856044a8080094f23f0a277e210e55ca1b836152926a7a4123631de2c7cd894b117059d4acb57c5071083f44c2d5dce1c9ee9a429d905f20546e84cc94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfaeacc510148c55536a0138e33877c37dbfd980c2d48cc776410fcf0ba895e740e685239213ea159febcba3c3733e5624486b6fafd0d4e99c45e6b916d82a2acd6cfc12b86fe50e903d83bf17e3a3770cbfc93d9a658e156f7a551e47265ea1f31796df098a3b17e4d3dde12a4548067;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43979575d65c2f2f0dc1ed07c39971534e261ed0699e318c096a6e911e824b10751d9ca47270afe0b30997be63988037925ce5308e91534a5e3397e286d4a0c8d4d1089a94fd7e4371fd050652cc65a55c3da15e23dd9b4810ba2ec67e546b45a3b66c86cf3d01b4af588217fa662610;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eb8bfef49b61d41bf9bfad822544857da7c43e71db42cd860580d670f4a9b50922da5060d0dc35ffa34efba60805aaa6d45cc12325541f463db7c305f7b41a396a94003492ff21b54fd5a7aa7d6c05704a7014659e50b18b68fcbe723d60f3670b39263e7a01af67f140f7876183a42a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha54bb72c74e2f953229a5ef79c17b8f4c5133d3828264337dbb9e92ba13fb0989710ed519de97681643c2ef01ce8448a06b827d533e5dec995bbb05e2eaa1ae65e7d2dda851c00bbfe07f28887a0334b17e36caee38016e306ddadada31e399c920570bef41082170dea5d91a1d66cbb8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5289bdb4c7c3df24ed569e5b8683863fa45e31dee1a5139e10b478eb4931fa1427a752c21db5e76c595bf18fea4ba4c588e09ba2e601a7f1857feb27733fb97f10125c01d65825487007d09ba9f8b48ca97395480d16ccc43617c72db1db619121a6f27cab15e816af806a022844c0ae4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55dfebb80944cdcd29d00a54cfac92475482d0335e7f2f961c67e9cafe75b0569dc4c64268fd2e5cf2a294b0cf840c9f3922852c2e6b05392543b1aaa8ba9a78b766edb208daa3d039fe04b53c357784d04afb1a7701320c581491f6727c21c167a09a309d6a2701d10f0ce64a2ae7e54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc6e35b005485c04f0cb9602a011bba7c72db220eca8a09aa04f5db9930487f8dae8da71b0f7c1bceea1dac91dcc9bdffed863ee8e4a9d84de0ec74eabb1ea40355fe922be3a265bea67b3dd0e4204ca1f912910d5cd06fc0d6a29ad9e7bc693a08d97ed06796b3ce65d101213d6648d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcec452eebfcf9d3cdb5eccdbc52d701d473fa3707602bfaf99673c0669b0f514eb72b9e02aa7abf67311dfabe8c47c702fa61dfc3cf7938bfbc921f80c45b741f62cde241417626ba348eba659a4c19f1587bdb6c081460f4c7416dc267b0de0b63d138ee95af5b62031b88b9beaab08;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0ef5d58c150afdc59153cefda9ec89b3ce8aab8159bbf546b4c8a4d7f4bd8bca50a62a60d4c7e396822fad3faa463e67568a0dd2c0341adee3191511cf2bd0291d83c399c02c20649fd4d4e42f7b5f8dbe6af216208b6a30d4827f3e0989a0634c1967ecd8c3e181ab2abb9ec1a02146;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h463da510c1d171d2f07dd95a43ac03b41d71d56a46a4db35cac725c46f138e826e986deab8b48f901574773285ef95855690af787959538eefc69e95ce9a5e59f91b15152aca3ae6a789971a7d7e101f4891e1ea455daca2df73bc07968fa28c65c492d51f4ffa6af74d7bb284bfd13f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b5a9c5bf39dd19886f95c1754fa617062e467aa8ae60dd4cb42606a0dc3090026368965a6d032b8d484bc061ab0aa98499b0a975c46599566c2322cc0101fc5df26a2f57c6472987bd66f7ade50f86557e56ae071cbc469a11f410676705a4a90b14430da5b5d96e53fb424a25945102;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40360f1319648c1362db7ae0fbf401ec9ba69783599e76f6f8c4511270ba3e570f4c00b71cd9933ff4ca1f6d8d6ec7fb93e475208d18a64cda6e6de6e9621fdc58738a5a3d4246a33bf558363359790ca865b2293a826ae4438f58de8a13e62ae1f2bb19e5c5c9c8a4f1a9a5e63d330c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10d1d5265d431811b7c33e8039d17311a4e859d26a7bca336c1749ba290d731e0bb6b5763a80347418e4d1004accbecd3414edaadf303ee2a21dba68d76eea3ad678f107f6a41fae7ea1c12d76ceb4c2a8c5e91e13ab3dbf17b330e7af76656a2843b294f912118190171fc34c7b3478d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf986d819644c22fb6da1585f0ef758a719b91ebccab74a3c6ce2797a1a5b84ac2b9fcbb90f771661fb1f951e8f98b527fe2ca93e8f671fbfa9625aaebf147126eab214ab1a251374f9301c4811bf1a81b43aa93edde7a4487d96a01d8d863b7d8c651fc144201c58563ebd89121f560a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe9987944f5161bda7d86eb6782348ebabbcde0f43e6a60f3296635e6914f72e2ea8090be0e68c868e564270cf800e3fc6d2e837e048f415a7939420fe31752fa8b390ad014d48df381bd45aa93cb62e5477dda17af77c0acbf0ad37cafc114436d253ffe0660c8ee04556bdd0d06eb0c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd470d69d80040877f8f981f48e03b30e542da1497dea7dad83f8e35d20bf43582ecbec3092ff6ee70ad68322256c06743cfb923f3796185be7c0b4dffe7fe5bb9273e0c69ad4474b9515efde237ba42a801a9cbc413e53d0ffc49a4868e614f3233eb422cb4b8937df83c108120e3b9f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd365f4cb811ad0826537bd6bb272febbd1e674ef6c58f354474608500ad0f87255e3b26423195f1915c65d68c8e90e7c19691415de2c177b6af7d143bce3b059daa013a417553e3625f29def5d71ea6fbca706ae695fc8807fd4289f26b50dda537eab358b98119b38ebdcd69e3d46f8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h577abb8bd47e602aa46465e7662efa44872ddb038d5ca416755b65dbb52119c25930dbb3a582c616358f9d74e42403d6958fffd89a615d5227f1048553f2064d3b2f9c8b2b7fea36e5112df18cc616c9a54f62178db8720a5c70fc3625c8118269d38b5225eef47885a0945df0eaee6ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4d028a6495d2c09e86ce452448904c950a445c6f03ead5b7ce880e3a6ac078641f25cff512710252e7056dadde359d04a4ddaf60e598bb1e178132eb893df66d64d4c41df4175a664bfc36ef55677ce571383b6824740597a6a19ec8c32b20d6b8085b88a7f7c803556b0bf1acf734e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde32c1f6937cc4cb8955aedf02a35dd7af4e17e4c796aef10ee84ab39f8464656726e358933845dc72822bbfc8f387fa584c78ba2dd2e951b399db8359bfd2d8cf3894b18093680fa2a5495404fd11b248a17d0356e02cb221b7afb19fa7942377f0bd0331df0daedd92c4b3be94b2eee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23045c0b25446ea0014f2fb029c1ec45353aa3730d2b92b53a2cafa624d0836970d9b9aab05286bb52cd741357b2800594706b03a166f0885ceb67c6349b02f50076684040c040207f5070cd28861305f636870f22042d6ab6c345c3808811ee73d71f8067c45069de0ffc084e9590072;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2418aa18b4c43df2734c6d72f47f0f55f7c5c785f22d725e74149cf83d7b5e075b9808799a779b6b2cf2fc9e9c8641e75ead9707dd39e99229fe857c7b724178361d440cf3f92ce6b0cdbaab4c931b3df5e4e7979e834d6c71432d5f3369dc44888a6790e0fcb87763a0717348e8ec31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0509684c4fdc9ea22e3bf6ec6d7d486ed73e76535265b0d202c32b65ad6f5556f77c62c9fef3dc5759a05852dea40d5ae903a914e1587d9bb45732e64c3af74414caf342a8da6c4ccb0e6c5afecbc2c3a31134eef115da53961a5f36be42d934135db7a5f88e092858bb3f08a7f42bb1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aa2394bf82679bec971bdaa399b2f449201695f0d9d5a9e3001c77afd82533497714d1a4d63f05345c45d7649830c4b2d29b5a33dacbff72feaea97b16ce313e916552f22dc46af600a980410fca23bd550c9f539501809ea734e5d9bd62cf64fb89e56c6c3574f972a32f6d299a124b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7b25ec689522de3cdc7df9671a6eeb0198e2ca7a30089d576f7d148c0c1d6e79c9cf33710d329c7f40f19e5399053138a725d144bbd0afe0bcebebc825c6a46a50fab869759272cebf8a97baf11e7516128c4ee5e8c7e3972fdd9bdd2ed35109f39459da5b8c9364c4ec547080d3b032;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26d14c0970cb81bb994ec0866304e52b28fdd9b96f4f3780d22d19ff4662e38c17951bb2f6f8fb28bcb64e3e39dfa87184c48449ad5986f724d3118d44cb8778e1350fb8069b291f6c70a542291abf77149e5e0f8ca53ab39e6324a59a3eecd09e2c9f8be56edd2330f91814e869f2864;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62487b5e7a5373118878ebb89182ad40e9c02ffceda881d880ebb70242a6ce2e056042598f36e012c309a9172ae1f0ff44911e1d7ab466d6b85a31976a168feada5fd29fb30b4a8aeb33020fd41aa25c9d7c75b434793d6cc5b7d36da5d3de90c2b361173cdab7ffcb6963b430c4401a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1a5ff56ab2eafd4ab7be1b028c9fe39f95ebbd73e96e69cea8717568c85ccb5fc9ed4b95836bb6806bc0d0200901877d48bf3a3b19fd5fb993f6911b4f2f30c9dbb4a1b435b070be3483546e7f48f03e119bf57f49bfb7f7c074c667839583d789bd064cda05bae08dee0ff6338dffb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f53908fc1a4da89421ce3801fb182249575b4109c9663982e6e2a14ae9955ed5859b2227781315a72c34719fae10f4a1dc56360a68327f1898e20b54bca84377548e82fefe4eb3d61beff04fe39836808fadf9407bb464be06b733c78a5f550c57c03e37ba005f2d5a4e939c83afaf3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h289e470cf4ccaa1aaad716bc520637f09a6f7c4f3fe806c11afc47bbf7c5cad9c8bef1b04db1263027150d4d13cb8d537ed656755db64c5bba21316b6e8e96d976e72795ea684b6c1d8e668e46b742e43c447684aa95904e13e6d6d92e40ae63c9f4651671d9e6ca228e85e0c7e7c1660;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc099c83814759ae347013ffd796ab0e3664c0672521bee28b517bfdcbc6671c6603c572bded970b5a85d1c098683d83ccfc3ccf22298aec93eb51167bbc991de56a6a87e5319a8a462654b60ff1123d377d13b5b6c90c86e4333b7a1a4b68ebdc368f315920132c6bd6923163d93cb94f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c45514d250f62444809d3d3e961d6b64b1136cf3831e1681cc6a80373adbc2a747393e519d37f3dc352f428ac04047c6b2cab37170d573f5a56d6ef4d0d805ebc93674f92662f7e00a02f062059e0beb09ba79dbec69f5de730f798cbb4516be7429900a42945ef59faaa6b5bba1522c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b2cf83cf5ab448053541821d5042fc5f05da68a2489c0e95b24398c4907d59056a55ece0fc97db0d3d1f16a2a311e6659edb306d62dfbc225a59120c2b94db09531c121c289be08d91f9f00ccd503c5fb21cb5f2bfa503c2b353f391553ae5eec3865d82b916864a09d2b039ad610295;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h332a9b7cf80bb291db6930096a39e2dfe0fe149033f1f011cbcfe6976551f226d1072b64636b8ec0f6203904fc9edb4dd7f589130410d56d2bd317d1bb10772870d7c5ba495b4d084f97b95dbf08a53a7e4c3b124c9992d14b81ed20f7da5429c4d1e4dd7ea73f6c4d7faadf733907b10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b7ce48ade367b8be99bc92f3188d254b0f557eb43f6d1f532f8e24aaff6f0a43229292cd0a2fcb09e57872c78c9d604badab8ad183a7d815e2316d9c320a32b4a1b94b40ffbca21a4a816475c5b54fcf2d45834ff611898a277edb036300fa1c2550093c1dc3f8e4334bb881a148095e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80f90345cbb9bfe976761da2af6a574ca89ab371b683809384f0729809644acf7c885d23aada704f835786a7a05f9b95557656e3a0600caf53bd65c609ed2af42c2ec094b85d0e1ef3a37947d366eacb49e28c1851ac97c867e2469ef66f6b68d0563827c1632ca8707e31cd212815f0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aa4e41fd2f955dba7e83137ddce25544e7b40f83942f17aa46dd94e23617d06d0c41c3ec3f37c7a11c8a03504684625273473f5162f8ade69a77c30f9888eb632b7df5af619ad3793c26f4830e9427e33bc95bb8e9ec1d99546480535c200497a83771f5a0bae5e8d386f1b09a461e66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7213dd420b98c2b5bffefa84d76556b8db9069fd61f4cabf5ff0379b0d3a9800f5b079d923d7b6835f869707a180631b0fce2353d2edb7a3a6c9bd33126614a0a7fd8f3b16f5ac581a9c5666e07badf4a0fd1303eeb2536ede0be963f7f0711597775778757ed1edc4bc4c5dd315355d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2050047f8a011e04f149ab09460bffbda00830a4ba1c4b9cd3fb19d997b18efa7952982a34e8eeb527a71e6d06b51e56e6f6aa35c2a587eaf5fdd57644dfbb720406861e3e258f6f7ced0dad25a59e91c2e9798f893a80a5bbdee58f6a8cd2f782bdb1ce601e649f02a6b81f4e53ab6bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbce2048099680a0e2a8afa5be8363f31c415d97b12be43919ba600ed3b627a19745219943cc39e31774b14b730fcade1e1ed271c4245f9afa2b27562f091dfc3f93be76e10c290e13060e575a4094af12990e010276eb957122c93fdcc41311c419537cd76443b5a04f621a1303284b80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53c3584550232b410a811934fae3a325181b88a50636ffd5bdc6d529b2c5edd4762bc6de029f625da0655809e9e33e18a558d6e0b6f43d007ab9b027ddc896550d09309b531f7b93c724079b80db7aa5b9c363ba0093a7dd3bce19d50d32a01bad4522899c13dab828639352fed83868a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h952ba300082d950afcf05559850e2d3f6a30b6473020217572e62453156344dff3c950e82a0ae732641f595f812d85d2df8ed0fd481ed83b8eebc8aa6176b3b9653a84da5d17cf31a1c55d5f822c052352c56719e994b2282b871abde9c837f21652073d4e0ffd7123f95190d693b98a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd541a434307aa28498b81c80f70d749336b4a2f866965eeedd120cdf9401a1b61ec2293561e0988f032c5d37c2ac1ed026c48821527ba6ba1abb4fe62dc720d246ff603292a6dfd1a450808eb79281de8cf2a2d316ebb9ed36390a06876713794e10127cea84c71829ec5072e5009a922;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0ecd609992b57a8a64b51c595322606a240d4554c2589ba070d9d93939a175e1acec56a11196fc5ed604e69d51ed55fca9ba1131c84245ee06228d932d3e218c2401d8fdc3813521a7f7d4439b2a8bad8ead4e579ee89a86fb1be1a0d15fd577d198a26bd111c1f981f30b6ed2c2a7e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5351e49a6922fb5162e997f1319de08b070f4e4397824d04979ff51e7c1b6ff39cc13e04b7b520e5a324d99faef769944e5fe4b8e93a87deed58304b39b4e4ac6891be54376bfd71879146b16df76a5911459acbd6b3d1e35c22c277d7d9f9b7f0760d6248ad49fa06203d832a50cd1aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc25113a65f22b0ed950a22d5eadea4284ed6adbf64ff863f43a3ca36e6acd295984c67d74374958c21fb36b3f344ac192695e6645635a2b4bae22bf41e17e423d62959472ab1fb1b03ab493bab68309a3d59eeb991b9df6e153d3adeb8be800b1033e230ffc5a400d931f36dd8ce9ccce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1650a3a9e30353ff265da848989201795eed4c431cb1ec75df1670bcd7cedd79b084c1528c6baad1238acc31c58a92498540764d1924fe209bd0e4404adee01aa8411fa556c26c902b932a8cf4a9d87175eba5e6834961b8486ecc17614cd66eb3d8ab51ce5b1439574c77cb2ea1977c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb60249c1d4aa23a579210ca7b54755108c8e3ac18968d392a87f754ee5c7875d263085d730da23871d0501ce995940f66a70711787786ec6120cc8ef62dae6199fc7397bb4995753993e17d39f509dbca5fda6246f7c8130b990ea3283c906846d5208b0567ccda067fcc0f46ff89094d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d7c0d33d9465d23ae112ad6afb2a322e0a29f589b17c31a6a833dd9b8b76f49efaa9dbd768d64d1c8c8d692fd1917d88a50fb7246b382b35ad036355c05007f7bc9a8f4e14b19ec4e9a3501f738bbe528ce5b531e3fd06540477389401aea7f2011dde832ad411b26314e4a315601c87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb16fbbc16c54f26e83679214cfeff7aca290e86a19b0c27e1a595599db63c387807f4a269b23180f8b83050cc8a0370d5800936c4e3f11441bc56918f70ec34c2177548fdde4d5dfcebe8c097b7e4f2fccac411325b34b3e93ffe5de64459a31bb187cad9db1b44823313a5bf1d84862e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d52dfac66e4bca81945384543d10b3d203ed42dfbda1c359a6622b008e304c02c443b982b0db85ab254fb84b6e5738687a106a39c7011340a68a5254d5d2408591fa88c506c16a4327ced1239187126c8e720c8f04aba0569171a0be11c0284eb9e419fa72e8ecfc27b34f96b6c57070;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebb66b916b17544a411ccc22e86bfcedee359d84a1d377aa4edbf4d14b2f68cc825de2f5f4bc90e370869a3d2c2948dad539660d2b973ec70bdf440d1eff4a089cdfa981f5fe522158277d00e31ce67f3723e7e1892d3c9a01e05e9742ab6f26cb48d10f5fafbe1abf351c7297fc576f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7c58e8b42dc4c959965bf8ff884947a03d6fa79caa996ea3576ddadfec2dfd156c5455503071bfd7cd5303170a3dc03332e18deaf464d0721e705210119353220c8509d0ca58aec68037b37818b34713a3b7e15ae59d4def1c804d32e2ed09d05660cf0a403a11992a8652bbb76c4460;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b8b903ee3bff8f98320545c5703d18f54ce373e9bfa25c06ac3a36522234bf22fd9cd0bf8f4ca76d5b95cbedddb66937fe6005b878b6058fd698d32086b5e2c77648e14b96cde3d6e871a8f0235798843875f18ffc9c36fafbf1c1f3f1cadc1532f6e53a06475b8523571afc6bda6c4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fbc4068f9466ac93476a95140b4e41fbca89d241235e7b426fa70c0e3624c67e16c3c460a4d7fe15fb5a3ca0c47a5a0e75a83222f9f2f537e6ce7a9aef7c6459a43796bcb5010bd852b92449ca26362ee83e11d5107987b14d1a9d45cee5227af45b47dd3516749dfbb9f79fb1f1bce0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a14f5b3d6341334e755fa01fe40c789d0cd5457b182ccf1767ec07d033434547f068acca9b20400a5dee6b655a1ba2c4850866d14b6a9fb43681226119338daac893fde179b7eb7e02376452f9863dc9c6d4140724e7120e26d7ae6faa2de35774a268687928efc03a25184445665bb6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48c4d35a8bb85e975223d071ef07b687746b44362b0eb369ad31bc02ac0b99dc7a44b6551dd3211dca58a4275ae7db36739a4b78cced5a4e0b35ef2fb1dc08ae41f8d3c380cc9a8bfe29d3d13b3bdd0a8f5bfbe00d2ff1c99979838c7d5f04aebe2e303e52909445bf7c3e4ae2c0f8d99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f0525a2f961a367a5423a58bb1aff6c9764178768d165da1f10a912260667c2195b94f9281fddfb9b89082901c61151a7f19482c77d30946fa1bdc95df9ace7758e830c00f69ad88a63bae1ab9ac91bbd28e1a05a1cb0f5201db27669a0e7e44e078938e4ac59ac30fa4993dc580f4e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe8043c7cedafb154352e977fce6ab7d07aede03d4920b7393e429eb5a1a985ecec2fff98ec928d4656cd0b0e34b66dc6d311bb28f0f2d890f427fb883064cb559112f4f7c0e2921a508e2d4f77c097b71a7284a2a5a961f679d4b01ebe265fd8d51a4f4def62d5df63ac3d2dbb49424c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b555d6d44fc1fc50605c9952c7bb1486a9ffdad245d3e36b031360e948b09ea45ccb84954ddb96f25c255cc19130b778290e2203a840842bdac65225548c4345cdf7d4ec3c99c31afc1836625de16499976844b2862707924b6ea81ee324f68a223d420f56d4a6b2c4f39b1dcbf3b7a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6bd68d574bcfe53a72219ded4778bf83b64ed78ec3fe7ef47665c2fcddae009e0323b5abf69fed4e9437d91f803e904ff58ddebe4aea8b69ad389266046b9209615755182e4868c9f8da7f6db398f23aef98ac3e8a7c157b62b8d91aaca18db11f0be52b07b60f36943681e4beff81d39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fffc9d200f1904e3387636c69f7df73e57207091994c705a8941af4fe073c373aeaa61221d9fa8fe47ea2fcab98410cdd3cc793bf4a58ff185a57547dcfcb1b25bbc53e449b95a8ed08df6a5f6a50bc7398466b87b95b812a9d317bb652a65d08d9a1e4460bcc3ece57a34078512e871;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40d120650759d9d29620c6cc7517a88665815ee9af9215660c2bfcb42f07633448bd1e97e1d1abd9fbf86b5de73d02401bf9ba371bbe4c363cb2ff6671c6969b23a3346a6fd35c5ab412d211e8cc084ebb79cf9deedc03403b31037a684e73467d51272d24902562219f7f20df9bf2587;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2ff8eefe72bde1a46ab0ec846433dc3d459698c50df847487c9065c03db859a8ab7b40fd78852745d82e06484df452a560378ba7e7e12280ad7fca585d32f592c4676365a002ef0da4eaaa7138d0fe448e91aae2e3217f70ba9fedbf95e96dbf0b8bbb15d8c58d1826a5ada8419bef1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bb8ac7b7d9968df89cb31afb65807555e23af2217a63fca0f7653d13666880c590023519e7cbb8507f0e63fd32ac7ffa24eacba6d2fb1a92ec5f48b6ca987cef0e6dafa25c16bcb85b59001eff20f804930f2606c9f134172840d2d43d5714ba954897bddea66ac71336b146e714601e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50c5462c71ac4c9a5eb20016f0c2c7408034b5e6554a24b188411e8b327d2e9a6c20f96efcf2bfb76240bc016b47e7c1b729880feeaaf6b7c7c1e622e1fdf11d26e53f03946e9650511d1a034b6d572b6073222971a2d1e89839b2d07bdb6b34ad581f65ef0c5bf5dbbef01a3fd23ff8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6081112028583cf5d10c6e7cf8097fb9fae6fbf341abf4cd7ddf33b563c6f0392534d4638d5dd6f4e8f649e9cef5f9272ce829278b8f4d6f2faf69625778999d92294540e723dba9139dab888e08b13eef55af9e76b4524401add31c086c02a3fc71bfcc5ae65ff7f4e3c97f849d874fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21bfa01828a133c03ef5c0587c0a3122840596c9d19dba881d4c50c9e052f7f918332af3883212aa900dfc0104a7008574197fec93cb474d119348743eb23a2f832d49ed2cfcb363470821e494721d6f3f5d85f8db9c4b04a0d6037615db024824b4acf15faa5a54ad9229fc8b3171bf6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd18b28081c289a50e7198dd958c5eb403b17567351e148eafaf6433efa9d904ac3b8788b63675cd2a12f9746a273e537b56f5f223c49aeb3c1831d1203db2e1c36f42d6fff4deb8ea14e940bc5747a5bafc015a09af69cbb32dffcf7f8216b68719a39abbc0d7d8ded4e180d7e0e17bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99f9e049e9e1375017c46bb25893e2c1490a304537fc6cc938bd10a9d6869ab7d56f6c4b40227d01c150d18f8d8caaa2a15603bbcce352d161c69d90150a547744a16e49df9591b06de7726c0036a391a0105ed710350a74df3f1f8f51ca3d02ce22da5ff477c048df75b5dc5f2779a92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h839b8f7615643152d2df8fdedd338297943041b3dfb9a3e4a2d2e1989b3f98f0228cacba1dd375adc24d6724bd97497e4816a0fd33ff56b0e8a906d02901090b4b136f9834ee702bce2e5e5e924a8b8466c155eeae92972c996bd6bc547844199598646d8e117f3ed2a2137f19350bac4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd63119e9e2ee5ce78084fb64117f091b3b2909c2b344f5b5dacad75a3fd865835b9712c262f10ff5271ddb5cc7c9f677a6fb0d7f27fc3b5cbf85fa89faf4726f60cc84d983221cf5308db2dda8cbaf636ee6cb3b8dff561ec90d66b9b51087635709f930f40c2f7e43f92cce5295043a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e80cc5db8dcf2cafa9d90e81bfe755c73ab7b5e78a30ec82a95d2418d2382ea1169078ad7b3e4c1f2312c75484af66190f4d9e4f40d5ada4134aad2b600b36e9fb71ccec68ba60fa527090446788a7358b750773fabc687b15088021b0b1953008aa0fe915b328249b0faa939a84554c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf4d03d68908a598e4b316618064aa50059ddb973e54c280d97ec5af262a9ca28f88b0b8016632a26ced0db0ba65353e537ced11d3d9615552d9f0608830c253ecf919a998081dbd0cbd62080e7cb8695e7cd08dd026171d04137610c919298cb442dcbb1cdff21f5b417a119dea5ff97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66e866fc19a51fa58ccbe21433e435c57f5c9622960677ef9a6d3f6e98ada5a25f4a26026de76b3846a908db339935c62332e5b935808dd381f7f781f92d36ec3d9619eaf309570b0e46de78bf948d5c2f816160d025566fcb13db4d2e7efa24da178717b53f71db3e6c88a1833a08260;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e2ae56a9493fd8738e6957fcb4182c1032f618a2879c9b830bcc57212121bd87a11b7e5a3e2cc15ad092846e932df67c33cd5be850f2ce8cb001f015ccb449b936af61d5804b11f9103a7ba785c1d7085e0a8b6702f46596bd3bd26db5e749ac379514d8f0da9f0ffde4ef5bd54d3f77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h404162620ffb76de4a0788fe4bf0ea09b4e375cb323b69b31abfd33eea9012001876a2e9a7d1f4073956388368425d5bf447da8cf8e2bded3da0f292a2cbf45dc92a93a56995988125385b16daf420adbbaf640774f14394810341530c75eaf4b8931da67edd1ef8df63f83bb3f4f855;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5789c12f48e016e539c6a506811b37474bbd2e48a56ce4100d578a02413d9f89bc0375a0f17c2cdfe2fc8d291a02a0c5dd33fd90f0315146cbbd055d07a59e3b8813950940ad7071670cb8ac72c51df38582f86c44cb8634abc10ec0b939d55369c8bd6d0badd8ae505b916d0dc47cdd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h750523bcb813b46c2f1976a92921b2717437308c2b93435aae174ee3a5b1a1289a2728b1d2c6cc6246fb2d7bcfd4ec4dda774da2ea3eb0b375e0b50eccc960d79e876fdd869c7006405d56b32bf9e75aa4e8512db3e3ca1ea0ecccbd47c288cfe1ea595fccc1216365e51ac2c72b3b9a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e8d6e188415f178cf404c1ee97b91eb3dca6f0fd2db9726245459523c114f058cd6466abde8f1f8854a1f505ca7fe9543ca2460c914e79cc9044b378e103af5fbd15b09c1b208bd320ab69eab786322a027c462a0a4395e4d4b9d5c3cec0529401a7ba4c93743f9939085fdce1b00ce6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78c0d254ecb5aeb5365e2edb364c6cc7b317b881ca8673a7a98b7f1c95b2e5824980348ae71c1b19bef0b1e84c22bb259762ff47e087a76cf9f5045468fbd178d7cf7418d157e0a79eb85b77c4ebf7acb6197dfa349c90a9668f6cafc5b8494885b144c40d2f73174d6de470af96f5c3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c486f1fcded95cf06a23c9b4a839bb5653c2089bea34336b9bb9fed42d96b495b6e5b93d781f52cb9f073c869c48d529fe2d4c11ce9cfed4407d477a4802e1b6c9c82fa171a361f5602195096b6d4715cbb517f9b12e3e34d2911e306ce579e270ba6893e32e1ae8a51fe2792300709f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66f3a064e0dfdc5c8f52c91c9acdbd65fd6be589522d31fedddf5472e2f1569200effde2039acab33e2c0dcce014b759dfbf44ff67ed6532fcd81133dfc7e4bfa34fe5eb3fa6d473beaaa2a8a2d11359e6012c220c11b8ebeef8280864c0e71807b10a9834ff205d244f7f554bfd014a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f6a6f9e8ec8785ee5fe9bbc7a95587035ab4b9359a3cc635d2ceba73d75827a7f224e696578eab6c3c66de1d24c3d35f21a1e67d1e22a829a4cd167e5e0783267ddcd0af4799940f8f3b538d40683ffbacd75d1c5e7ca9c8886a99d67dc0bd1da62886536e37052e9951ac838e52954;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5ee77dd2d55ee9b70b77fd668355499e07e54c1e2a1acbaee1dcf8d62a20f51d51e49ac30f6775157bdf0787c75cde447f5572e7cbb55d538c569588080f12a88d8ff6ff523b3de65ab86b42805b2f1f63fe588738a270555ae44ff3156bd69fe3c1ad1f7db239b080a5dd4f88b7763e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h439a94919a7216f7f4830625c27b95617e339f2b2d7daf2155a1a287d1f8bab6ad0c38d3bc8b0f88531d1385ceb303d6ad362e4688471af28ce4a82db13e0e0f8fa00439fe4d39385c87ad055ab745e1894772e1762a5738227303282bfdbc610ce822e2093a70507a0d8db4cc954a4bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d332d5b1eaedab7039caaab094ab6e61aafed19ff21f76d94988b31a1c41cd4d0104a57af1828fa8c60ff91cd60404b3e43035f2c514e613af4e29f5f5a4de921b81e530ce648ae887974ec75fa2981149e8ea06b81d65b5f500f207555d751bf5e7b4557a826bc7b26aae0ba60923c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5231d35d2a074763845dfd7207e069f18ad62297cc5d138dc25c9c16f57fae6d4b437d453e1427a1ec356334e161089cdfe26d17435af5f54adcfae827a8498193586d7a90110ec54789893b42adb44f565d640c618fc31cde5c38919569797d4bfcfba18d8c2badecd307744480ec7f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafae33f3e9e1969fdd9d17abf3d8ab8ce6cbecba880520b2514143fd14fce3a3e4d510ea5bcb2c51c3146c620597b3589e522d258120883401661f55d0277f687892ef9b9c9e0f424a78620460e3328c3d76679ad8e479724c3776ad5140547b575ff2a3d5400c3fd53a1fb583acf083a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bc4dea6895f907af59bd1318d5f98f7dfb6b866ff2bba0016f4f6ca1552a9c67877bc5999291557ce1040c0e91e9713a6fabe0d3d6df721162df368b629cd76242f2423500d8b445f2669b04a7b75b88ffaf83aa151c17a062e2a27e9be42c6352f4c9e9db7c191c6da400fff251cd12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17c5d24e24b2e042bfc9f4c863ddc95c55b2b5e6b541e40485d3877f7ee731163c0cab29d4160911e01c1495f8201158f512391885e25cee2e5d35868d7fe69054acbfe0027de8ee467832b3fce7cb928a8fee5eee4bd7d1d403fc9260c47ae566ad36d51933f2dd6db557826cdfdd35b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d610cfb9e764a370fb96086093118f57d148130201a322f885c8c01d9a0ae021914bcc779508c073eda10f3b9ec31246eeb061af32e830c0defa84e46f9a93d9b1293a72638fe43081545673998210e150503878796c163d4806a777ebc39fd4f5a7513b056f5a8d8b9b518eda5220df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33ff8d50a95967f75f588d78144c2db97c4cdcd2a1aa04af251d95ba4a3fedf123f0a3552f2835ffdfdc5b656d6ffe2bcb089779f1920af1764a01fe46fd8a1d5d5d3b8c655fbc1243153535e47736067540ecdae9960ff2a39d19364837bea0b21e71e6cf428121846975989fe181983;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48596c6709380ffa395460cbe2d5a04e084723d04f0753565cedacc2372496d4dfff4d96ad39011ae76280ebb4ac3812e24cd51b66fcac2dd024a493d110fd32cef512774d442bca75ad5da84a1713ef0702e10af9060b80a22ebe85de1085e6dccb589d14ead753fe728bfbcb214b0eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93567ab0ce867db088d241c29d17d318b0e9dbcced382ee1f1a34dc251b841541cb7e669896b588ca371a0be5475d711d13514ea991eb7a80d3261d1219e73fbcfc8bf54f846263c0d78a59c0397aafd1c8dba3b1cc5f4e10a7b00f4206ce99e9e347cd87a3a7102d785c9c871d523899;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb754b3be2c638f154667c80d99883defcc0c32cb3f152d69d9bf63be182b86efd7944e086e4f4bb375771652ef4d2d084af1a7f8eed9fd5895fcd2cff35b4c570e3ecdbe4545a50c602ec9ca495c453c82198f05e879ba7b59d0913de0cb125cb276cbc69318caca5843923e18331c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h392b179e021804a31bc69e93784294caae6ca71a7e7d738692f4beb1207209bff5b772a9aca3e2a7ab4bb5e176c0abdd270e4e5c67244f869f2bcec4cf21ea3d5bbf14abd0db6f01bc1f04f14c83fe2efddcdeec71a5548fca8f11ade7fb5422a0cc53cb4958d863d56c398952844012;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc2c27b8ac83d1a63911cddcbecff8604e580f1bf5f5759effd3d24f1ce673f7b485d9a8b67583f1c730b237d126932ba7afb71b17cf4be77fa32804383a46bb4bc648968722eb7bd42ea8fbc43a7bef7b87e4014499819056b3ce9b51f0b7f68efcd4ac7ec544860d062d14dc1ed8d82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88f4b4d13f99cfc3b4f42b77f3aa5dd57f6d50810b931c24fd5564b973168086e7fc5881eff0b8e26b100bcf69a2497d0c598a2e4c686ab43c25311ba9c39800cfa159cd0a7c84464c963d175f5684d7750c437d1ace35d902de72f8adcf3639b2d698419b6230caf4fd25bc9d6667e40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22891683a5a69aabe0dd5024e30d1a6f211c1fc7dd2a5769bcf43e9fb7f1522f6f35494053b25e8b36622dd1f7b29b25c1f5a8faeaa2e28810fb97ef98c8bdecbedf388adb85bb280fc6c25ed6d81efe0e3aa38b290dffa5d7af8b83a06f111f8fa957ac435030c83cf6538ba27a39031;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddac9cd15332b2d3c4a8b6b944f08c0f6499474d6c2111edcf17fc73acc82a12e888c310dd620888fe98d2c18aa0795487a6971063c20cf9943f5a00b8d1a16766a0872f2fd2af0cda0c93652892665657e000a1980c4682f98997888778d5eab0cf63babffde78318a20c30841d26ac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef89f564be022b9b7ba7219b14df07341eef3c453d2d06d34fd1bedccbb410876c0c49fbe24688312af260d07933721fa045563d15a21c317ba709495092834671d37bcdf39776f789d7a04777c1ef9b4b509a557a992251004179144289f28d9657317e9c0cc829b47906ad2698f1060;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3de70c1835f5af90ecc01f091a1416f9dd5b0493aba7aafe4b49dab308895bc547d0dfb30ad71d397b38277e1271d9480972ee811d805e9f22395b832c9ed3cf0fe5bc0a94dce76a3574b97533b22566c555137cf4365be7f2767c7b692516b834d84b378dfba105f944b22adc336e0c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc25d9fd984c92857c449a30b9f69639ed7a9480b53574a17f5a19cb738a011fa77bce9150b6728ade3c192ce47e7360748273637228ceeb1acfceb41d6fcb54c13820acb8378dc471ddf056d25346e6c5391a9a24ba2977aea6c5b73c11cd660415409dc23541597a0e5ecdbc7a5e8b1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ecef9c89d7e184e30cb19ffeff9ad05847736844dff8432d9c2267d6fd5c49fb1a05b94f14322c23485a072e8ab0dafc28f3955ba41bfd34d258ad08e21e355baa48ce5ee18413a4e05b46be40beea7550e5a44a36f605f102f49f5e9f4aca4078ad9f735462ab6664ce3da3c109e71c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h166e771b0fb4ed45618f6a41194dbf027e7c82f86e79cd1e16a9c21c2ef2712e8902c827f802f34a47fdcf3cf100bb4f3608ff1b06086aab1391499e07731eac074ee423c99261515155ab9f7a1775a27e25fcfd9f45b200ea82988093a1cbcd13a99b14e44a3d5401121c565414342fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb882ef0528ed959c96a24a63a761a77f67fcc4a3ac449de6ef129e133088863f21a9f13bca01d163e6cee75d83293606f397645e8ec87be73c680916d6395e4c4c7eed89201d1437015859ba44b41a4dc0817da4f388d2bb4bde890f93e77ca624ca93f3565138b4d50dc43348b6c10bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb07cfa1286c7cade2de338eac70ab9036096647554cf0a83787d8550a11b8077d459440b9a2108b9c10774421943c002017154712c83dcad2164df293d237ac8cfc7d10873c3782bcc97c34de099fb9ef34d1a35f72244c415cbbf6867162267e802f70ad2928a875a7986cd7b58703a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a1434a06ca64934d0165dcb95f77241312e23bb480ff7d32687d2b53e49acc2b2b735fe5557a87c4ba29853e4c521e46940e60e14baec2c04bfe4863d0b0d616d090fd11b64ee410cd3cf57e2ff45fdedcf05bf7f382986e19e7a24daf374b35c486278faadbb43b5b18c539cb2828cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h234bcb32e9c172bc7ee390e0177f533ee39eda6ac8a6fb10913e87cf0a6c5a51e420cb3f0ebac436264876645e53fe9b3103b4f809e4b76493a2a214d26e0d5d05f7c8b181553d283aa3d66f7fe92c09b264c5bb08f6ef74d2887be35d95ab765cf585373ff618224fe0532158905de86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94c3c65b8d029bb748f54a1338cd81997d70f52cc6874086d1a45b117ce8565cc6e8fed9f9f7125cb1192765b7b03c6d2f0be14a396736760eac932e42ae1694b58df46ad7509280d28ddaa1fd6ef06251b493c9b961f1b9a7138ed2966a0395899ade31d14d8c527d3607d043519f612;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c0666acb95dd869b0496a4a0368d712d464a82a2c0b584979db42c81ea47cce71b182f9ad752792f9cffee005d387079b31b893ba545a4052e8d4c8d647c5976d54e6f44e216e325813788aa85027e016323434afd572bc738883d8195e240dd43e33390b32129067557bfde3dbf1627;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4284933621868b5e5554d1fe94b67786687edb2383d820d85e711d1ff28c92a9b1acd3f91311163939e1d20b9ef360178dd1e8da059fd0b2392440730252ab5d9cad2bd640b9b1c676988599db9d19ff2a638ab7725f8f34abd080fc673185fafafdc02a0f6a753b2fa6af8b1965f49f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbe88eccc80454ab36b0536aa1bf9c11838aaccde53d925025b15f753f76e103905b3432ea0a723a4ac9ba06bf03c73ec0013465b3d790b4549feef50c31ce6ae98f5e3c6fb0c989c771697f4b411703adfeb36ca7b4b9d111862378d28c3aecb6256340b4778481f8e6bd45222d9ad6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h831fb8f1f2d4faf6390b38bb13aec713fef558b0ef2da0a510a64c2ea7c4243144c7ace6dbbe9911c7269ef2e76cf3a71e7c23c73d010cf1f2d74a9209bb8a9e74bb3be21bd576ca71f21bfcb77f352336fea58465557b92373f74e92c6bf6f634c57a322fbe10c9399a7f3a9ef517110;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7780fb38ad1499914758691ce396bd7caba7097090c0465ca54af09830bd853d1ec7c8de7e0c7a0828b835a3fb03174514c7d718994b067b40399d29290135ea58d591485acb424d59cac41fc6fa2d6f4981ace03338a0947656fd76aa8b7933283ce8cf993547388cbd6618c231a0939;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92f73e0ac99af6fdd508f9223762f7fff236663b57852649b86c2bfbc8a30deec86c0ce93364a2b19a91507309dcef6c01d10ac90b1302cdc49cf1baa74a66bb0783a999d9fd339d923edd03693a868c5ac917ba51400029d19df99f981652b3d4ecc4d4564deeaad6011154559ed1124;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccb0143cda670035c56b94f0d4ee73647ac63cd3d3ca4f1d143e9b4ddd315076ab4f5d4a44917c833d8037a62576eee07c561238ff3cf0dcd33e09bb3196b9f9e31f9c8238ced3fc5910fd0892d011842436cc127e409c91cb0d9d21517cbdb734237358aec49d9ef853f0ced86e5b6f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecc24cf15cd0d3050ceb185a4efdc71c945d6629c6d0fd525fd2fb78aa869d0415890762ff2a1ac7462e835f7704bad452af9b62d8ca0f085af56259c276800e7b61e50302a526b3b19f2ac83346b81e88f7843f0f3f117c099c7e7062e91abafc2c39061be197f592a6d5d17bc1f6e0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8343170ba5e355bce60f0f38fb1c649663a9cf076f020a209f9e095cbcd0df23b53b3ec557dc773da89a84a382476a05066b6056cb67271ae3ebe5899c51e9acc0c6068e4574072ec3464731af7ab25f54de47092ecd51f3cc220af0afaf4d03529de48cb17f54099064791457faad7ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3f091ac7de484658f5c0a1d2ef1ccb6d72cac12a92c9b4b91af6b606c284c305dddef029dc39d751d71131897625601674a4bea9d9a47e5559698f1f8eb70b14091e9f623114ab724383706c88fac1f2743e668ea9a1b78c1bdd79b04e335432e4997dc05f1e583275227750eb75a392;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd46a8d4cb0a0043bb9d8980efce63c9e4b06d8717c16a4e8c64abe8e9350fa3ee2d0eccd1d889fe14589fea4b76d3d2807744155ef20fed1de4c78eeeec8a93c8379075dfb5f14d294a36f6202a9f11f9817693e4a3869bc0b09b0647c3409ac272cb33cfe0a795ddfb76df8744f31f44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he838353e1e52fc367605f8c53dfbdda263cf6159ed7ec79779fc79f8b6aeea97cae54bc72d5ac7bd578a7cb9ceb0f14645f8ef43365ac6bd0a9ee18488da52914b563bda86807efd539a4346f85964ee5a650213fe29d86b18de56abc1368e8d7018cc77ebd9e821f99b16751f78a36cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab52f8031a82b3b4d7ace23af8e15da2dc588182bab97696aa40c6f353cd78c8d9663e8afa16991e23182f79f76fdc47fe19c476fdd5be7ff3d982b83f4ed784314cdfe2453df2829ca3f8b60b444345e4d85928435ed41c2d1c9b9d7aabdc2afd4f327b53afa2eb322a5314e50f55264;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d306bb1213a29173c42c4ee542206636911151e05de8f58e9998902cb71526e552f1e87e2d347793b729cb9124226fd92fba4c420656648d92da2b32e57913a6f7e7c6a945d04f3897a3151118bb224d18fcfe5a476c334600ea43eb21a02925a4eaa9cb2c2f7dca1496a4344c288b98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he82eb81807ba6a9a6195adeb2112286f657fa98e5b277f05996ccc4ea0c25beed95118cc17576b38c17e9b45f3cd55664b28c7329d6c01afd374945d1682d2196f84a0433f0a0f33a557f110e6fdbb29b6a536eed40aef3ed2d875fec4a3ede91e7d48a8ee52e45a55aff6cdc804700e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6aa4b6de582f5c999cc9378982b0a83709e6a845f6ee555094fd8bfa2845b6e4bca568f61e0542210f3ba203fa86ececf41261cd363ed9cdb0463ac0a4ea86fa7c13fd7b330612cc88926fcc85bce4876af7f1d25e0a9e6dc82ba6603eb39cad0ebcc93bf92cdc7e2e7397688347a6431;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3866a9a0ef396228f054f772cfdb6c149a59de9f0c5e75502f19038ddd3b7f47ea38cd3d35bf7d0b419ca63f7bba251a942b26d456f206c19b304e48fd36b64cdc095022e4e38717f7af64ff647c8db10b286aa82e52c79534a67e6567de34e9213fbdf952146d0831948f210275a22f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he08eee8ce72adc2d34aee5b3271040120477229873c7aaf7da7d050b1c1db97066326f30cf1b66c458092d3b18de1289d1202c56600e9e975bdca10641737ef1948b784d5790b293605d88b110a42d7463c25668d4a6a1219143b8b55b0cfa446dc50368591b0b7f165cbe64854a81f19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc93c62f60ede8de41757e8f285ca15749081230c1b866801bbfe43e038d2b16acb445214259dcc69a26c09a3bbfb4bcbbf00f8c746022b2f958d4eac686551c4104cb3e587eb08ebe5a395e20103ab75224c0227a15ec538995eddf128945d065b75a18d5747349d05fed98030655df65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39358c83604298ad67050d3ce07afcf32b4d8da2e255175c63e82d4fca1acd4b916bd18dd6ff07af2cbcd4f62383ac8ce3ca487d177d9411c40c256e33037986c28ba35750a9f4190d2b5c95f0fe09eafae7b9718c267a6fbdc6056a417636f1e8bbadd60cd4f2301938e16d87d1e655e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fe4dc72b2080c2ae14938d496b9d192c5a71897e4716f0366c6e3ad12a1fca513388030343c2f6ecc0e96e0effb35bd8c232d6d76c031aa5e285fd49c190fd7a17a54669532766b703b06c3fccb6d3be8b2b20dbf5972a49cbd7c01a3d5566540facc69b202b07a122982663a9e640ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b43d36edbae23f26c78de9b4f339cab91ce36dc83566ab29534b4c45dabdde99e7aedf956ec3a88fb26ed916d1628ce61275866fcf5b536a9d636c4bbc16511519ce497ff8303d1bf412339b841351e236cc49d0c78a7d21cae9bf883601f4309c5fe31bedfb28f0e403a1455767c072;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2815fd4eba3b2134b89185d7fe9993ed9a9c5c98c69d1cb725a9675ee12cff169a4fda86e70ec70da99a3f24f5cf98bd55a2292d509459b4bbac90b06387cac2de68eba18719a1175b783c3d0669dd956d61603bad80da9f418fc70a8d0984ed0bc5431a59a89e65b3e1b381d2b74aa5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd38f0bf089456893c2c6d6a31615a1506c4d122f6a066274c19769c16e6338a56622c2ef8709d58379f9465bb35f4971d7641225ff8a4bb64d06a6b94d50fbcc2985a73626bb72306c23b4b688d1e33c481261db545972e494be2550edaabf20f106ca556e5a10415e797f714f283fdee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde7fe77402c2f39d2868380b5b12c900bf38c85d7b00fa582ebd7402759da37a6fcc7c8755c27bad4de81ece31ad42372411b38e1ae788f981fd0f9afe21839c1a06ce2f64ddc29c09229c38ee4f1201779e9005a3207ccaa099e283465c7bcb32f9a5909e391513e5a2f3683fed05283;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45f19c9c1eee0a0e60833da22d7932e3cd7f2826c2f0db729dafe8342c10fcaf1f61b80f91377ae4394c288689529c9b6a8520bb80318d7e2ae9851f95955849fff3bd3d4e1d6aa37572097f3379751f8580587b2c24999922a481a63a1c6a3345393d8eb5dc263dda53fdc7199c9e7c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98183acd921ded7c842967c89757019b26b3c39cb0e56f67006ad3f22bc5b092ca0071462ef1f2449dfee364457e50518891a2244118e0ed9108c488c2a55609313fec1c0e946fc87a3616b847b0cac78ea8dea9a8a66c42f1b558fa05ce682409cf7ea388f6ada23e1645c9cde2dbb1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha37b355c0818ae4596b09a9854e0bf5cb037a072085665d5dc79eb4d8ef9260d120e432686edc283ff059ad2c686cf4f0648c5311f51c1508d5058d26a24322cc73b83d971cc44bb22b16bb86e9e2ca27a5bfd54c1445c58025a703dd0aa01a2b7a332776cafacbe059bfcef22b995ebc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc145cc2241968ed3252a9e55608776830bb1a28ffada3064e8d597403d01563d9ba69159178120753ed365b286607a3e0e90ae48e6ae6b1876d424e11b4d12ee2ac6caf2615034e743663c5ec86ca761ed5deeb776dd43a7c61441780fcd82370857e95a3cb99d35673283fcdc88f4567;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb13bfead60670e86b81d376ba3970fe4342891804b56b83adb4114b60041990aefeda3bdc6df9fbda1b1c249cee617cd61f1f7f32f2a1b78dfa7fb7356427638d53c289b41ba9ba578f337cfdb630edfc53bcd8ff7521fc59ecf18116f43bd8e9d659ca870e9c2a9fede38fe239ba4b33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d69e955b3793021598546394ac5ded51d7dabae4562782c7ea0d23acc598db4a7ba559b765f52362db6be675f09c67c0f31f3d1508c46970ba16043b25dc410d05d28bdc348579c31d4afa49f1fe694a63baff967672355b2d7864ba2f1171933c053b65dc54909ad3e16e3871460e69;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5efc83dd1c79f063fbe3d9338f4119939f1ea7a6277ce0bf1e71e94f9918ae35728aacb505053338ef2cd84204bc8db953813c49ebbfb6b3051730f8c95aa742de8be08cd4a3320f3980b6ec080a0b72415189f31236293bd8b551cb1741a31b0a5ee1640eef3374b52da8d4e122ca60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91c21cef087ed8378518d6c40d6d525ce0f643c830931c43b718d61108923d5003856f4258dcb92fdf73e1442dadd0ad2827414276cbdc4d10d250e7e9a31537fcbaf4facc201797a70b33780f414f76d00d6f0faa08db1cf149d7485fda29e4c07f99b45a1ee709e759f6d17e4cdbfcc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5da6b1afc67794b8469587c812c509f5b5210084cc1c00e0738d04dd743c571b7ef2322f739b58e16a11278ca785061f9e2c08f08d1c6ba9030a12f8ef3ad8542f9a493baa270673b6bb5b01d2d9b0ebf0a4d50f09a7052a0a66eedb38bbab52d877debaefd4bb8e5ce1cbe6184750202;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b01848196c0663f0f3cc2a9ac71c65e60ad3336ef2618c85b552c226c53dc13d16550da45310858ab76fe7eaba5d03c5aafa148e56f26370e6a46bd6ecc41c19860ffc74ed592c41727f9e5dcc91ce4271220596df8bfa558064b5e6807b1f265c7711c022b14c6b2cb42686c151dee5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcd1499857d961cc01ec42147dfcf3550a84e88abef0ae4e7e98e548474af5679fd61eeae15baafa9695f841763bfbee66386194dd662bfe02374967a43d6f27d416ffc089fee7252bf82f66db66f5d50741cc0203e143a6de3f3fc6505eeacfa5b6270a04623e93737f1b9dd31b27861;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17cb86ec8600ac4837dc9a2c139e94c286b48707fc4730c462958c0e3a62bd3ceb7ec9ce6bc0d694286abb2315e8825fd929834f64602160ac13481bbbf63d5e8302fdac0e474584c2ae7fa911168ea3771ce05c09a48f09afcdc2f3d7e079d7192f5276ff79847ff20eeb696ae890c9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cd9f781ef03b16b7263b1893560e57270886dd2f50b80b02433763a921ed7b30acded0054dd172be1a5e283013be0c63377a32b2486a2ed59936e52a2dbfee8db1faf941593ec0967685cd8ac223eaeb29a1db92f77c598024f275e53d3cb0722da8b4c8ec148264032c0f8426a59388;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ad08540a2a48c25911c0cdb57addbec96ecda35f81b3c21b1171453a537bbcb94ffa14a0df6850a84518fbbc7a840be4baff0ad802a01cc9d04a0885ff008224bcecc328a17329554b86d7a15b60146812e45fb3da2d2a9b5dd0b6e13bf385a44f2135dc8c69e3a1317c154cb3fbe390;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3943187ada4df6ff93fc6ae1e89b925a7e66dd8da1d27a3b923522d12659d7bf6838223edc54fd4f79e726d82b960e674a7f32ced331c48b5295dcdfc82eb79683763aa296d1652d5628fd170236d7b9312194e77740a9a53024f09b3ce48e41f6f4aa87ef7019c5b41e1e6218e1aaef4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heaef802eca0fe2c51f9889f188c03fedbc83cfdf499fc2948ac4bbec24dd126873a482ada95e0682d56601a2d4cd2134f8a40867cd103fa666d096053441f31368c913bf296aba34486cc52980eeb39ca08b8ad368c61b18bc4cf1b929180b55b342a2cc73c160d234cecc1baebc89553;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ea2d4a0390d8e71d62bf2d9056604dad5ee306a4d77b151fb473a85d0a9d78f953dc328575f42743ca5c16e5a327253655c90237b38d7d146077b6e4c01da11e4b319971d14865496345dbb603f2644e045be9c429ce38ca655e4759a073d99da3b1214cef913af809add2f31ff59d02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd11c5a709747f1ee93f3f895a32051895fd891ee11d9be7c1ac2ccc266fb97fb15cf860105c992b2cafadf1f6e4cbc0122f641e9ddbee689caaffb69f34dd91bcd7b8e205fb7e27d8afcf50a7f292f9ed18437369315402769a56b3a0247a98767f066532237495c21bfe32bb1b2a49b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4df97ebdbc306eb1e111976c929eaaf9f4ba9da325257a5fc77dd9430461eb1a3019f56837c36f3930cb0dd953f5244cb93e5c55bf0b14ab1842bdeb6770672959cf58f2f2fe2e9492043cd69c06d3b36f9b872823573e47fdc39d5835d4900d2fcacc471ce066b07bfe2b7ec7ee1fbd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heccf45b640322a8461e2a0788c151eb79f3b31125e80ea84870c328da69ef6bb2ebe026aecf75deb085d82b9e0d5599255ad4c1f1f844b30225854a143a7e4b800469c23aa21e582bad6805d5bd6770971cf3f17106a1cdc516004c59d963e2c76a35c571eb74311c9abe4ecd6ca011bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd65b226d554e3651932ef4ec0608e7ca390b8682f28164e270f5b2baf41a1c8ed88182e4491b94a3621bb580fe9036a7dd7bd42e8ce715ca27dc4707081c56179ed5c6d12c1bfa0eae940954f1a2491626cc1478b04539dd3335299c878e62797164f5a493ec9e0513ee9a99bf7feb0a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3f4e5d661e74079115bc394b57f9f31a3545ac1324f23ea3c2a8586a63c49272d87879f72b3817401cbb8c8a86f307b11226fe2b0ede6f684f52e5c2654d36c18917ac87826fbd5721432374fb26335941bce145017f7f58410964abea1ef799536751ab2e1c45c6de78b30f18fd0a0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2886a1a96bc2d5e69fa74844d8c55448e4c22d2c43cb81363d7219898217eaa6473c0a7c7236b5d5e0bd0fb99c3eb492b315c094ee8794274c7086414f60c5f912833c57ab8b0949ad4ef9f3af995c9c37e6d0de151f4057ba19be99c5fb22106d1102da43c7bd0c79b06249577d95b79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed5fc3e17de099e1caf2548786bdfba701f5f1baf158cb714f876555989f4e224b75f46df7696de37d584ae80c355024b9ca6d5e6e90aa23d380db21db467c47c59dd0c7bcb8b61c3fe68975fcfb15231843ff3347016cebf6956003e8423279afebf7887f56808f0c570a5b520cd47df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c35d038a1836088f6b3fc0a0019d61945891788952efeac00347d065250f5de249ec7ea0cceef0c618a185e3c80e597ee496616c4ac703ef42d66129558e7d5c7499bdd5675e016ba4007106eecd2d8ef41d0d521c346cbe53c1bcbc6371009acf57f0703255afaf89336f1eff8450b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f5857930f452f505526e353a16d76827e8e8e5d921784d5fad0aeec98fad7ca8bb23352694ec995e059305259b3c2bf1b998e2af9eee85da02117a201542ee0579db49a5aea28372d59caaf7ebc85890287f1fe3f77eb3f608c007f877ab9a06da1da82246fc7567ad10094267f756cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39892e60c6b77ac150439bab1dbc25fc1890885312db5d8e00c91c5eda9570eb1b93455b9e466694f494664689b62468bea350c478096705cdaa23b3b08ab509e0e7db775519332b8f1228333db44402780d53496f847d3b0b99d06a33f84914a20009e42885af3b39ff435ece46cab3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35075d1b494e1389a09a093a5a2362ee7cf550f638091d0d048202fc70ea3668cd003f789d51de7ffecb9deb2f74567ff65831750022a71d429b80bf4d62de367aa51115f7fb3cf357baa52861c66a3c067eda5f77b54b639670537067a556ca02a047bc308ca0bf9e6fde5733ba3ee61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68a2d86185ef25ef8d90e64ca92f822315e1d81a6b310f421e935ccd91a40b0aa34de9fd32bc283d42b8439a8b77903914e9675ae696b82a29d6d25c386eb4f95c6d94a1d9fb9333a7cfe90edc48ecad629343d4466e24499f0175d8b14793aa69dd2c1aab3814acaeb5877a07882c7b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99800d111c2ef54394dc5fa75288251c0d9b9f6bc5eff108588a0fae04ae3b88b217cfbbcbdf6e8e5afc07a439ea2f88dc20aff30d8048c95e6ff76a47e70b5c31add895fb3e767299e6fcf7744cf4c6cb2c946078f4baf585069eb282017dfd7b70fe15fd7c278419264073a37c01e19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4eeac575711db57d5b8290c0eff8d96adbc34e7474ddaed961a40d1c69fe10ae146a22df27eee150adda68ae2e9f1e8e3641d7334bbd42d89f8c2024b9a7ee4da7609f8eeed14d7b6bf5f72b9a130bc95e522ff5f2b14c60a2bbb57858e51ab1b3e8590d58a536399067eaf6529c5949b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6025787305b6ea16b3b4eaacdced9c484c63a568e83a86f08350ab702cdda9ff03e2daf3780599b5bac9d8e3311dcc0667fdc960e8a779023bbc3bd5429aaab27e02ed22961805f5485428143f6db8047bf5ecb51200c9f39feea9feeba7a16056ba0bc3bd6592758c3a023e968d48488;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h725281054f2088485ab0358b77b9633de039c48e9703817a4d1e9700a2edef4d89310e7338740b9f8582eb3a6139368262dc2fbde1a81b3352d19459e1ce035434cfa7cfcd3677facf401d3884f6f5576e88d9e73c3ed3d5ed3766e8d4d944f430a2ea18db4da43cfbfa8c5631cc4f5d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb3117b30dd5fbce0d45b8d726766f90c22bc8f2c3ff38d34170d0f19ea772f51f5ffaacbe5ff5bb64701933e9417df62a9455f146c4c982652a2ac1097a132b21afa5e6f9c7ff5fb2c5c8e65a6484f17b90b4f80e16b2a6dfc15b15262bdf909ad40c3ef9e7cf31b4ea30387d8f4a98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h212d2c5b9a79c3010ab62bf372fc1e542e6f3d225882f88f558225b2f64378a01da9e817d84bf2230e22d4a201c193d9ec095e9bf32a82cec593ae67d39129ee77e5929d8eef58783a168b05dfd3a42c125b59b43cf623723b34e9065338d8dade794b43f938c2f22211f39747891a7f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e3fec5aeb732c7d895bda2b11fd84d267b464fdb2182048461ebb0104516bb47490f1e6eaf09843e35ad2a49634c0ebcccafd40fcfe87be68547e178465fc4085ada2f4d24d92653052c8fa6a0a5ee626eb5716efd59291e3a0e490241e20dec2441752b8f0df2886469d13cb6460e56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h899fe3b68379f1851778ce2ba8f93c221691d5d36ce38b6dcc9c1da2d0dc8eb4635d2ef8d4dacccb7dd2c87de1faeed8df652d2d3515ea16f1d43313d4128f34ed5ff96335d333fa8850a1c17c65691535ac311265ef36465ac80774e07cc33de06ff85985e82f864b454533b1daec5c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb04e19bd47061833c789a262f705761c245d5da53ae6f2937729e365af29558bcd5ca168f6b017968d54e20b4e3ae82e1ba674ec3979fe4b8d0ee2e927366ec4bfeb117566f444d518946ae04e64ee282961fa2f5bbf995ec6cbeec976e45b62fac2fb422686af32765a181376fd4a5da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4baa87a5f008f70c59469c048183c93b840959f59db98d4902714a375333ea86c071eb4c1037f1655bee97a14216ed65674a87fbf2a08bee048ff6372feb2cdb831f481bd354add1d7ed423f28e7786157059c307632242735ad9656c88ad3266a39aed7c149f70e44df0d291c3d238d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21e5d12ce80d78b07cd77fac595b07c016835a2cb29de4191a90654f42194612c477a03bf90ba3da54e12c7e864fcb01e005e9ce546a6283448d673ffa17acf315a38d4642cd97303dfed2c8cf80e0d5887f7345b8fce8411c5f6630b9a63ba0d0f7770f9e9f079ee1297863d2d3ab5e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9a1df6ffd8217d5a98d53a8dc65b4644c1e84a920b641c48f9112427a8f6f72ccc84e1c4813c04e42a6f1db2524243809d2a0d5283f1f53c5a7d2a509b0aaf63d3d1f33d87bc1007078abae078ecf45c3f089205a6c66a3aa55face9ac9b9b4871cc837642898c4633da3105639ebe88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4aa4abed09f6bd1eafcf304d24a0f8b91d6ccb4c36d26c4847bc8473c17cbb8ad73b4622efb218c7f0082d9a124f3f77be3eed0ab9e9042bda76bf8ac56c7ac2ac75ec8b2eafe396e1ade1bb9773fdb025788e20ef252e812d82e0215e50acc4ab2180f2f1d7993fab9ae0ba1849ca1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f14e23415bedae6edf375153c8b6f58fc0035d245d669fb982d7ed51eabcf64796ed57942420ba4dcc765609ec12db783822f393f8e211dc46a9dcc54a0a0e52bbcf7db8cf5d0178a5c73c9eb8bcec451096510b8ebf67ca9bbeb877c50dd50eecb0d3ec811c0a5a0da2f63f990af738;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb446b8e02a1194edca16c817735f2225ddf73d1b8e363729245180d583677eb19ca646cc52a61ee8dbc5d3a7424995001453ffba4512364672460bd777a6cfa28ed8795a7ee4356915fdb81f027f974dd3d1205df953cfe0b19624709dc0a2e768541d6ea27f65d414c94a41ce3d7685;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb38b5005962f1237cbaf5911d1a6af9fe59d174db4e2f364eca445c1840d585c46cdc15b9a70999a47abc189d380d9bf2ad7c1caefa1895198ab0ae7f36f7e7f7b1e0643cc68674d0bac9d266dc0c4d8ba7af6e3b5a69841677b221f1343a65fe7835a14ab340c1b90203789ca092332;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he20525a9c3455421832c74253c0e1451564f7c148ea9fa6440f30410000ac74463bf896211934194bb66e0c24a4669e53c3934cae7ff4a015313250d1c048ef185e7c3055bba5b8bc46ff80fce69b738dcd64c0855315faaa5c443c0127378ca49657e04322efd7cc9266d984aa338021;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae0c1e8a187e3d4e353faf5463788086d54d3e781b22ea8e82108e88af0b0bb835bc9f55ab161a2e6e0e8f7e3e768ac98129c00a205eb16d1a3771f2ad9e837aa5730b451e1649f761bbcf93fe0983329b5f1ef2754a0a07050a6e5c820ea4a1a9fca9f8d7a3fb429de13c8877c15ac6b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf39389dbcbe0397be4a3d9afb5de8878f13bcdda2ac921c1eec138433940b8295fbb2b864c71aa79be87cf692400171176150ccf85f3f217f07246d757f46d64d2ad32c23b939094f2d4305004e739b5c31b7ec8eb6b7687d3d8849f7f8779a29ab717888ed9d95ae25d1a9a162a169f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h633002f515e603b39cae3ad85abf57f5e0ec2115992e2812e61e2a844ddeab0af29bdfdac0057e69dbe48888ac07c8e065296b07d886401acd12dc5b13febda7698e4ffd1215e74b13657e41a3bac3282f64653d7ac8159dfea11a25b1d23bede765c2f4cedc07db9084d92401fdd7267;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78665cb383ddad2693cc8b0767825110a3940d0dc7c8675f516a6b2984f13699020686c56fa984c82ee86a562ec73975ff5df2c292288b881eb839f04369923292f057f8745758fa75d72f0137eeade9461fcd3e15fb5e83aada83bd93289a21f2be84c1e80c28b7b017d5cee911db836;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e7d0522253fbe2871711313e6a9812b897a634e0e0e8ad167cbc82601cd3e6551007c869ee19b7d67edc0499fafcac2e8af60675a60e58843ba0385823effff19c0cba3bb3415dcd7cafd374b959974f95a125876058b3f969d86f617777a316081fb234bdda99ebef2c0e1787a86600;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3e0a45f3e0773eb33c0994f2a54a36425ed1c662399ebbb1669900043219cab479d926d58078cb178bcfb60e3444b3c4ef3d0aa13e367d02b650fe8b6b243047e92ec72e9314ec88587285c0e124957778000c6b52a839ccf3a5dd804df16e40a98ecb95457b325244a3c5d4ead32406;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67dba49b3a70d20db6e7022f79d5fcdca261df56996ac7fd8cf491ac4aecab50a05b9130aeee5997424faa3b960a3f03d251a76f04f426489b2d765d1235cdd5409bf9145f65836c9ea3d4a0efd73b3fcc5dce5752fa699d235e744ade9a4db183e655f272acb1aba24375da360c0f765;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10b70714fa4de54af46d62875d9f5e45c00cea2addf8b0e30a0a0f181028149fbcf4cdb4f3a0636ae7e02433b219344869fe5614426845520f549297820d83553b13257581fd183132a51b175dc110b127acd1b2c4a30c8f3ae77f3b41fcba5af379df7a7bb6a081454be4ed0fec3b0f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he927630d59bf06ef1b2067d255dc4d796a3c26eeebe9fcb54579b7e3b5b414af813c00e6279fdfddd9293ab31ba3892aa792ef1a450308a401b4bdd65031cea96d7bc0204e21affefb49f5d92f7638c3329522dab458a9de8eba6e8459d63f11167c87dd64d32763f33d3414469b18ca0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc62d9367bd80bc9ef7411df049c2864d8a24d404cc0565c473b436b3ffe27125b6cee7aef2f82eb59f4bcc8622a895005355cf00107b2bb5d1c422edc09d0a4d4f5056ab27c05d3cb3832fe785bdbe1eefea87b1796e858213dcb48c16c18766d56e282a2b0b07873196c36a72e981b9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h532b1722dbbc83796718411f83d83540c4903553be7fe2b9cef61aeb6b3585617f4d15e665d961043d3b2e5a0b125814814783e5de176c008029ec1f8460ba52a9d0feccd767d141520a2dd1bf1098ac04a6ec31573f85100b518e7430dab71c6ea2add19d1d066c187d4dbffaf40fac6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8af001a61ed8ccc0a902d045a04e2b407f68a5e950f714e4d728d0156720079daf305a91d5dd551b56dfe56d9b64412bf076c32033b879fb7949deb4efca52847d9100050cd7254a4c8412c886e7f46e8f61004032950b2f7a79a2f5c7df28c4dcb28eecb1dc8a176ade2ec5d99a7e2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae3a17b394b0c2cf42a61ea3cd41f63cfa608a040d4f6b7599b66849e59e7b961175da0392b03f34acb6441b796f2a462385e5208cd9cbdc9a5c10401ab23f1555fc9c6ba1529151b6cfb145de5e0fe340f35ad7c0d9a10432a701c630a3108b894e30929f3c97412c3147383706f9f95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he47a127a3e52cd46a9ae7464b01c88955a65ee7f57c06309017b96ab5662142ca72626e5d6f160647c0ceec14ae66af5f73a77250198b6d53b97619279ea009032c090ddf17590db07863a79d308ced5c8a78161a4894c30d029f57964b082295f27a0120e897bbcc65b044a635d387cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc76f09eca2c32f23a4b0fd16f3b200a43e3f916e43c29bcfcd4a4161855c48fced19df9357cbc85155f3e4cda0324b3f868a6aedd7bc38f9eaef7fbe86f03e82a8ce6a7fa3fdddb298432b8ad9714adf9ebde4abbfaaecc597fcd670c57de20b43125ca1bbdf09f679d125ff2df8057d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e5620da8572bd3b62071805787cbb181f89617f5ec4158281db03b1e76ac07ebab70bf42461b978f7c5544b8873d5ae09520c626b74872ce7a4779adcfa467b5e3f63450bea3e9bfc4e32fa44384930daf289867e83b64c7d3ae512aa0743e9a41b85d03af72d1201420e67cc348503;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb443f7d85c2eb3a95ea57a6e20d005b45f208c076fd655afc70f404a9bf546bce43cf4add954e15dad3236e488a2166a202bd535e279772c3c8043d4e153b9610b98bab6aadf07b1091fa2aa3d13404dad2a6b829c63f529ce3e9bea07a2da7e5374761ba2818c3b1294019770fd9565f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fcffee6c954044d95ef633fbface879dfaef3f8967bad3fb9e0a1fa5abf5356d47709c62df82f6d5b5d318975dbd8818f6a1c4f2b2d2ac09881bede963629177ca74a84b9ef63e93839e7c8e0928f14dfd0c26a3bdc2a9fa2fbec06acde521dd6c27293252e7e2f8490b6d6f07dfe5e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf36b99be900d53d3d332b3f2177a88fb31dd970fc005e698acee4bfc65e54e9933b9a3e2a33bfe718858a0072b0bb200a65c09e970e160a2250a24161c6df44e907a18aa93e829a7561145baa2458c0b7730064f0633749284db258540040da743c4ad1aecbebcb7e58555625e95140d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bc2aad9ed817bb14d8f5be29f4970fd45624c9377cf919713e822a91df55d1af9b8644b4704eae92996799b88f7ef1ed37df6c9295cf7bc07dfb899ffa07ab6c394d9a764480d64a2cbbdcf264a7e5a08da85e8d886692f6c442c768a1f3d221d0829de652f7cffeaa9fcbef84325c28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49e4f6769aa513aec3a5463abdb9d2b72e0bb4a78b5ee15c852c44bb748af63b175fd969aa61f17ac24ff35b7a061e762ebdc7a71d6f98f5909923d7dcb79fe35126cc2b3d30e5dccbef01e88ef22778f533dbb012fb9251621d79536a0fdfda6e47ca4cf2b93afaacda7f25e05ca964;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e9dc33879e95ad4d95050d5ab3610fc9e956a1915686afb977ce4eafdc2e1380d0a1135bf85c3316d6ec3b963fde53f63f1ef5cc537b0ba401ccbf646271c55354a85803e3ea464be20c6dfb1299ceaaa21ee6dca463201d02df21b19b4dfd4ed92638f75dd5f8d5d60ca149a2db90c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65ea595f3e72fc394ddc6369fa48a43ab4d01f772c30846a3851b2db7dc4857fcc4749c23cc6dfeaf11f36e58723c83b04625648385d6a455d9e628e2916686b2d00be2570cedf93a65f77561b417f1742b53d34acc73684ba4c147e6e588b2ae80e5fc5bbe882abe52ae34576d011b39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf15deb2e9f23a9174bdc5b2e8e529686daf075acbae4399a28290ac43f4e0b6a2abeea88a1ce92646674039627ce2422edeabc2d2025b3d7114e998855e84a8a3d05840f99c344b130baf351dc001464518d435eaafe573f71ed8ad947631322f8fd36900f8c748a90f77208ac661857f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haff47a579d4850a384e4cb9479c800727df82a845a3782a9b44d9e7f43fc96118f3d6f9a4cb1434925e3641a1b4b4b32682df634d8f5c8dcbd35a51e72d38d2f50934cf1a116bf2b2cb365664ea3d8988e32c78f2110aff67279cecfe06bd6aa446f88938cd77a99f2aae525d3b728a86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d734c57f829db28183c0abd5e980b6804bf7eb406fe39e79ea5a2c29812c61421538be1b992283f79944a3e1aba9df4134642cdf9465f6f786ad9f11dda1e6c626878b9ebdb7d43d34b5836f036185d263cbca7c67738a2826765dd05d991b1c9e64735d07ef467ee0b64776a16ff743;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7067570115ef7beaafb31f193d88b19bfb65cbabed390a479324b603bf8a32f0b908ee9bc5a21e883abfb86d337dbd2655a2eb7b63a646113ee6e21a0cae8e1bd31c6da2f18175ed5ea97c7970acf800507c59cdbac76ad7d17ac1a1ce0ddb9e172d824c52a8deb866ad2efbbf9c278c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2624b817c38c823bf222776a89a10ebb3260591ee7e90c0001a38472ebee7c0cb90b8c81d5ccb53222ee85bd0965eb287f4ef16962d8c7e044f677796d25c11b5119be00cee14e48ff4fb70e119d2da11e0df40d487bb6a3dad07670416b3cc4234121578eabfbcba678c264c01e9b4fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac5b7848895c0d51baf556698585537165aeeaa65c7a78b464615436d8643fdc6cbdfddce606596244d1f0c8a4256437ee778e00196718af38eba18412d91a9f57781f4a351f3df05581676f7d8a2be18ba02771dd5cf05180d8f68ff659b724d4e07fbfc87ba6b05694ac7279b9b8d47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50870cb6770c7fbec91575e3d599e6769f335c21c0973592dae740700eb94d28959420623ad004cda72c13d074e6ec84fc4c6022d9e27d5c38d22e7c466df1ebf2f764f7ebfbbfae87843997f1a8a36748f700b8f17be49568b5556b156e34b88783ed40a22b7c118a92e2312b1b3cab4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3b26dcc8f8995efe51ef01ebb1e77c25ab2ebb7f57017035360c8d2b27975fee1fd88bc91d027b38b2c09602a3e0fccf5e75b6d73398c650ea28e2cf64c91b9e92df50f27d89e61f01651230e4e73fc91386cc32ae3a248afb9be9ce764937fdbcc650510faa37a531c8dbbf66a3a821;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c672f658953f46bd2d7a95095077f1d422ad3f7e0db541835f74a5fd431ad867763f22b1c160e4d4e6b9c1d4c312ca47a80235ea99dcdf9126d2e1098b479421663f222929a76884ceabf0a859104ffa780cbf84a57e45b2c9b79e89a08caa45330e27c03830b74e7a9f16c0520a7a33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78d4691d3fce77a36c9c93cc9168d6801ea0a56c2851246d9ca319ee11a3446e2e7cd4f52d239bcb60ba74ef7f8542b73c73e15ae0ad484b955efcf5fed58892ad20e9a1ca2ac41b931d556d26a1dc8c3f1eb12ae186446bd2104d1bd2a8d5061e80901bbfef89d3cf03dd76d0fe235a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13b7d32194359aeff406aad466a3a49c0b23010c296815908bf4dc67690143069343d36fcb849ccc3db75cf22a04341faefb49ef1799b62714e1401591c48acd2cd68c058ef333219d2adb41d5a350f9c5651dec89bbb8cbb0fd2b272c867ce45d2d94a56aa3c97fdbce415326c264df2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbe068a4c6bf0039871f4e42af31e092843c2e28d7b44244194d1a29e8e75222cddc3df09e75d26d6b45cb8a5933650b7c2dcfb9fff941b8697ad07c8ebc246a517df4c6c9a2661f3ca6d2ef48f57afadd3e6d9d8e0947e4f974bcb81c04395a513bc241d1b3ec25292c2a8f0f3518d32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eb5c477d118ea573baf1eef0f7d9e386e496a4cfe065a84ec2095fd18a4d467940f28a6f481ef540d63b22dc0a0985e3352d57b76660f9f2925006bab2a213b00cce257972c4e4422dd719a6a2d076aadc523d6c32aa756e4b46c73ce513fbfb0858e3306f36b05571da0f3d9a89b1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff42f48d0f065700f44620a14493fbf8a53dc298ca2da15b48c869e1704293fbaac87306acb389522b332b8862db46c968e4e06887bf92f3b603eff8315dbde108d02f33e3d7a9b7bf6bf65b611aa8d959ee1236e8029926eb8587b655f4d1d127dc9a1909f1c5d3fffb12b98b6eb5302;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1756dc64bcff281229b8886c5d345a04c67208b710fca7311a5167ca84f891e4fdfaed4cefb16260364a0466c122589a610a7c8ddf54fa4035a3123b8221fc0e00446005e71acb6a2a55a343ac60f0ae580eaa6a8d013c443dcbe0f7e58ecc3d14d50a948478e92723c560c3db63c5c16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3ed7e97087a6950422980b2d28af5ff11d51b9342d53ebaf9e9acc1d38a403542b3404e392000cbe6192aba9782e276302278aa0a8c012de61933fb4ba05c7103655be62e2fe3970e625b6c4325d742bdd061cc0e956bffb9862bca46789f19a34f2e403b1a4ef966ff505f8b8d4785b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c9b988345affce657a33fb05faa9ddd8831dee8f84d597f4dc2d791de27fef323e428eb6657043c92bf39cac92d1c21cea1bc827f1001cce1d934bafb1dc122d4596cab504474ed8d487cfc4cb8c3e845e3447ab759f770bded110593b5406c94f89bcfa813f7ea2a4d3c611c7d6b48c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28f4e282d6a103dbc3a4d9b65cb04f97ccb776f85dde70041b2c433e0f932bc9deb761b6a1ef52daafec4e06cb035659fed6064d57b4f3d9d1780fbb13e67a8731b329786434b1cbd093c71fd9034f3be826390f04b775f59169ca04cdae83b7a65f21e02a10da0b1b897a1a8a2a71431;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea856b6e33f5325a3a34822fcd52e2c04ec583dc7449ef93cbd4e356a8d06699eaa414205ddfaafeab5f0b255a00a6e1cfe07924aaca69478768f3a94000a34e0c8599beb52c2e3f2acc88c2e5bc1d86f50a3af0378f0506ef6fe86510898b0474b0c84059d6043757a9ecf923e2565c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf116e5a9359c49e93476067e13bce820a37cd58f29c071800e39060e08ca3bd55065b1b03b37ae86baca3bb9d7ad8fcd80624c880f8423ced038563595722252d868f4946fb161ef1ddb45b1bb749966e86c47d89ce9302161f25f9cb8f76721adb713422407b3661f9a61be05bf722c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb46793afc0f425549f6fcbaf6c8fc0f13297d0387e747d15bb74cdd02fc5584ec225f759cd9d3d65a547ee16339365b8723bcf0ec265f5a051b21f42ad253c0e05bfb268347dfa3bcc3960a7b3e4f1de88f90fe50daa97b4d82ff1fa365851ba181ccdacdbc5ace3c86354928eb8cb306;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc72062596ba4f66b39e07377cacf205469a0050865ff80999edd77a385066e8c752833701b1b6311543efb442d5c1a218c5a54cf8cef62fb6d1fa478e5a256d99ba7eae0a036b4cf08c4965b5b0405eb7004d4a07b257fb883fb0843cc3924586026bc050d8a5ce97f5622909b901f164;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b8e245ddda8eb68acb454096b486b63e5c87e941217409c99ae922945ded8ab3a05decc21dd82e1e32df46153bcaca4a7910cf70b75cb3a92238a14c0a68414e77ca0545e62388cdd1b67f440d1d0d85f5d275246ab336fb7cd74dd66e30d6a876bc3d69aec23f489ce22d677759ed51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2512325e78451dde1fdb64fc52f1e9469ae50c7e7e8d53e770446c586dcbe778a1a2781d7498e46e66ec528f15b722acc43dc29afb918c97a3d1bc5398fe84510fca5c25b4c2cbb6f1da3b0a1a4e3a3fcce361b8c0ffd81e948f23a450ad6a50b2777b84c2362a2701498b37eb8fc4940;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h487cb081f4b0c1ad44539e957cba8e92d5398bdf8769e8f947e1ece6d442554f4cb15bd90ecea84a638572bc575a9f53d64e51df16cd406a37dd4b66052fc75930ee4f063ef44db2defc6a9d9a35efd5f5ecebdcbbe8e0d0fbd552db0367c02d79ba3b02f8a039dffae0fe88b23eaa6a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdef34fa27a668690e72a8eeea9237b81049144a0bc6676fcc6d99c815ce6e8512243cad99e6211d4a550f9ffb8baea087291fd7c3b3f65d35dd63dc8d5aee7bc6c4dfe197f17bb253df555e8e14a05b8f2398beb0b803cfa7ba350acf5c679cd63a350cb5b0e0a7106c4efd25875cc3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97b0136e2e01456b20ca0de4b3e282e803aa9ddb943ddd249a80ebaf02caad411207c091c4b3786901d4893a14c120a7335422bb7c5d3aee04b3f96cf4f5e11518468aeeae14e60655aa91fe722796c33b275e9c2ae4aac567000d5e2d1856593e968c0a285deccdd7513ade191ad539f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5630fede841a3a4ba6442c3f0187b5fe12e17fe489c44f88182041d1868cbb0b0b41c96c6990c2d0a9b3bb34b39244c8c2ab2cf2ca8263827eb0021c8e597e2511532c76aa882a8a474164446e34a46473d5ee9e9b75b1fae9e77a5f0f7fbf5ae235ba0fb73dfe97c4960c1a1f8116ece;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd58011faee343788ecc72e51825aeff8bf3f552446c8d15d7e50a2428eeb6d13fb0a6fddbaf412167433d098a70ce3520177a13ec43f825e7a07f40d1a0721128fd87da92f46c8b57a3f498529df7ac0569016505ca3ab696527583befc99715404d9fcb4290caa5aece6c2c182c8d347;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbba11dce93eeee3234c78dbc065a37386fc47d10d17df187e3e12b5910008963606547a940244e97fd8a3d33275311e845c95bac95125615e904f9c38fe6b16166d2b49ff79d9917f2d136d922685d26a4905ecdf026010ca7d4c94a5ab12b21ca2278be7806a7b065c2f9c28b8e3a55b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ff0547299c45f45059e020a62cf5976516048d3065b159e584d8d52f34232e6a96ef8c343671c27bdec062f761a2fdc751ead3f9dcd488e83dd6e45ab2ca726c943d95c019fe37c457b2d04431d942b66fcfe6b5182471b22da0a1209a23a7cfd3c6ea0ff2a13ced68c82008c230fdaa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95bf5dbe2ae8a0d80865d72e803cdeec9c54d39997665340ab45853fe02e06908dad9a26733411c7f3f8b5a31968e26f4f65e5c09221199177893d4ab160e6d686a2396a0755ba08dfe1b8f8e8901cb8f255885663004d037fc92b976814d2c92f62d30d451290bdecb8200ee4aa2522c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb749c283a34a6cf76feab7debe0aec9d95eef159223351fb9f32f4a923f49d6c0493dec5ba8fe776a7faba28cef82a85ed9dfa7c088f5dd41221b6e9708664fc53a8121a1d0799a93d9ef8a2d829437337991beb6b0594f5f1a8b46f1757c2c21257876b69f8b6c0ea86a9a3b1ae4f264;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a603ad75991182d956ffae860be725efa575627a8b50a476117c10302401c7373b9e5fa74f3718905ad03cced7868e8bd8fc92c2efc6ba5a3d122ad11d9b44b7edc9a96959bb0bc892e52125324ed6e2a044ece831537207b17153247d3cfc01063d64c6097511ed0bcb7e8ff87ef257;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha73b73718f880501bbc81a7d57e620532003442c7d70d77a7f8841f4b87874596f1fb807298ffe36f9549a364b8895689a75e5688ada9f6e54075f42a29359b4fbf75e50e6a89e873329d12abe4d07acbf70b4d32909682d0e4ff01803a31ad433c2f9947e6f29567d3ad62912f72a20e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h645ea2d1b982b859f62714192a02c935487be5f5ee79114d289780ed63e77a4088f126cfc35c7ee04d8a45cf4ac9e93f3dc5324ca96d84d2a8fc90988a1f090f896654628e849e4c7cdd134de585f67843e7fdd0ec8f33d684cc6ff23f3134dfc9bc647a52cd57ae70e2a7abcdd7c63dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f3b863bc5fef74860df29ca171f634fb0df3fe049f52e1088a05293ff099f002e38a8f99fa0a118f03e301ecdeaa47ee0823dda25362bfc20c6c900da86e155eefe80795d810165fdbfc3ba3888ef5b8b7d6a0a07f77f58c19925dd88552ac41bab02ce3b7e95f0e886478e7ac28fb84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73fd75794c5f8af731d87ba356302d187415a6ab061eb32381b3aaf6e14849a95f5494a8311230aebaafbad0799c792d77ffad56022a7ef17edd6c4fdc72730e77c30dc6fca1ac60cf91e69393565265c4fb164306d9fdb209ed9e822721988af3641cecdc48710f19a89a93a0fb9a405;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3cc2c8af8447de7c9c056f78a0b6ef80cde7119fe51d9ab92701f293d4466e25a89fd689caa007b08be859b3e855211def88520b4c2b4782b01db7b033cbc5186f33a1206c73e779f486498887185a193220c7fe59b35f01fbc5cad0cb3dd4e55570c825c25e4a9874c4bc6fe3639b97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e0dc039effcf6644585dd741ac0f62e7c73fd257ce13efafe7373df5dddf593711e8996e3291f7785e12cb26ac23f8223ca9710e6b1f7c06a09c1a3c0ad03d4b7102dc192e5ef27af3ea46aafb325e5907ee8e1df3af8ec95bbf6a13dafd62317d3bed907430b906062d7e5a6dd8d615;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a84eed987cd2a53f90115781131623127ea3be853a105c3c433d367cc620ce071768e18f6f3c35a1c2b87a9abd8c596ededf6278344b2c4a8f47808eb4587ee0191cf189b8ca139ca369906bd410d14024123978d1c2d07f3858d17a270607561f17716b27affeebafb593a970a5c36c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacecdb713d2d4f2161190398488a06493816a64da0c48cf3821354f69949ec3cd22f185e857ba17a59dca5986aed4d3babb8bfe5a9fa2e55de997c260cbef01207576b1c4084281df5754d924d9db8abdfda7410aa949d8d914bbd759ff2124d4b179e2869cc017db229cb33a682a864d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59375c86a363c8e7c3de8b579fb0017a298d3b28ef12cd5062b262abc3159e30557d46c28ce2a59f93634744198bd62c62e29174b304cf26c4e007cd4b2a97f92361814763690f433dbadfac7c367f89cc5fbbbc5ba96194f8b7425272d2dfc53abbad1908aa588fcb97a84811842008a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h824d905631a31fe1b732e4a09d3e833dadeda78068f004138c8bb0c5d648bdad65fa01a9565a88dd4616998e84f880d8f865a3ce5d212c9ef443c90bf873aedf8a220d1e8a12cad8f40d1de4827a569eff72e55f9ebc430522966ed3f9874a9b09755c337d544bfc67e9089d20f31f110;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ac18fcf5a83fe34877e7e83f6f541368d8e2732a6a61af3e6106ea2861b04437db6729ae0c77dabefd3ab16a2562a87ad898a243f41c7a36a9817fab33bea11a39dc3626b4da4100263c55db297df0e47ded42f8b0ccb1894ae7e338000bccefd174c62b53275ad117f82bb94399f3ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3c563bb6e09504c8960520456ef4c7fb5a00224f906a05e2e79a507da6aa79ea95aaa83b8654c10c1872d4aa34c069c277a73eea7756062797b35f7580af563b7f7cf3f74dc157cdc31dd2d333ef5e147ef17178bd862b242d95418bb9ba83533a62cdeeece86d1b0e45b6124f2a85a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ac4b24bd6bcfcb87706f33d896bbff7fcfc25091a4fb9e9e4f87d61c9db502c4ba7a23331c41657d01233d4ddeeb2534371281001c3cf6a6000e983530ecce41b4f79e120da0c50b3c0661a762e5fdeddbf215e107c1e264315f214b4b33030c581060e5f765d15d597217e76d6e96c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78d9c2a9c69ba8558f4a2449359700fbc97318d20b026da71905df6f7e45ec87b2ba055d61849741d5a6437d10e6ec0535ce2e8afe9f3ae3ec3af34055306ace271ccff9dcd38bf91b91a6b7af6819f7bb21e2bdd2700fc657b6f7d55ffabdbddd78ea46f1963917f98eb0a2bcb431a1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h986cfbfac0a9f2a3ec5329b75e535df15d68ea829fcbe13e460776c6f0e96417fd1a11db1ef1d304a7f165a15e4c49673da8d5ea4f66b74d139f726b5b184bfeef898e1db23547535fb3c305e5e62bcbb6390eb554f7bc32671947a02f512e5b1920b2cb5369739b478b4e9bb7c38c066;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf770292472f0cf21ece6aa760f51336cf802e5ffeccbae85e5fda912b2cf077a281d4ba1c076d3292c199fbbbdcf2cea130139abc4b6355c2a955f7202abe1623100f03a2c67a057f1586174e54f43671eb413f929cabedd7b346d5f9791975023c0e336460ffa96193e23237923b76c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd40629f77dc7d57e3def32ae41cda847af982ca20d2d6cd46dd27764198e8c52181a8c7bb359c80c23dec1c305125258037032a4fabc1d8bb3e00a774be81239a87302ccb4ec838d192ae8a4594ea42c378d2d395fdad86506a6942a070c70bb824b14f2f599bd4dab0b54d2997b24151;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a98852cd79f776c1719937b652df76ebfa3cadf6db1a3462ac1b20173fb5c323a51c318961516eaa5e6a7d34678741d7712c12976a83b7401f24721bd8a90f68f0ac1ccd9e70c976b172ab043945cd22433b8fb747423c9f8c8854ef523a9b84175004c19b244d52a0c3905ab54e04a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7816d92f4588c3aa98658dd3905bcc34257915b5ce6a0652adef303bec0a00727aced1ef5f49a2eb0614e5121195841aa83a71e3187a0eb46c54059dee858c8086e1bcaf906cb2dad4131c69cd1e22067f8816ebdc8aaaec2c7872258260b0ddb62ad99c01389acf506c25efb06d6e203;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f9ee72b5a4e7a67aedd645685834fbacb4776d1a5a52d9a608198f07e3216f6ff87b187f0c354ae26edc74f4611239654ca747a33e8fc7d91d48e657b7b236be4cd7018a5baf1bec1fbfb60299d427edf9cfc0b4bc0862081ff8eb6d93147e4e6839e2fc5bca71f96e05c5b19fc5b600;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2dd1d4c09824e5677b6a58fc3d364ecf40e790208e460b02af37bba633636d149b6ab223fcc358a0b8a4a91c4ec8146741985390585277d8ba30eb24ceb86366c995f52a37fccdf87c9e001413978e51da09ac951912fa7543c27a85032b5f00be05349f171d36fd4ea9d219ecce4e3c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d1c1a0c74409c9011c81a7045287ff0707f2d85bf8fce96e4c406cb1ef9d2163dc1569dfa1fb5d18adfb9e8e2a8f3df156556dd284d946ce24fde100db16488e77a4cf76cb9d875cb52deefb3572d69275395c0374a7586baa5d1c65ecc2cad26703a9ceb920e58e9a6477291b6db359;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc20e8b66aa90df2dec4180e472550ec2dbe75d466ad1ebbb80f69d6f38b9a2c17e16195fe9562eb5b152dbcd120a82e4028d5b1c241eb206f8ea5b8fc3889879bae45de700037221c3868738a729c3685c3360a2ad7b9ca51462303f7cdc9c32be758f40e73b83d232044f72f76cf540;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc188ab7600370458bafdefc24810c7c469913f477c7eec4496e2a343ebb5a0ca9e67bfde0f5ac91d5dab375ec944f45ae0c0287084254d8814ab5e83e57f35511ab192b2b86a2aa2b72045ec0e91b23de91d7d9c1d4b008bb304765201053a4ce58396f21e32e15bf4f32f7611aa0678e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e04d9eb563809de003aba31386dfa7e4e726b34f4beeefb08f677af5c10d9c8f9077f14dc19a7ea3f0db6cf3caf71fa95d5f561ef606082744b00caa1d46c2831063054c24ae6ba6f1c84a71e88177d20232e5011c8f183248cdc2a5621bff2231985f137d98dd4265271fba88e80602;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e0bae69ed851890356cb4c75df2904aefe8ecef57511a3a7378d2c2a4d3482b5543a1d6495de2e73c5a944d74b3b3620dd4a8c9757e99fc8ef9ce777688eb93744bb55022df5a42590f2ea9e658821f940a9f1949100bf9a7358b40d39c3778cba2e78bbfd88ed1a3f27a8468971be87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h435c49e8a7c5e74f5115842936dc559cfcc002d41b9204864b73611da03104064e621ddbacd10b29d89e4bda86872295e3541b8b83a7b14b0aea76dd487c532de318dd0642f528d72be608c6d1b808b5d6ecae61d56c97b5f84980e956b1bfe437cc305bab2b25ee8dd07bbd77bfc6e93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f6e2e4002b420c8a3e386d6a00c118909ec745ea70d08eda2b4d1618463a161317edb83266d3606614eed0215c0f4cd563dd2225596a08220853b3a9c2a90199b25600f98b152ee2b7e6b34b466704aa459a11be385da0dfc1c724cf8575bc7367e1d7aaf125852f1860a22e97ccd08;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90e34cc348789a6c767829cc3b3867528a46d8ac5f7b517ccb9fa5108ae298eef93803355c1268434f6f9709ea3ba8a11d003014f4210d5f57987f49eed37b86f7684faf523a4a5d1cc57f7651163d273e20686d6b1b4ec45904a1f6121f35bbcec60d6efc34f89b30caa790de489206c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc061882c22c4dab18000d0beff1b0e473e0e131b9995f7d2ba7ba11e4e8c7819f70596213ec87b490b93b39c8ef03172bc4f8c6e9b23a6bf2e80ae685569e2c189eac0833b4d18f8adc1f424eccac50966469a128c2ee1db45a2579870c91392c7742832ddb9408fa5018469b1be3889a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3d28f72c22029ad114812840c122ddafa085dbc3af21711d475c7e9a16d3b150399feb204ea90d9a4148aff946ed39cfbd0e2b3bc6c76fc29c4dd9aeacae8d943af43f8da87b5643ec75b12c8de6804f849b3a10b122eb187ac2c7746a05aeb72d6eceac639d3c2aeb096acc12c638f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e29a9bcac07dd53723e93aacf6a809416aa5e0ec07daa3c486f4b1d28d0ae19709d14ec041dd6b6693bc843881944e2a11445c97a9d8af0d2f83569ae8604c17a2cd823dacf753c4d861b93c23384cc17e94f09a6d145f5a3ddb26b79022d1467e5b9595b1d7b2ca9c6abc442ce859a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8284b894ad53078139c91a5e4e5400407282b3a8bc99e9510708885352e758bfbeb942b06917def079c17ec245e0bde5d2c66520b484839d856b795974c5d37bd2f98c0df3d9dbd7931e10574f089f726c22b1edeabb066032e3165b0341e8e4889754d7e3ff36d34a66191c762b260b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd01bf77dc15fc66a0af1cbcd36b5c4460a04b4c0d4ebf7b7004bc9749d8ecf1d2ff41b9e9f1962f0f0f2dc92c11a206c5391b4a3c36d7526b1f55ac60093a41218902067098ceac3f4a29949d16e30909140b710a0df9936a2dfef85b4fc0a3f1b135426401e08c69288e1372f97feb26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bc6f2434f2c8a9cafd5a5c52f91d0ca7ea81a3b1372cbf14894e21c537994c148795c8df47104ed6b99df5a63197be99819605084109c92c74ccc8b6bc60446072126115a27129120486c1c0eb2767bd93eac09dc575e11b3aeb5f9fb1e8b3bec5a2a3f173176760341a97f0c49b7e83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd614a4c718c662b49aa912617810ba529ed1212444d43e3bdb7decec04a80470e956fa5623c516882d574af3e013bfcd48dbecd3866ec7ffd77bc85c01e528351b0e848dfbd0265aff53cc7fd60d4d00595ed0618cb3b7e3540ab43e3fda0708cd6d066768da58f5a2f789d407efefa24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb094569aefcc150227099f684737224a0f089171f4a72dc41e7824b38a7c0d150194ab180705ce98cada8a1d97df2352da62cc6d595c50588dbbb4d1802d7b35ece49efeaa6b2e792425669bf9ae61283b5ce30ce27512eaa2cb67f85a067910f02a9e4965eb9df72ac60db947f0b06b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7303d370510c12eb45b5ef29054b8b9c4d4fd380d4c435ae40ff10779599c341725ef5168d8105f5fa2cb4701c306613b557e17c1f819139cf4551aa48f66469b24b9fe17731ae4098248e24f5f99f94bcfd3bdfcfdcb5c4442ebb33d6db4bce5929d2e22d349b875e2035bbe50fe1dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h852f00263bf8ec85c3357fdb337f300ae8473d82e440201bd30a3f1f547ce06f401a063f8016edd5e912566ab05e607f5925ffc40c60746afcf9034a8db6c208e4b5d16b8a7b3950542b81390960656660f542631df7c7d4ff415382229688a75ace62221aaf890119870375f816d1725;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30c3f7a9abab12219320c0fb81396243d6018f5ea130d788df2e6fbfcf9a87e74eeafd1de20a539ff0e7fe4616db64294c7accd81b3911d177b76c4fc63feb7aa517563a6356d298ec40ba826ea133e62c66914b792c8e4343b5ff6efd1af9242505a7a0f5ccda2e77a08856a5cf22fa5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb115b6a6258d63317e30f88f7fc95156b5cc2d37cb7a3782490a71815e687e6c30cca2d6851dd747080dba7778a8568122b7131746c7287fb3bfd982d824832a1065e8e17386d1b0cd7464284c756497cb03740ea44d84adb5028ef01a4910da59685b3f9466a9a400f26891c0d2701f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bf6337510ddc03ac1cae73efd4cd687b8cf0137ba92102f5a33cf0060eaaad17afdd8dd25fc776bc7865bcca134bdd2ae1b941ce477c4e571cf6a39149ef76cd1c518415a21039cbae02e42b85d71d35af9a127349ca14acb4b019784ad9ae9e386d741c8f8bee114923120c75e4709e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h933fffa7cdf0e0f29760d9873073e7d505d3178bf9c27bbcea81b77bd1d11ee61b42ac5833da38e1ac79abe0f1df24da0fd1750aa15b3f0008d5a6ce1c233328b553940ad7a90e25a3f67c6d547258e85e6c9d4d5d466183d117fb44cca12618bf78effa8b3f584c9a639077802f06d92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea7d6c9c4b3aeb39453da38c3002041eed5a3e8e4bda4700fb7ad6aad61583787ec6ada10af682d9de45008569941c0cebe721f7997c6f45fd9679918275419322daae3f5370fff23164016f8e696744b7fc1c4435c4a325a5b9cdccfae9f5ddf7e184a55733b1019c9b0fafc7c0e5986;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc51c004fc42c47d14199c02c3a3da0328ed31fb79385509a61cabb4ce918b9834e79b88f692a1a333413bba5a1839fc7d98358171f671db8a6a206739246ebc425a3c1f9faf316f74f54636ec0ea2497f807c0df770f562dd6940258243c6ee6710531c700522a2c73d327f53e07f2256;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed33c39e75d3abc91916c8fc668ec0647de5be450c7e9c3639abd38aa81161dbd3e466a5687950d65bb7983d6d6cc12152e578003ad7efcaff38dfc0d58de7aebc931ab2b9ae6658618e4b441a7af15d4a7ca72120c29cf4072229dc9dc7c0572f4f08af47e20fc08523ce2063da59d79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h244680681f73939bceab1319b81671184b0d7e0104b694771348678734f08d6c8ef4b307658c181236ed2c6e2bd167ca9172f003d76029cd0d3d71f3136183a0a95f1753fb679e0815e465b62e2b6d7d26641d28f71914df4354fb3a90f3006e61a50a8ffce266e1c6dcccf1f0933cb3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h177378ee8266cab34f2ab4122fa491f2461575aa2e1c8d6b30a88728fab9e1dd8dbf264023a519d1e14979e00fe02803ae06267f513c3cc3a831f30c924940cb05c2d3c80ed3378ca7bb5eabdf4f018cb2e925e0e27a2a1438286b747b6e002a9746b5b43f2afe04d5aad031f9a1e7a3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf06d381b0a4f9e6a5b42a0c9f15e52784e999fd3e9338be0db546dc9ee76b3e05e23bb8360efabdbdf31596862b5c9a9ca3ad657d409ed8d94d69c568eb7c62ef40734e46437d303bb0164223ff110b64c27c8b3ff09e4168d92bb193e4b53f6a39d9b08cdb396cc4b4a38f701a724c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12cfe768cfc1d1ae38be0ac9c4e9ae01147c9930f938aaccbcc00450e022e434acdcd8b31c450b26a68a41c2e3d01b2dfb5b16c72d55e37199bb1ef3c4c954d2bad8ea61f65b27afb0364518b0a717da7997fa94cf008935c4731dd18eb2eb6ee5e743c64227a0c4ae4ff7a763ce4c02f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b891be639f5e795d50f88f59dc65b61e8f7bffe0b7d02a68a8eabf63fdd6a98d460b7ff5e2f20a4465ec40c6c3ca7cecc01f4e4566f383373787777de3c1cb56355c43f46e7af1c902b33c5468a85cbc92c5d1be711d50c241c7206ab2d29b9f1c603707530cb77e0a9e70c6ce9362f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b7edfbbb497039193afc297f3b1a001f25670cdf798efc34e2986e4130f33e8edeae1e6a6d78ddf30eb8d2d96a24f40fd3c68e3979ffc0fab4b538a3d25b445ec1631fb865fc00ad0c73bbfc01609b660cb60f7a137707c02f1fdcfd36c42f9cd5f918993518923482d491f79540cafc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20cd6d725b70a0ccfbbd59f35178f25be481256d2351fe91390d38b017de368af8b63fd7f0a81286779fdf649f8c19fa5b96ce7bf53dca22940fde2279bf5775c476ae7040c3d7b1bda450336ca00efb55be322d14d633b1a019665ffe0e0b0ad4217c240523786d5561e7808006fe8ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4dde7c0bfb3421e2a4cd80abea250aaa11f36ba9eb45b3e6c1c6ba2dddce875e7d71a9d8e6b49b176cf687437c750f185325663367101207e2d9cb5c7400e2bf1259cee52943db29cf08038185cc0a8dbc1455270f0f1b779057a01526631035f75d3ad06d6eddf1f9bef85508f8ee7a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf66cefbf5e4fdd3eb4640776da9928a72b01567e656d6727a21d2a9c0d924a465b8b9ebdaf43d59afe877f5adb95c45eb1ce50bead09d26880dc86afe9624e4f96390c6e31a0c317c185105ec5cd7fd3e9c2c6cfa8539a22b3d886994c72c98e4f014663dc84e03791411ecbf69a1f14c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f95123dafc7b9797aabf32ada1b3f3aa073482aa19629c0555b098302cb30609db8053813310aae47f3aacbc153ecd2cd3097ab06710ddac17f6a952998bb8682a30cb1a1d1413cc061f3593649c56389672a1a8cc22956ab6afc6fbb4498bcb001970d1be0d9416e2add034f3c4e06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0437d84f5bc43db11732d74cd279a3d48145e5d7c009f089a6df1f300a5c27d5a815bac948afbdab5629b18468a681bdf2b089d60990e6da7c7263c8b13ec418d7b2076c227d436a2297d2f869a9d7ead016dacbebc45736b71efa0fa94885b11f2655dda660c04f46e11de819dd8ee2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha98d4a69a3c8fec6c5904531eea16f29492ad140fa26b55b0a4fbe70248b9d60111a08af18ce888dc0707452953adf3e6feedc930e529bf9ceb8462344c95390d685b4bfb714911c07f124dd45e31be209c487d315f021f51b4b808f4b0068f8676e5ae09c8a04330bc80b96f7ae3044e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf170b1dc7a6109d4b26e61b050ae4a5e48407854d63747b92db4d777fc45aa2b24cd5b32cb7e546258cde54802b6d97c64ddd631adf6eb8f9a0a101144cd5e59e48dfd3aaec42d9d7ba71c2a7a9281cc8cf347b9b8987b6ddf7273c5b6892bde84ca20b04a22d494b1c7b82c5b95fc122;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb82b93f937a7943458ed376a3d91c91d371699d89c374e6539ea675502317e7206b2e2e564df19b06559d9ddd84e8b2505316085417484d21e3a786370c5f86f0a7e29bd9470fb5f1d45002a61e62630868d0111f1b7188632cb7a48f0d4f45fe236256cd8803cbe4913253196b555cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b673f8bf40ae8cc42da32de02918b556bd9416eacdc32409d7b490d6699df829a78e22466fb2b4cb64b8e821c85b59e5092ea0635d9f4f2aebf965459d67bc611e59fbe53a70838948e11be89076a7db194f409b98a1d3219869efced83569170364b20b858451ec03bf1b75845da4ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a059a5a8f025c575451cbdb198f491eb1a5d39d0b6e8f4e793403c7be8140c4b31023c17843edcdf8f9e2c5fabaada1d42c1e89a262152dbb3a094b47a8f9607087c4307df20638896d360493b30918709e38ce1f873327012023809125554335b64fe2557d79aa5caf67cf57d54b275;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb73f76c9cfbba51417097de4c91c728e07004f2f8b66d18a66bd6cd45672617e0d500d4884cd87027ce839baf25cca0110d29334d9be2e7baf70bdaeef5e51567899488080abb5419a9d661418c6bda7db208d4297664687a3c490bad870f5e5c30b26315dee8d6ae25b66c4245e94e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb32eb391edad509f2796b67c0f02b202f43072ff2c1242b9616790305d595a378de5413cc3770e89acde6a814befab33e7e312e6616355c0fe6387b7de6c759bee444bf3457af19399a5403aae6c95c723ff7700dad3b409d30eb7b973cffef8631dfe6358c001d816cbae35466734cac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b3b01968e99d63ddeea5f47739c17a1a840a0b3637f14ebc0a1d2006a3a36ca578ef923d8aa360563dda631158741ad9e57eae8b1e37ea4720fec3a33ea5159105197aefa4524cfa5218388a614dfd956b2389dd72c7c48b57739fb8a30c14ffcc24324bd46a257219ff917d6573fc9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9feff5c4624d8ae79b6a316130e3ec9725b65f367646d31477cede18c52e67e40da946a08c3139f410d227ee9afb1fcbf45bcd11da23cf2dec6d8c56aa4c4204d872af1b8257373a171978d7896668d64e81df711a495bd3087d7ade0a94dad0ee70fcf00fafa28e3008d68b05cf37d81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3262d174c1245934d9661a0ff029e37b4e3d9ad2b21267090eb8fe002b3b66d391357841d5fe0ef5a7591299c3d65b9f987a8c3d33d1ef3b96037126faf7a9c6b3759c9542d4bcf9a1e1a6ca12bf622cd4775b31eb3daa077f90d30e2873885169b6fdf167551d7f58c68d1d9e09f557a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54d0a0806f275f9f631b737fde30b30e962d39ac2a39fc249f44c37d7672d9580433091da5565c0fc97e36e7fb8aeb18f2632500e9fa9cd9fd1db7c1ae820748752a4f07221e0c3e3819423497141d7b655e426c452d5572d94178e9abd1488d14437fe3aca160f944651ab9fe46ae710;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h588bb352c2981f81a8e55469f87ac26f9710ff1127bc3e5f60cc66fcc0f438293aca158c0baea86c441d5c422da5e436c303c66be7cead49fbd72bfdafd9873586a958a64953dd7ca9b6b5b56503e60d71414139647d5177db0f5c800ee3c817e4957015772bcf49a3e45c58db6a5c556;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57b019ab67d0cbf9442e165b6068ae95a2a5904fcfde37424fa19adbb24fd93127c8407487b5d1166596c35c1c96a148c4d20bbf02a63e3a965a0afc04dc851c559a8bd965238cc09eda2cbceae86de5c3d1cc3e3eab11ecf13708de3fc7f910447e0e3ae41d54d905821df2e60ff6fb7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a0c5965e66b9fa4a8b42f80f6c0195194785a05e738ad15ecb6b0ac8b30fffaec27ef7a60d914b26c5cacef431fb0d63532e3382c8d415dec3f3b5eac345f7ec06a722098500f75be2f5614f170e38f55a716277e6cf75d56c3be9d69ffbe5aa31100d11d9d23d7f779f372f1818be18;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heca6e15757d21940207961f2f8b9eb7008674bef52929ef73c910d3ec3732515407ae05bbee83d12ffa6b3acc188ad9be6a90e2751275993abc2574626a434694feca01a59363726a79862dee64ab852483ae6005662052d066eacfaebb0ebb756e2bf98f8a8c8aa7e968b4c5b30eeb65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd835d238319c9733ef752a3208727c8c336140afa772ebedae5b47e2910d95410532190ffc213b55ab140e151b6c38bdd5c18f97c1f46e2abb2174e9873ef416be485ca213026723997dd976511d48d54882675399740ae98a1b27bcc6e965cad713383bce3004984f71e998ce3313050;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdff7ec0dbb3c55c653a4be4d83ce93898c3083f407f71ea10712f3dc2197e0fd811f33d571d9c72be7fda2507f8e52154fe43f0bf47a7cf4c2d6375f5e35fef8e2a97c02fce62e83cfc0c953e3923223f57cfad6982662e5cae4afe97a1ddbd1e6cf929e2625864163bb50afa4dae9638;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9a6e8666f634e75e07b096e18d60410f5af3aa50d8d15b9f958b31b5b4b5f57a57da9b007631d114cc71806df2d505deaea715b661eb19569f23eca4f401ab5c7176048417f97873850250db340e37f8df0e73ab0c13261045b641a5653181f3e72b65e77d57b177ea352b4a9f65589c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7e323b1369242dbcd31e99c0da50e2a08af029815ea851da682487a2bb794a27c01b60afa286d227e82158355eaa4f5c147a4b9b1d28018df935ebd5d291b783829519b92d56850c0191c1f418db2cb7ba8e5b60e43c21d0564265ea1305ade0db2f16d9cf771082d3152156d355304c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d66e0a5324058b8d21c5ae3c9b881e92253c11f0530adff68c3efdb4e7e5da7a4fc024bd625d1f452c34fff0a4f2237938edc50f156690fa35236c2f3e2894b1bdbf43e5d134dbe621b8065596ac6c0a4c642e8e06b272c822b627d1f01a5e80a2051c0716b60e2802e4fd2c96f90eea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35e0dea8cf73eba19713042c43df4ff9b8ac5f1ee89315e725cc1bff6bd0ca5fdbcb41206c0e531a98b449afa15e803c017d9b0ba2b442c390390b2413e1b725170f89fdde2d079f0cde9da50d8c53b699e38174fff96f75127bf3f53bf0eefea4b2411ac2bdbb2137114b91ae00c93cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69fba97c20b454b51ff0f6c4ed894d44ae77011731976e80bce037b89a4a306bafb286e6c9da7c8e3ca4f063ba36ad39fea22d107edc9ac7e3b9decbb79acad7c8371f2462cc18eb17261d789b5fd7448bc2bbe3d2d4ffcc64665650e751e577731458f98385f32fb4240fe6348a0b51d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7962ff59747d42cfd0c5e97973397ced675f782d7dddb88b469f5fd1e98377fa6e4a1394a8eee75155f2032d2306501738f1348db8e408fa27e9461e0d8d065b30a70cf36538549cbde779908fecdf6d83d2ec6cd2ec9ae532ff1a4967301332e3ccb0475a47edbc455443259130ec87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0b6a4947ea7441ab7cf078a2ed2942e25e7914ff79efe42b3ca291571d2d7c331eb3136830ac78a8e6c7200242b9ce0de7fdbf948cee4c8e989774088e513dd457ff9da389f45549e2a93348054ca16e5fbd058ed6e0f53dc93f7f502918d3f1f99d537ffdb51ddd9356ee5056e970bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87a39c76ec75d7388fa18250020d8ae472a40ea5784e58ae37e63ba8704447e89851177d1e6c519bf450c848e2f3612f271cce23765b463a31d46356935830640f5aa060b5bf8ebe8e845c6ceb07b052692235f8b89301abd55e2c20ff8cda93aa155d87ed27f9c8b5faa0269861bb50c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf25642c2fadb87f954d16d23678486a6903e6ff2b72eee4f2d7ea5ab8053367996e655f0fab3c5730e7f6c541c32193b9cb26de83bbc746e8a013d15f18a2dfb4ec8c2abe01bca346cd33c57e89478fe0048a0594c870a243e0b4e6da1c5b6dd91bee3ef47ad73ef526e6ce88e89a03f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27cb57d6d1fb2315268a0de282ab59a2b218cc1f01f78d84a1e1a92a06a0ac61dbaa322d2a5928031d0fc41c4b0c5262663b5fa8ffe88c84bdeddd87b999ccaddd7c4a256066cd01e7d218fd2195dd4dffe8b4a5f16b0886801e5964a7e3805c4e7943f464c47e32546a16ce4b91b6c4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h998c22dcc6da10b93d8f190014e37a7789b973527f17d5b780872d11e8c43f1be412804baf8dc0c801613ded1288a059b0f4a923e40ba42e4934d2af64c7c1d08ff6ddf9a1e05a5df2a5a8999cc15ece624d3f7df9f833c54dd1ba884488e7de87d173bc6c2d4eb89b78de92933ee7da9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h485deb5ae4066e4b5bf4d2324bf7f4438b347e537fdf76755b7e91d38cce84602a9189d7208a209a84da1cce40e9304f7980324d7af18bc921f7265051eb551b403d2b58a1cd9ced49b37da40c8ce8216862efeecd638eff4d05e9dd0505b8c94cd2e7d9265965d90d015143992e589af;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c836f307f24bc25142ff17d0f782fd788693202006c6dda7708ccaf6490f5fdf0983769a9905bcbad449ff7b51adac51379e543316d546d94d6b84c00a60bd0bb7027f3aec15542760fb2798db6a55b36801068995f2aff097b519c084c3cd9f90f6ad023809f7a0d9d022b8a21bdc00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6b423cfb6d18db975d7552dd979dcde8ef1200c4d7023ed5e0bf9563b9a35bb8e8102fb47f7fbb12ef37ad19c1351db9d9c2c92f235d9ef9fdb1cccb21f79c61837f7cd977e20fdf2fb145dcde761aceed56237533630400f06b202573bf43a9b93d087ba12b03d5840c244e07d61f10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c957c50b7f19588f726bfee723b73b49b390783d8f41aade9963812055bb6f7914e041e1e53d03a33a52883198c115176f57a3245ac579f7e3bb5a0fafc0f252aaf53df9c8a40a572a54b103b123e0b9d9d3b7ab8ecaa7b4ed5ed64bb701383fbb909fa7b8f86026368d2749d5682de4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37ddc4db34f6cf8c9a1108c5f2a15c5491c02bb4272256edcccf36d736e96b0bb168c8cf8315b6e9c69080b1adbe7fbf3681f3adad28d3361e52a61d1cd63dcebffc292fa6663e80cd55833255de667457b915ebf5eb27f0246e736c150050430fc9aeebd4c70fd8c4b89739ad0afe2cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e175c67520f525f179ee9508f45ec134e04996b71c1b19be750d9d7759a4faf43c3196a3589c3c50da99c6b2711dff792149b4d5ae7ba76f16e8ced1ee36af7e6b27349a96a838aff124466d02a88789ef1049a0093cedd4dcfa1178a64eee361bdea0fc33ae1a259a31c42cfe38a71a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ce06d51f25c29cb9062534c0c5390eacd0e697cb6c1a4bab55b0d484074434526f7829701c8872062af0a3e3cd8c1c0845255c1f3848769bf9b31a921090853b6d0c38936e5374a9c8e9924d91c2f1c33f99732081255d9cc339d13d7d389dc64c2f98bdb15b0f5b6caa0949a09b352b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h560926592ed504f828c5170880f2fcb84df629f5c34002cc7ad2fd015b750ecd5c1b0cabba2647a758c602d745d0556cdbacc7f0c20b5b919ec85163575e5f8da6e9c041e37f5b40520a571199454ed54c426909af563169ad595f2ea41fbcc437f32e2fb96dd6b760f08141c9f32840e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5f7f2ef1942e62ddb2ee4bdf4311e4e72755df5c036fbc68073f3b8ca4301163530f5b3ef7cca254b9b1cdf772cbe4970f7479d5d56cbd0a5c39b1150cabbc445602f32c39584fbc81f730ae785a1d0de52c7835452afe3b99d97a30a37e238bca7d072b8903a0cbbe87bd40eb284141;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d49ce5ecb1a5fe5906857a903ab0c8793693680cde592d51d94ec24a04114b02e308c8bd0475476da8d6e711d2fd124820b81ddc69c362fae87b4a30e33a2419036905400aaf736aa7a54052ec1187c56d825bef66d269d10c889d768a0b1edffb5d44500b300504f1f9c0c9a3a8761a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9de68b5aecff087b17fb5a9cf18172c2939766ae67256a5bb25d34b6a3c24caa9647615a43f348d486de152e0b21389b176852c7bd4e1b77aeb46b4e0255617b23d0a5bf1d933cb972c8c802fd7207c3509a4996a5f81c100dfb6d62cd30db242e9a21f8331a3cd2bc935295c7ad71931;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceb3f7d0d49e1b1dab3c850910ca09bcc167cd1c30a80b64d558946317590fe4c029ac2e8bf91fbb4a7d56c88c6ee240535ecc84183403c6a8f3330215a64c928c2e3a2daaae929242e9427b935ed118da64604c87a16ca6c740ebd15626577205ee3157548800370ac7af78deb8185ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38c20d28e6cedb31f94e4d89660384509cdc8d278332d409178df89e55f94784c17a32842484926ee363289e7c520550eb2cd32b903bb8ddc0c6d17b9288e98f13f45c1c02e29cb12e369df0db949cdf0c3974236b8692082329fddf273d055b3dbc3dd86c1d6d4c6aca686150251b7dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1dc78d93eef16671796a309b6e110c4ca364526c60a95056a9da7bd3bf1bec564dfde27f303de30e96d17f62f8413b690037a57ca41af5f0f43ae7fa67f057d01b7f6a473a398ad8e5fa76159495af165d5472684a5408712ab88b9383c0d31233c6ce381782dc74dd5646f135e560c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10d4a5837bb17d031e9c238cfe979adc40217979ed48c788cd76eab80c43ced727412f51a78bfc0a5387f6a7b9bd9349074242852d883dddc47bb9dde23a4b1ac2e0c3db0dc18d773a546ab59965e54a6d48e6b89c3cb663e23f600320fd931379099e81e8092c24985e315b775733337;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdba0f628de6ca749d93d4869128df21e0f51d439e1fe747b433c10f6b6cd58d722d3f24f716a53c810dc78f450cc06712001208904aa455d9722e8317c426393f02643f43d9bba94a42ef2c7d573e2c5a1d43175caf7f30f856bf4c63442d97e046c72142f63b0f7dc759537ddfc2068b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he57063104763668ddf2d378f4d5d8a24387523cdac7365b78f6ea21d39cd0142207790ce336ed061fb9384a3fee73ec3829cb255eea7b392d77643187bc6e8031e1d75295dc67ae803ed0fef2dcd1a5fde4ddf65fa11f5fec3f11b601843961cb78a9d638c0666a4996685d00858be699;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b4f93c63b8f180a3557582781edaff8411a578e6f9e3aa4c24bf0eec6c0658ed817461f507006c3abd0d3b1a78feaf4465845d01d5c32a80762b767516f00df54d667def231fec9bcad1ea24d16220c1184d9975c5f55098e61db8e0e108eb341c10b2e260317a961eef9e0263142c81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9dab4abd0cc4abd7adeb5e5baee6cc825215b0c5385cc414b3dccad31da6dc06fc0509c51159cbe96d64a8159e0235e60883f1b22b97144b433b90ef35a3fb674e88249537e75ac8177686b8fed1127310e924059209f328591beed4d9d376d15a86701adce2d2b903eec092277ebda67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha231fdf8e092f08c532db66cb61ca4e743908193bc4bb0f0677d49e3ef8f1377be8ce120aeb2ffd7a5c8fad5606275e57c2f73df01363448a80f4bebc659d31b7929f7f464b5e897b2a19bbefdd05f9550c7e9ef297249207c87310db7937345274f323dfd6727abc248ddd4ee8c3e6bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac3b464c022d6f4a4a799ad00ff25e6128052efb2d58b911ee7b3d960aff4929103442d57dfb0e7d0026562ed57695b355a548e6ba3da55075f38b506a27e4cfab9d0198817d97851c088ee8672f44284153a6869bcf592b2bf1cd6faefb14cee375497ad971c62d21e779b78646bff27;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1272b7fc95e2e5b688c197d05375bb54966bac4bc4737f134846241764e83b7fd229403d2cb938f3d5cde1d4f296f4ce82859759971e5d10320bed7d42bd1fe65432691f3fd5ee61bdde9062078588e17e661ad0d646f788db477c3f39c998b56228f5b47ab93157abffb6f2b4008eafe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h778113a73efcd4ee9bfeec382dbef00a67a345f69ed4948f3968611a054722210a60e18d6cd014b4dc788d375f892e7539348851b8e4dd98a447f17703ebef28d1ab2ba6e5f71eb61576c5f3789b4e5e77ca6a5144a7409bbdfea71fa494de909d642e75b5e9ccd4a6e3406b54ab8924f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a2204dd87f1d5ec59de9ba3b531dc4cc94387a0c9bbbf22f04384bb00ccbe792d9e6384ef44e4fd4d7ff5338d1d79056676621c7e31d31676c4134f32f588376e8e65913f8a2156f47136a3c92289f5e83e8a3e39dd7d5167d6cb43c9ba4f7d0b0f0b271b1407aab71c5fa3baa597559;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67e0c2f23b1a793ebd7d31e9ebeb938bab7a070d52e0c9af19dd5bd8bc04bdb7a746f1ea9fc8c7388edd32b49aa0b2132288f9e73b50d65f237db8da3dde52508365e05bdc1b5a7b50e80692249b7d3f5c6b97ad1e7795f4862e7c571106dac2c9296ce14a3aa687282772627a0005233;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70829a63c5ad9a69a2b930ae036e7853caccf9ac9c536c42994320b96057a81cd480defa46384300c64b95a6f47a1f003cc79c724c63dd979fb43be1780270375a9b5f1d993aec8ab28198758a90a02cfa86a565e17b9726e1b23b895889ec5512da9a14ab7f190f646ac1db21111dfdc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he44c6db3362f771be30f9d7deb1121dd2f37d4784692b24da0b8857b2a15da311ed3495dccca025207b5f8492d99abc67ebf36269f0851b894d05cb0cbdd73b97eed5beaf47c3b5bd58e3c0f81c80f8493e1b1397d41999fafad74f03bf0db686588bda248c02860c015783a98232ff66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7930b4c6e095c1928bf745f11819ded7e77a30a58be6ba97cd3103fce40ac2d07e2b7f12b7d2b582e04f45e6a5aacbcb3911af4a21113d7d7088c0a578cb54feda2287c16143878e1175570150b586ffb2aa24b821138b63924f09b571d9af1b90c0edc9b9a20eed7dc15c0360249a85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3320b82c421f978f7d46b72100c8a3bbee3b748f810e3c98a0b90e043fde0e6bdf533c1189f07cb2762e5c68bc52a87350b9ba869eb43fb54ab9cf333598476ee6fc87da8e3ce57b345ea29e371ae5468d1a3a79ee6adc2b39f2c9467c37b0db02fe0b5e45d8280ca53bc6dec0c5988;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ec2afcc18e235cc6d540cd55dce7060a514c343ffd48ebff5b3cb88bcde247be50628f7a3762dfd4ac1e3593b299b3ab6c6f5ed55ff94170f5fa50c927aed487ba276ea73319f248799a03beb93a4c53903207af5a7d128ae6b974369c9798522e2bcf7d53ae71711b2e17a102be0ed0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd57c7c7a2cb9ce8fb343510a3c2efe08fcd9670af15ff9793e86cff88ea85fd53d8ef6877cf52402fa8a2d0ebad54586cf5a566039ec0a754328e76c9de6b7e22a160e3b05095f5d021a0a084762df85b81c05262d53bd52e1e6db02d0922f66b92213ee9098bbc5da6225c91ce74da16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40d56fad43e538b235fe5c901438cf9b24bf8cc6864b0f527b26c72d898884c5eb4eccf39761ab14d38de25c00fe8f11c290c7ac64b7e054104cee874455bcdf83a2e1cb06fbae34e7dc2062f48e37ec5532230f5b0e3f612fedc775303a38bae366bac0587ef3dc8f2b123c1a4075201;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84c05ecb2e53d4a40f0fc17e71e513af40b95025fd72c318d3cca8a7d010482e8e446f8fb801698ce9173e78ce8786c0ead353b8d617f984d87ddd37ffb128aaafe38e870d4d03369d0634b367d89c7bd4c2b18ef88552d916f21da1730c649c8a0266241eb38a8a6bfcf15fcfc1aaa1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6f890a5c9d97171efc28501ecf8e334d54957727663805d4ef9b7428346e5242f86bc253f02d4db555577fd623617f10e0058721da5a07db151d1121cb5c770ffe5fb8175dd6de761147cc72cc1bc960a8132eb38fdccf1695c4d2b8b918b1be61f2e1b18f44bf69531afb48468fb10a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3458e39dc33db0248cbdc5f7e7dc4cc7d8588ec898b45a7261f14a047653d1f0043109234254b1e05befbbfc8fbfbaf1ccd570f91a246bde2fa3348365fa0559d97d8f97350c66f51dc4215ec3f4f88cb715da86df8c5fd7f77b777680a9eb640d67fffc16196fe7f12b469dcacf9faa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32d409b9e9da58c4fb8ffe9ab8cd5f51028af4c91630e3fd8fa93d2dd461ea6addb04d6804e2373fecb42f5b473480a1e8b13e101b5e53baf568b88ad516e3d51bb08b4d4b6874021a4def0f21e8e896dac13e7721daa6fd8d7d68cbf2dca9f5877529725ca0bb850e873817bb64ae400;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9598f814db8230e910456685eca4a44ed86296f29ae3b791bf3e888e54753af4a3451c05bc5055d9b9aff5e18186af0954710d726f816f5438e43057d694d26019c7bf486c82f043a5feb3fcc8d28af3447cc4031b9df03dcf685ef9921648d2701047b48850983706d0db8cd03ceee35;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf617efb2ca4da95e4641de5084a4e2cf8594b321ec39ce7f44731b7037c1b49c46bbdf89c8048805ee752052e7cba8b6357a84a3abad25a510114e3fb33e2aaa94f5e44cf34dc5d4ebf9c07f7a3bac642d0313b2a81e8892c7e1d8df98668d8f59cd1f4ef53a836246322720ccb6f5a0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4db6af45e9659ff897ec4a0695174e1be5e87127f5f9cefa421a74c54fdbf07b12f100565caf91c5a5cf6c248182dbf639f13dd3f8c2983a76f5521a033d5844f4da4f489a4a5020e99d021bb052751c887a05225eaa5299a1f0e3e0b44598aab88b419764f54c32be11e67c20bbe463;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c3504ad92d0f9c043c5e7ccd7b1d7aefb566f2dcd0d5891f311e646c3690034c01bfc3047abe21e91cb6ce02adc38bd766515e759e591bbc05d073031c46dd0182ca187a709b84babbf0864ef432d72a7b3dacd49687f582ec62c928faf0950a8493e9b69581f9b9b97115c867cc6818;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cd56aa9f526e9fe5e98d5a5ebca440918dcc129ca131fa5875f680d5cbad1afcf8309b5d62750d6ea7e64ead92d549b20c428e60381e62f667ea62f8a94530dcbb268542e47a1d8cafb00d69623f01ac5500cc3c80fd4969501633b5453276afb44413ab850f55dd2104352f6ec18286;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e7dabbab9b8d1cacab51d1176612b26753ab86d831bea7527b8767ab0ba31527b8b8ec74615d3eca4068ebf0d94f1b297e3ae80023aa26c83bc387df9a0277045acaba7507643a1f687190daab821991b80af0fb55e9cd41fab8be03f986e08a8ab48b35b6f9d1c1dffd15ccbaa663c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6fa2fc16f96709700dcafd2a1fbca8b7a851315bcd5c65bc882ebcb7e2d878e767d8c8f12f267fb9e7c364b78faa1af50e3b64e8a69911487405ed2fba9a35797d3ed04a43dd05e631bdb94fcbb8640502bd1380148b2f2e20047ddacfef8cd9c8df91b28eb7b012f28a56a2bd296a23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68f495c55800f3f0e8557fe7790facddb92d24e7862c0cab4f1c2b45d9bb726a4b2df2d2af53fe90ec3f4827531bbe731a9df3f780875abe3a326f32fd525344da29d48aeaf9d12324634bbcc0ccb01a40d9a0a481eb29f40f2f85138235336244b619217a33564598c4ab005a32b6253;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bd45573ec0ed511174790b6f8c92cbffaf0daf7874bc06d2d9c9b45a9ca3c3dde942120df2c4d4802fcfe4e775daaeeb33685f46814a060b473c1bfa6061350d7e30c30386715476f66be6c8cc2afd53cc30daae98dbbe4614ec8a2c2e159d923ac339d41ebfb63afcf68139b5ee2cf6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he72c8e048685f03010f33e4002a352df529ef568504e0f39d7c7f6bd669303c37b02b6501f48a2ec64913c8c68ff57485de686f79ed028d21fa81bacb0aa624edd8087b7befd2c523c75f9a7d778df8d7e92cd9ffdeac72beb5e85fa20709e67e3213c01a8e56d6872936b66d4931f545;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49c39c94148f54cf75828788380c589283d69cea435f21e7f8120b492e6597da4cc920f46dc231e906ba5e73ea1f96b142cb193993029caf197e4c09c50afabdade9f6358c2bafa66441f4a45e695b42c3d10d4401444a7bf67e76e845e19a57725599faf4252ee0e57c92331b6021bee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e2acc159ab705aa910985f5d75e39e17aff4b079c38b2ca310ed3602358aa290b0f807cef1b4ef562f508883ad2a050623324fda2eb2131967cbc29e64b27bed31fda2a16cc0c4e40bd24a6763b8e2345afcb2d26c0e481d0a0bafd4a7a82903889361bbbf5271719c67f43ce41be0df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a0f8285bdb37663104118e239da353de96fc77c9ed232d5a4b3cb7be86a30cc4c419fa5439e050340ac511f347393e86ea4226867def39b6eea09f615d5884a821874e033e9403d289bb4ce809189110b2bbdf1a0979ed08ca1e3ada9002d6846d0dbb652f1221c15d53ad1aa65cfb71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7b85f2fca44f5b4d4fcde470fc657deeb9b2c292945d0a57d461e78af126831aadea02f5ca230fe9e989aad861012d579c9f64bf673cfbbe8fb43e1043a4622fa2978ff9e6d5cebaf5bd06adef63d54f9589c0f6d00872d4e68bfa017591c1e7c3014cda1fe8d08d6178044a891f1175;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d9850fc30d49951bbdb7d5ab774410bfb8a38ace1ec7bac8c7fa8ec48f3cdadf1cc51b813ce199355abc674f3a3e77f278fd5468125390fd0c6a44b8b104f368fb1e70183ac0b858d881304e77c04791760e2d17718459646a685853c090cbb2987d08213c87670688ed29e88976ac33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74234a61d21b2ec5c05ac2cf401ceac97070a10610d8cfcd9f03ba8016bee846e793f0e85ece9648ab4ce8ad313500cf481fa3d55616edb3693e90d577afd2d111d2d480cca3422791a76eb20e4992933ce03f9ce39f6b099c6537e88e7ec61f09744c39567d549a2811a6759ce6f5bfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a9935c345e8f85af61cac045486425f64f9b1e55500f9434e69c18eb144235051b2098cea29ab1deb728720b22c22fab7cbd9685fad97d500fed0ed6437c6c1922e7133b0dc4e5cc06c403f3b1e04baa863a939266c07ae8cff6f0041fc7f26e528b8fe29513a46d3d3faf114b8ebef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1a1f9048d3622206b9028adb5ed6b40df3fe9251b32926dd90d9876103eebb728332438f21be3b98efb6c35f766426bc13741d8405ce127e1b260b3657b86ee7bbeb3c9a3b077468da11846fd656af37e2a875a0f80578a78264048e4bb1d6a797160ab6ad5bfcd34fd8a96b317757da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3761ca7d0b83c450e6586d81493a394757976b1053bf3a63c354e094df767ac716e888d8cde5ccd1cea1dd013e4bdff23aa9a064ce1a747c3417ec56b0a115b67b2c4ca57a7a393d25880f8fff4bcc5adb73ba32bcde8c42271e869a31d2bfa303d39107225e1ba7211c43afa2665adc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb418c11d06acadc3dbfba0dd3a8655e45348e641d625096ed6728aceb5c20a6711981ab55d303989da799b0fde5cb5d478ba917cac8a2d9e1fb98c0f74f4cfa2b7350f7989b09ad188024736a10db72c2e037e2ffc92c5a54770262eb46fd87a43f50f3e8f9b44b27a524efd94d37dfe4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe3ffa29e5e029ddb48b6dbe0a24fb2357ce2abdf89debb942099d2c635f23be42952c89e0354da3065fa0944bc3383c2b372ce92bd9412efa9e74e2beea3aaca5d5aeffc60c66613d9b60f1f063dc8d408794e4e2651b59f71a6d26b4f0a5482e59c5535ed8c706a4b89eae97e4451bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe60e71094b5546bf0212f1b2bcc72c3b0932f5de8186d3db417b10292154a52f0dd6e58ab38a9b8e1c4f4bdc7f543dd9dcf526474c8ce8e8ea8b8c2eb66a01e9a13aa4eef62bf32d20641236e08f7068a630192ed59778272c4ccaf9c19c0d406013104a9829d68d4ed3c8904e207202;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae3f6d25871a08acb3c6771bca747fdb8e1141229bf3133d5029a3ce33b9e79bcf34d59d55054fd8583632715ab23c9c2446c5baa39537b316ff5f60a4e12d10ee31a376f30eff36badd0e0c97d5ede08d943e081f5a3d07ec2e515f958ce4daa2ab28d975bb15071b969685ee4e22822;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he29748cf2a79082c792524ae148e36e031abb5554ab8a70ba002f6253fbea61bcb2dc527cf1ed90d79ea724d520114f3719e2e1c9f20aa0ffa7222ce4c317f3b1525ec1bf175389d2a0447c6975f932d35687436323263daa78ab4b61a1a0441d86b60e06d77e481b8413b70d61dac6f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50de2e1f752ec64275fa1a5d8f292cc31f3b3750011777c91ececcf72bf257c9312f7d71f7f791d245e4c868cf4784d99fe725f7799b5e8f99bd48c86837ecbd021b5fdcd92b8a5e18dd2dcfba35f236da55815d53245a5fe3382c570a687fa6e3fb320aee61a1c0b50a858c6c31089f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc66fd22127867ea9f7ad9df7be3a5138062ae82541b48f14f61bb41a80553f78e66d649de1f09bb2587662b990d7f5a04046cb3b2e05f6f2c346b2d7c5978088275aeeb33d5643af759099f024a9a8b2dd38b48b977f7d15dfc833bdc2e20ba955164498148b9e78cf5515c49fcec0c3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcecf06fbf2d659d9af1c9c2a98ce8b3cf092f3539f0c5f4dab861467314989df6d9998c1c5ac5fc1a2661a946e659f1cab251ab35934f08d4c7c9cf662618a1bb309a12ba16bb1cd5981aabf2d8b9400f45806bd27aacab48a404552f7107709ea3d6edb54b81d4f5c297469fa86d353c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c0515a96ab83aa4e45d4050623d25ad26fbd986a34a0789f0f4fe17a94421ec6e131e2da13f4b0a16078074e60e2b90442c46d2975afa169dfcedb760e19e34ec7feb687909dcec51d8159f68c9772a3c4d5db8c8c0110083fe31d791f63d68fc2dadb58229ce0a7faf971509d41a762;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95b6b7144c97e96f13c6782c2379ca3aecbf12ebeb81a18315e090fed17a63406d28c7f539894727304df30165c8c0ab0960922ca9894b4ed7351b14d3321bac3888e3fe66e94c06a6553178412d8959f3518d05cdee049a5b43caed03d0d26032102859dab07ccff013eb60f9e8291ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66af9b5b51e54d34f3b7a25305b4c2106bc58f6a83bfeb0b1ae6d507c64fe51eac7cd7a8373472249d1735b477feba7ff78a552f613b931a11770ed31eeb02b213141b434ca4402ba1f4d73c6cafbba125f29a36f3f7d0f13faf82ab57502bbaa8ff31fef92b716799b68ee2fa17c8f88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h660d91f0f58aff1eee9bb29481de5cf00a5cc75f0ba3d9358c2b215d38700f1c260e6640513a471db8adfa634ab31192f2a526e4fb94845649864c0fabe174d2e6f631743b59d577d700396357b7e3d15bb8c0116055325ca8a478debe92cf19cfceedb35ae8a87b317982b40393c2446;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3411041bbf03443017b17145264591e07a8ff8eea32c10ebba9fadb5df649815f8bd8a11b9b4dda6e3b7eb8ebd91b91d77fd42378e4e538b36176187ff772aadd132a25c88baa2f7d9064c32daa84044d84c5c1f9c52be652e3c5c9393be0f597a4b9fbab1d2a8e889c123fb010cfbf9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d4e762d8e1416a1760fe50c8e02a9f15567b0cf75688d14ca04f0cf8060cd4d41a5e24aa903260dee8ca0539b9ad03c4e9367e5861e88c9744a32c0c6997bc3ba1cb3b84fb7a2a0a3adbb433b9c2f881de878bd8bcfce2128b3f02e0353bcd84691604c18baa0ced471266682319e9e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc86958d23388a47a5b7a1420c429f12c2e57bc2677131ae365e23c88ff98eb137ff87f4e64b771c480316cd3e2baf176805583650e5f786178ec7d25e746abd9c4815ac855c4c582b34a29b3fc70bac606c9f765f8c569166f05b476f8ee9e071d441857eeeba1db41b44f659902748aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b9258c158d6dd46aa4d346098bedf9fb6ba21ebe0dc2d5a3d26171d2bc7a7f876c77d0791bedb506521d6a6c955959cfc47ea085a3c9614456ce9cf28ec9460e18a09e443c1e48dc3216ec1b4c60e1257e81499cee4cbedaaf097d5f7204a53a32451b85a1108ca1b4e4476fe14fe544;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6aadd1aa98fe759e52975453bd653e8a0ce794efc17c0bb16bab2ba897f42d7b352222e8f2cd925efda3c1c86e2899eea624c5cef32af2b646086af0727348609ae4308193316189f216c9dcb9d220baa6019570862fa8608fb4eaad2dcb9b19f76cb93462e79a851d8d41c8d29b229d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfd5a0b713e1bf1ba5f1631df67f9227342411f67c638b8f9fb7d22302a22f5471f20affb13a416fa10a64a9b45ccaf33b922c512bb606266820ff7a943a253f1153d6b712bbef8e8beeb692349bdf63432110096e51505d1aee6a54916b399635571062c0c08b8949095580dbb3727fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha98b62140a03259946963d8ab602ea172c0cbf677c52b6979e79b7235ae7a5df7c2d3c36f11ee11c9fac3f27c0fe6c3968474e72aacf65691db8d02ee3bca413560a28aced26ecbe08e950935b4eca377a73a77a5afa25aedfdc07626ed86946a28ae8cd4836681b6d136365980a2a8ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc22e7b65390c45819887235b1219628f9c746dd369856fab8789e288a0475cec1bf46eaf65c10ace5e322a536ea883b5282b5090bce19dffdb0d1b7aa6a1419d58f416f0a4a4cb371423c7685db53b7495e5ddd0fa43ca74ff828df50819154077c33daf75c45d46d0846a9862059e04;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f001bb36f199425974dad2c622c7963df8fc5fe070e153028760b6546fef8a2c1aa1fc884523f0a96a16a38f60bdff22f1dbf28e54f3e6f55185761d7733be6394b8c8c0094dd86d0cf8d5782d8771e738728e3b0956e46baff619a4b3c9c9d6af56481bd2378f2165ef1d40c350278;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36a6057f115b54c5c5d0f8cc89b7f908f40978eeea8331ecd0fec37fd0d8e051464b9bb669a96506062076c0095c99df6ad0111a5b907dd1b2fdcd237ddba1c195def2a7a33c936af37ff35c8c0c479bf8ba3043b2cfd4109f13ec3b799b3312d0a77dce0eccae6055c978f4f91508969;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d5587bcbb80e5c9e0af0af9fc516e20f8f937f137e086047c1163c73ab79a0546c76b8dcb350dab4fcada8e09beaea5a1f3a1e6c253deedbf1a2fc0f5d73e9cc7459d52b74a76932dc75a32dfd4689c93bf70d22b54284110d89355f2e0186173f7d3f59a066498d03224dac378fc5b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9acdeeeae6a21c5f033051dc450fce5516570a1f8eb5788f7945795030292eda2041074599d3cb13e46d011b9d6e7234c9154950c39d44a0fe18195882f88b2b860cfdc509e85d6fe28f6f430e8a5c0e8a257d7d094d6397ae05b94ccd73ea30ad2dfe5bc73e7aedb67593ee8909a784d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a5351699548317c9267b118ba7abf3fafae9e1e62391d49cf625d08c954ed93caf76d4009c62304c0342ad21fc4faf3105eff4d1aabc7f01be4df361527cf667f2ea63053290c746b3fb147cf158c9a1d16feb65bf7a1a259f7eb4267b228043c22b182c434f53f21e5f3bceed2e0a4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83ffaf9924f997a35077b0f643d36dd15293bf88304e5affe15a3ae21d945e4a69e08703bc9825c5ee55b836950a53978c3309d2e76b7cd7140a74082b8b09e833a5b21caa9781f2c18cb58e850c8da5939108fd3e31822ab40d7d32d6f779f5857a80d935f4843fdf867ce2371d5cfc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h497fcad932923c258b80da5f248dde44c2fa2e0a506e7847e9dc9016486dcabe764c636e687e4ff64fa6d59aea430a59432efcfef0b4cb960689d6096a4e87ffe582213f368c118acc531653ac4fb3fcfd2f9da536cdb15e59eec3495e9d66c8137943a7cdde6c6bb028cbc6f491d8690;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55934f5d7c3e07682accd4318afd45dd4ce7dac2b83f6e0f4a815fc3a3cb50052c7948e408eaaa60f55a7999622c5338ab8905c798df8f8c86dfadb0feac60ef459ee3f45a5c9e6d2634683414b179773d3449ba100120f3565e305c26e1101c3799db110403f607fae7e2145e523e33b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf24355784c27827299135cc9305c11f127a3052ea76fff9bb6d4e1a0f0ec7ab5b892aff8464c7931a169c05515933201ae13aabfc9f56458a7fa90d93d810fb17df871df15a5bbe8d9fa6f185651c745cfa52f322f1b3678a3a133d435ab22115ae15cf1ea66c8593a320608f32d95dae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ed3aec70a80fae9f13857d763829a2b367894c80a2b06c1c01ca24516a3f32d0f4b594d716b92328d118c5e6d7c4153a2dbfc15cfffe2702c2e27f2ba0f01048dcc872174dc02222f094fb4d1f6e15deee2845c390f5c860e01a4f697257f0c1d045e4d0e48a38d27c50efa24ad66a53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32e142cf64d10c93f0493f91225014cc99a452bfc0d12749139c1251c1ea5d5de59174e280d3561ca036b17172bf0b73117791e8da4139e5ba80efcf28b11c46fdd75426b8bfff927560241b575983dbb0c45578b3d42e2202ead8edb90d8936e20263ffdff3d20c140ef0fefcc683c82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc81138620d4ccdc2b62de6fa0822d218d9f43ee22c0368442109d287a4eea9da167f50a7630c0c6d054d0a8ef53e49d72852ca05275356eb9076d45358fb6d26b8ea3e6eb616033cf4227032ad38b29be7a41e3440c5ee59d4e91aa313857163e24cd189b74065c59ca596ea24d850955;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1024352fab34b57292cab7c7bce3d47a46962f1fd654eec21f8c701d1f9a8aec39d0678a7d0f6de7e6759a92ab6bfa958ea8181573351dcb5f6443ae832929427cca3db7fc661878ada2fcb88f311f215667d4dd7f109d1cc8afc9080205211ed9f4515b8464eb0bdcba79d5a28bc7705;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ae4f1292191321d1f258803e6856b855729bc3032b70aa9271ebc081555031c72cb76697591a0f1239937c736ff7dfd6b27a6900d20ca395d94cccfcd2f916f859d5239adca25e124033cd104c711e1d1611fd1289d36f413fbdc77501a0815ba317e5a0c29779bb97b76eb0cd9ba33f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc115401ec18be5f17918ee509e342eebbdbf104902d39a991e881cefd0ad71da360444855a445518af8508e6a4b6ec81a18626890370d74bdac34bc7cb9dfcd31e9624676a5db637bf4ffc2dd7454066b027bdb348da7808c2e1c671b8289899fb3fa4b6a962c2bf5d80280deffdccf87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7315df20ab63f5afaec1d0f5a79046cfe0440e5c2c6a476993f320cf9c7a4e0e56130b709fb5f451c52b3572b68d7e804330925617eb558c0330b71294aa67bd3a0259cc6d7c99844057a30c3c08a96b12a72b038a319446b01813bf2a981d497e76274605ece8fa79e8b6145893846e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bf37c2a814b66a15ef763810a2fd2a59c3fd6e0c11bf960bbda19793e195dae5b9959a3fe8850be9d014e7dedac33e83dba446604c5f3dc398295d70e6cea5c3552c605e72a35fb7c4979c1b6d10c759c9a85ee1bd5d94abfc7a0f7427769ccc7b6a1425f6fed3254422d4735391c0ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23c6ccb57ac3b44843e4e99bc3f2a95a7a21855e30879d7d0ee588bf1e5f6f23c7bd7ba35b9aa14caeb28b17400df47f8ae57997527b457a36286ef8eeaeed598b0dbdac7c0ded00d29622bbea01b4fcdb054453cce7e854dcea0a0d28edd65ac8f757b9b7191022c0f279bfbca7edc4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59fc98d9877efa2f629800db549fe5504d4b361fd6fc46f1018f27442978a25c94144122bc8e5c0a0656e6e17d3df3415cff4c3255058ca80755697f77016b568dd365c484d3446edc4494a3ee448fe57bfc761fe67143ac8e01a070e275612e688a90f5aca558289f449446779b6b7aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he74e25ae314e7ca0d33697135e4eb087647f9d565d2ec42e6add9aa78d0fda45b255d9eef6cbb53a77651d07c609aa8bc31c88194c2565b64b2e08bae36c76915e2e605eaa47027018a7071648d2db017a0ff72ecfb4fee227bcb7c1faaafe0092f91382f1d654e44731945d2aeb035b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a29465ba0cd7ac7b9df17039db2ae8c0fa80fb57d6ad8bf5b5bf495d5fd9ea01f5bad097da4bf71452c86b075fd303ab45a83e8f92a85193f509d856953d0b0aea87787aaa661ca9b2103e2a2ec96a6a25b9078649651e6bd7f538c2bc116aac4d72851e26bc0196a881750496c8214d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2644987409b76635f3af3091d9dc89bc18522f05fc8a87dabd86c617838df468506fafdb958906b5df649b3b830a0733655d70db47eebddea391e7a60c10471f972b4bf06607b1f959404dca28b54c0f489e9a71d58ff4928a62aca1182c15ec0dcb18ca27d2f1bf0b84bbfe9150377bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h654f2db4b3ad20fcde896f8e1d664394c6fb38b36dac9fafc0b575f029e9a6131421e266904977ca17fa9ad31f0465b61e92043ed9aaf05ca79499ebce1973671956acf7eb80c2d8402bd74b58aba0c6eecebb0322178caaa86272ee0057307124057ebc24a424ea456132b5535e29d17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85376a25adcd84b20b56f1306a269d156f0da95cea7406d3fd74cbe18cbe645c49bea13e6f8c8aceed36c23c451619bd33573fc5864b45ae01550414d191ea37bd04058e08fd867178caac8e90fb81ea486080c931434758f76ce4e02329d14d122e38f51b988c613b7c856b8698b9e05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34407e7c9cc28d984895b50569261493396dd0d60ccfa6bad1e3c1ef839f8356373d193a83c9076b47e1099cb4a207a5a9b77af0a00984f1d6342df2fe74684af9087144f95568bc636071214bdaee8f9286b1dd99467ed724028f32eab444db119b5491171e95858ebac1de33c2fc186;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16f4cd4cabc857e700a5785103d13d0ec77494b328f215d5e0a9874238600685641ba0ea960b324cbbd8d0ecf99b47619af8506f8e654fd49b9bbb83489a392e6752bc3b4fa09f4c8a2a58fca4a1e6e8b42585f80b7979983de0b3d0b6c067468f467b24228b65c49f0f96c3655086fee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf01bfc8c4e458d8561040f1664bc6ec8c0cc8933e01708fa4754ddec1c27ec73ed25ff875efd6f503981ed00fd1e9350b2755f20bdbaab4970e4392a5b721a2dcab3fe09c186f7a023a1d106bb1e8427236767888c723af968971a0a3208c8c869d05ffb5e1f0e6c9a28ad484d3d6afc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda0369b901649bfdb58c4e7f85d888203053d517a725d99ae2ee3e90de9b88d1d8106f968cdbc8d7d2d93df951771de8f7bf0935fc62118ea5453d8ea9eb78a5120437cd323a40b6b2c581ce8e925fc4ef7d15c7894f97689e9ef107a531e463fc2e7f35c614b7359deb72001d8563024;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc791ad7274b8023810176b3ae99ae63f32824b91f73fa0913459f727429b017855e5d6f01d5ff9a65c51bd4765261478282120e49fcfe27402c8c2e2922f79edbf32673032dde8b379ab2b192c2caafc60ad95ed0f456d9347444643faf998ae99bc7d060b9d04256ab4970d272dc64b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fbf8a16d7d11fd24bfdc274fd058aaf5eb379bd122b825fe5ae01d7a3df7cd555c11eff16b6f36f9f3ca2a9fd1ef6c09d1132295aa58893921ae952b0ffa79e12fc75c1919ba2373794fae307c564d85e2084d01810d5706c6dfd0e5f6f73a55662071fcddcbc13bbf4a55011ad4c91f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haadfc912829cabc9ad2e99792b94965790861e88488d3d10dcc034d08268f0224f4bfbcc10a099ccd6fd79a37dc1e94259bc9ddfd200c66446dff9f7b21535c1ebaa8a361515de4c8c1a551976be6e7902fa5a3b9570a069d72ecbd5aa21f5826fd4f5b79b68f8b9f0e6d77f5e1971eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71ff9a91063f2772078587dd0f79ee4012603ca0df71e445878d53307e7febd421ec22a35e5be33ef3f080c8050758df7eb528d62149c94da368584c94cddc0b193e1c9905a79b5798162ccc7ffa60087f16052f8b17c08d3641206dc0734beaa6986c9a081dae9f56e23c803d566cdce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h397b64e6ae408fa724b0f6ec55b23703f915b4ca753d0071b1ec6f23057e69c42f3a837988a2a9e5cba2532706d611e59a3846372fdd34f4ce34f3d665e80da642db4115ed0553c1d29f2fb4aed4d7e11760bd554acb12fb52da473e48d4e19baa21838ea894698471b9ddee4669664d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41da97a62a3afcb729e5f1b0b28e81d99d9e4e76d91b4cabedfb2a7886b47d372ad4853f84a1b0b836fee52eea318df1bb447ec2b8b8e98ae85b3e7da00797a0583704f0de3cf7505609e471930a6955d4cc3e3743c23d48761b117a6f783aa6a7e05b0ce286b5460449ad740a8d4cb1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39d3722799f24fa95bc6c45ea5e7c227b47d9c34f018da91ef8b176b9b7e967287956b76f3aad4d3592e8d10446dcdca1ae9228d9cec5744e8f30f7d984503ed793eed4a5d075a828bf706bfb43035afe88934a9f3558feffe808ec3712b0b0708b55ee2ebe87e5dfb94aa21e8592c870;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62b018fdcf979d81baa01b90bb157536c2845231cbe9c8d3d6f453d3ca776be8dc6a9c6234e05222f24419cdc7e2f1d97d52710f927b6539ca92e369408e15009919e86926f16fc3ce14234a109d66b9e4396212888e3e39f496964d44fd5f74441d83b684a14efae7706981d70527321;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7e131785234f5bcbc95e4ba83fc573cf5b54711441a4dc31169d99744e5d89c2bab0a6edcb7d97b77d0f184e95835f52b86d91891c7a033a135a4bf1adb0a24d813a727da218deea98df1bb0353d638be02e26d1f633479ac1d94d08deada7193933bd17712c891cc4e4e3c864368b87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aa8b3d848aa8d6e422c0e179b7a1ad3d69dabaa3bbef7eebc835b7b3a6cea77e49714c16be3dd534078f2ad458f3443c3c54b1c97b2654268cb8f81ad71fe000c9a4a222716ffc262a9f1c8e13011ed8862a68c71e94d0cf721eee0b82c307c5e08b55b6a900687f62b3091a1cc6ea25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95e522e80acaeb463b29265c7438e0e0b07cd24204920958c15c20f336349dbf9e6f385de83856a789a7e6f47f6bd2c988b745729b45ba2e99209b430144bbc366a0261ad6ac0a0b54ca7639483fe96689d6fb0763f1a0b8132f1a17f62089cb9338cf26a8d87d24cd84fb4800713459d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h880f578b7dc2f4e29e48399587c2bc01a871e71fe088a55bdc5c946935b2974a1ea35038968ca7f2b549dc1c1846c71e1ba17c9a930a8e5b8adba01ee93b4ed96d3ef47fd08e373c748ffcded37be9dd4e0ce6810914a1419e74521d4c55f64f33bcf477e61ffe02c8d2406c1d1b84643;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he63bc933435bb2de757f742d0f40e756d82e603d22668f8cab3f57834cd1284af3a2ad9636daba848e771e42eaf4ab2082f6600b253734957882afb78cc1f1704200fd04a5407356cf7c7d0d7fd7f6fb0de5375e92e5a094bfaf8c0e7e7f5b8cff6bdbcca370639e235192bd16c319f17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dd1bfa91fb52d7171d37e60e0a82407d7c2dd7be8a75aabf2f4172ded52768705ac980cb011a3b7df829a088931865d38c25c19a0df13576657e6d06048112e4ed2a032261b06196966d1603a7393b7e07d9478e95ae59b0b881e1aef1f0db2c1f6590c440ecbed7d0d4bcb472e13555;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13128d140b6988a3346a1d0ed8385f9bffd4dce88e484ffbd00a354fd491b52ce23aea1cdbfa501b13a2fb9d35986233522d54cc449bb80fa842c47601e6fec560b8ca0cb070a7c4f5947d7dbdc419e72c0acd5f52e78b1401e03b6afd250808dafef5aaa5a338206d663339adc2547ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe15befa22bf7fc7fda7ed44bc6ef4cc79cd0836ccb341791ee072f777ba85a4fe29d74a4a1ccc26d1076a93ffde2656fdd2f020669dcc7b068948b772f8745449350d2218e08d3bae6d108004aa0517f8d6da831d31f7f7117a87d06ee55a918ccf68b6316f0efca8017f1ce54e80382;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeffc6734926bae5084769833cfffd9575938a34328d4d668050d969c34ae6974da6f9b4d555422a65e4a5f49c0e4a98d4801797d769950f12b01327486b21b6e1ebc7e7fd97db5f3d944b3c4c373f26c01f2b4dd02b53725a23e7c564207577948385f43655868a1fe262782b4768c93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b2299ab3bc15ae33d27f7dc3983718a4358eb44c192a6a7c7aeddaf9cc6ea312a11698053fd6f5ed11ecad4d30b34d5908a3acdb60ea216a41382c08b45fcf0c4c0deecb7b5645ea872719c1b0359f2f89bde723f10dfcb63bd9328b5afed5bca72bc9992484ddbca1ac1db8e7e9b06c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ab39a300237e773b0d958678c02c8fb899651928e692a9a912e19e85f8d42e9d9d17a07036280c8391e612803e9998d028df42317771097b8167f750580fc50c0a7891adf9af323ee1ab8530e11366af56d9a415e0fe4a0fdc887401d0746c8ac09c2103d0bc5d3c4393645b7cf86141;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h716fdedf5cdf8651eec953f71b0b323cd439ae12ac4bf713fc5c6b3e10691d8e76191e3bd3970b7bc7edf8dc231a6f81a1f3a5fc7e365406741c1164ac2d8c41e38889ed8bfac46d7d3a1de5bb081ae128d918a6abef439e01acc7fde044af61776c32a22036b0e1533837744e53f0659;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbc3b2dcf476d9eb0f12ff0693132f3443a9ffb9cc2c414260b27c3c4248bc9f3bc8234d0410162f5b65cfc30f7e077ce3c5dcc6404544253c4e95f012b096343dd5870637fc1565ab6c7daedc4c79037aabb23fca53148395fa39d7ed8d7726555bc5d05651870e37b87163310a6a6ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd88762e56225b877fb6e366c254408c7861579f847835cf65b2bae46a1068347fa09b48ab748dc1582c85ae21bbeb2469eeb9052119ddc4089a2616a12ba321d39750d3f0428c442f1118d2b3a3011c84513e8e12649eff14e7b00b42177534c1dc588a2965020160310449849d9f8818;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2a4cdf809038e8eedb1d2e5e2af2b35c152c56cd5c9d97959d8f1e552bf10d20db1e97556b310fb4ba52af5b26d1c63aed4b81ceb289b4bc180b33d207f87ba0042e7b2d431384c1c40426619a475a957a11446b972bfcf454d06c718e0baaa90ad0b46c3ab8a8898d53cd72c6758668;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31fc9427fbcd2855a9d0d8c3ff4547938bb5ab325f6a13dcf189d68b613eeec200e2fc3fd4a3f1d264c3af9223a5e190d954d86e979b6fc465d2e2a0fdbb637a9fa6c18300d8ee1dd2527b1c4c2462fcd07aa14d159a7741c5181a1cf48f9a0b547db1325d58ef25c46eaa6c796c395b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8402eb72e515fdbba28b48706a5cd6bf1b42e218d3b6dd2a26ccbfe78b1e738031688076365e7fddd0352fe32ae8c856d7ef453dcd3a57788e84029ea3c5dcf61f3fe84aed4baeae0196d909a92695fc1b381b8507297e6de46de6a2a6868632d2d926eced5040b19d4f1be2a4eecbde;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha572d3f7ecafb84ccbbf92f3ef16b0f200a0c25247b1c823f86594518f4ba2b7c3b9c331bbeddbc65992b520aafb0e9c560869b672984f02ae4754d263af450f11ca21b314b5f68f3dbf798e4684b535ea57391601fb44ee31b36074c56bb0b0145427371ee852e50a9d083edfbde9221;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf0f2c5fbfdc287dd8a7545e6865bd36132b92a3e2569a862ebec6b2e1475d5df270db555da98786f6f01d2ddd780646d812a9fb370569adb3f07e64ef231b42d724457aa1d3c465227125450ace3c6e6c835ab095b9f883cb721242ef819e2276119c169ccea939bd739eff85f076911;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7694f2c20a6989b48b9a7e7a32811c4f2ab046a66b33e90811f8012c583235e965f4536b770d07f5f94b6da1713cfaee382304ddc95dd82c51c922379a8412be7f3556a0e40ff65c5711846863e4424a07bf4a9e9c88830bd06ab4877f0d2fd643535909161368a48a3ef3e48098c3b4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47e06d8895b5ad6871860b11fd3daa10d340d2e33a8de1e69a9fed29c4d1a4a5312a166e0d8350a5fb6f473cce0baff5ce4173d1501cab3a68135c65d00ce7c494a0bd0b41f4acaac129944387f34c0f3fc5e0bb993945ac9216e691232bb2aa9ea7062cf7cf5544ce8b632cda19d8402;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab5ebbe95fd2c61d6941d9b67a3af4e1d6bc70ed0ef7d80a2e61c77dfbd2088fd7d69c723f1fbf2b6c6ccd03936d49cafd901527820ee3b3c87e6302c1cb21cb305b44d04fb77c4a748b9bf652241f0625f82b21f162a3619f8d5d7ae9f5901f3fd79e5d6992e652539209f6719b443f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29285458e0e93e3d748e1b189797582054a4229cb7b51dfac1e01dce022c4ffee3e4666bc0b5a90b868eed5d27d0f9d5cee7fa2ad0d60c4b43ee3bab6ebe1d97f542397dddc494445181d0fa8e17b61aff90a40c1e4c67f0ac5b2489b2ce8e9271427c458f21ebe7ec93049ac0d650af0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he060215e19cf8e8aa2685046868cc060a211bb9f6c87990326d3e93af353ba61ca524cd74ccfddf33e231de1f4ef41a27dc92de2ed3bf044bf73e313ff16862c7e38adeb9b110c0e966ee4b97745d74224f3518126db73a539aa7478a9a2d103157ed17406f09a65c1ad21eea6ba9ccb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49651c50f833ba977f0ab0046b26c27b7ac44d3329f26f6cf3bea3270b84aa8dd19b1a494b33c9566485986707f73273359440d80ac20aad4a71f2dd867ecd567831f99d35d62b202a73b0a59457e1e6194541fde869e54abe40b6388ba7468f6fba6527f6658005a48e29ae449d6184b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4929dfb7e174e3a57769b03ab21eb406061991c0db1da989541267c58543cc11f88acf11d5f119a77987c98685afa71b067d65b37462310cf75e9e60bea937ca3fe2067ba31aee259fa1ae3691608ee6e8dd34c377cb76b5aeda7651c381f4a879b8898e4edb5e728c0467d94026229b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eed0f98b213597ee38ae00983ffca60d38cd0251836bcaf211a0b70e7cac21e32cbf673c81cfbf4a748d037598d507122f9d618a0345576260d431637b9f3768a666abf92776720776bd640f4699e6de533e031ea532fc5312cac7edb970aa8e19008a3540896fc982d247516d3b7c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h660a443937644ceca06f9b482fbf8bec1e47c37c5ad4fe212e1b2d5e553d4f3a6f22ec96af86426f43eebf427c4a9a464afe0aab3acb10a17f738eb0fff3fc8fed3197ff643ddae1e160cecd2a4d245b9cd36857652e0e39b9b684d78f9b6be7500b8100a8251c784b8cc9dfe284888a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h482658a34f18a5a3fc1414bc5f0995d809445512c860e877f2f5595c31e91874ffe5500515d58ea4d73e695659d9298b660cd7d74c73fe599d5dd851d6ea4e28f3185c2c9fd49fb977543d1eace889495647f96226ec4ff25806833e080ffd42b8f5160f83933d9905b1d3fb1e540fdfa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h767fe31243fd4ed968e814469a956b7696dfe058488e73704cb256a6e30b5800f8e5768396b65b1243707c597738cf6d186acb7e8da1622df7832866a3e616affeb7f7df32a9b0b5f6710238901d76effb655b8b8a48dadd203b84cd59c248bce819aca4fbe96f011d425a9b0d6829869;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde95f6ade008d9a84fed6a1df12d7264715b8a73fccbcbad02be86db57e050f684508a42bcebff194733d2d7b5144f519d048d5d0678141beb7f164e01352f7f011f47183d01a862471c50d42898e83018a0b16f96665d26c053ff0d416e3bba9e63a6f0b95d6e01642d8f8dcf00d7255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h335ab0a1352fe069522275b91b85906c370e1e65e9346a46388539c2d16abd9ce9282ead8fbce3bd47fb31ea0a8af9416c9469b6d239972f88120964ba8e2fefe2fef18ff038f11388d5b6fdf99fa0eeae0be8f623a32ee49830dbb9fbaba1eff69885b78e0946096e6aa457dbfa8592a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61a8c29c68ff9c490d029e55807d1ee7f14aa9300ab37e9b41bed06646974b1082eee6d81a08eefea620fcbdbba87d26cdf9437272573806680e1366f14d2a97a53c6ceb14e0a7f77d96c54813e65534c230f4712bccb3a9b537455c708312c856343655adf9e3bd6fc1a69c1810fb694;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c0da9029a1f765ee4aeb9e3864bbafad4b5580b7e4d86c6fc65ee1e8ce5caf04ebd8522080a9531eeaa5309badf96153da3c163fe564d185629bd3b8fdb5c7aa4b5ab676b63aae6f7821306dacbe9a7269f646632ca68993f36ba5af9636616fe724fc43219c1f445c61993dcb9f5e4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f10974152b50bc565e17e37d7695da88cab40e2d0a314054dde6f92adc3f50bce292f853d79c3ecc4ff081c5c92e69506de0e7b73b032a6158156a246756d45ed5d4490e3cdaef646d8f9ef2b57e407640a2834fbb98b9c964d0cbf645d41ed60c61a5a3f4dadc9d41c33a428f0b7c4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf65fd0a08b8e2ca34e6510ead825ac626f929e4338d40a119582ef85c9ad415317295c8fa5b868c9f66420841e2d667fda68826f9cd61f614380b1ded65b642cb7897f8743d3e84967bee15537f4e1b2c250883aafdda34b06e87d3f3cd39833715f3de1faa792e5e3eb77e99c358d03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4738ae98b5fb7869a21c240c3bb4a59b8999be85a4d52019d4cfa0e2b13de0ae6bb65b601a75c69e347678966bc1de90915d52d0f7c6cb7ef2b48e9dff0001ec88da6c93cbb07bdbe5d2fae21b022479390d72a15edca4cc7128d5cb25513f8e98b3955ba4f5d62ab749bc2daf68a20f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb325e7ecc003d136a6c2c651879373361300260b2d787ea3c00190da0e286e62efc6064e18bf3e098e01fbadf7c6642ba6ccef5960b76a873314d98d9e9acac4d3db90ce4e92f28f0c9d6e0fd2092bc23acccf2ca87491df76c97694a116163b7e28d665bbe29701ead5ae7bbe2e8c7bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ed2cc9412fc5bdd05712ca2637b5fcb4cd52dc7dabdd861e784341ab59e2c8488cef07c2ea6dfff09ee0f92beeaf34b65ac4eda0542220c90740531bc4461ae724751ee59e7d55508951861e824c6a1541d7c1b120c2471c9b4122dfdb7a208ef4bd4dafed2c61afd7f432f0f7effd26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e33b7c99ba4fab8248111a02f5946f26494f4c5ed51c8a8615f7474f2b964ef8d52bf23ae72d17ec264ef7d14e091502483ad5818351f38cb47d0bf217d773705e5f65571fe012f100fec8e413903370469a35cdc5c92f0c782a37086f410e4a833b21f1a6efb4a7124f2ba67e40708f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c443106908d14e6ccf33c978c519d90e7ae1b0ae1737e91f1e5eb321efbe69972a9e3b3065dc08f1e79de58fa2ed55d519e39dbf44025df744f6068484a8aede33da89cfb88c75c29a570146a0a22742942bb404a5976938c5589490e44784dabcef9317fc07905a03e90e6eb74bf330;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3bd0fe8e14559482784d26c1d90e2a22b437a52ead7fdedfd2e1164ac4942dfb3bc7bbe2f4dc9dcb54031844be7c9d386d1608fb99bc6efbf62377f9c95d36358dc172b1cdc7766d5d7f9b9439cacd6e7b79f53b44e74496cb3cf6f0002f58ea79442f5b51d8caa49d4e9b6d7ca5739d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92cc0d8c7bdf3ee7279346953ac36b9bf3b3dc11f0c03f93b518bd1f7583771559ff66aa9e502f868dc79b1f55940539afcf48db8122947911b253e50acf1f50232254a6538b41698b3261a9638514f6236a0c180ff0b58e0fed256a383469d04d2f1f6847e34eaab79edfd876ff0b15b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4ca3bf5228de05f24b07a982d6e2bca1f22e877243ef672f9e19d888f433c0b84e5c23e2fe217b8a0c09cfdb8a646439d6a59e40e691a4139fda034ad98ff91cb29e09669bd306c1e5255e60976c0031fa81db6be577b40f5910a166f967d4b1ba65a2ed4cac0ff1829ea2a612628d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20ebce1ff3a89b92a5e03cd511c63ff16101b913658f186cf47d77e65eea3aee5912eb0499ec4cab8809fa2f6e08dcb0bebd411d113d83402e90928b20ac8b028baf72cad0f8b240c3bb8f51c0d4b577e5300d381c0dee5c8c4969f67b963e35fda750a53db901a4605d87b44c97d7231;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2b78aae706646b9de16fd19dddc087b974ceed309a956b97e4ff2901c28050c2cecb25c8bde62a657c9f03a2f1f4bbc88803f7ee9aba26085fb2f21772ed53228928d87629a575a3349ba3c5a2d2501190d0626cde8dced2476e43481b1cbd18af40ad84212622b69a765f8ed74c039;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd21234449476d103b085dae5d28cf5b99e9a71349ff34343e72be55407e618eb5de230cf2f11525e4d6ad63e73c28b7526b418b8ce147688c7044aabfce27ec21fa9b85c494005d9dcf4cf9fbe0c9775e6fc7abe8353db3488daadc0951677cefb4e0c55b3dd2a831417e6ad7124cd422;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h747cd5a593fed8d2f42f496ce1ca7e3f8ea8370a7890ee07a2e253db0c724e33700aa07b15e02b6161df3997af88755ea003003fb15c10974dd4629bcdf74b8e1b115fad64384200c7a5724bef8ee3612b60bf0ffcf88dea1c38cacc33bbe84a1389477720104e7258a1f91696a62cac8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69ddd5f36358e1079d0542a1a39e01655710372b2f378e96720301a1433f3dc8fd36691aa4d913d54124d4e013ba4fd21dcbb5c90642b009e318bcc8d5559834caa5a58bb4287fe58627e8702e3353d92b225e8924e12e22a69c6c2c02e059c4c890d40d44a1d01c488e4b28a988fa46d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94b34f273e1a17dbf6a770f7ec43cb39335bb8489766af64ea48e15444840370aa439a7f711e7167e05e5795a48751c1a1523dc0b53d1a3e3dd59ef919cce20d69a0cc49f500ba74bb9fffedae25cf20ba7d9780fb8a38e19b86f0a653508ec38750e7a799df1a72f070c9217988203b2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa0781e04999c99ef276f9ddeaf47e35570282926bb31d15f9ac44128cf80889d293b25c2ad758ec875b1d823b2468266746c981214bf5a5f50362c8006876bc784d752d754784176b6490fde4862c2173517dd5d22e83bdb43ab2b2768008ca1e8a5238ad04d700243990ea7b2e6c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71cbf86456a36ac1a180701dd15a5b7aead709df663337372ba5554b53ef78d2be75a8b09b369ac56111378ab5cc06b3a93bd6f6aa77b171237884fa24110aaf4f65e37e3c75f70d12f666a69d65b51b3037a1d9ff869f2a3bf4b627361ee8f58375e2bf8bdacbc0f831079f4ee9058e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65f253db689f640b16ea8c741ac68dadb2899991bc2e59579ff2e082f593aaa6ff9bf68c6a2f85245f956a788767d49e09e544c08b43085b25c790b9d031e7d0a52a5407bdbd1c9a7eeca5df09070a902e54ca2194be8b93247c460afd1ab37898ffc42b500d0355ba2fda4f6b0aad6cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had5c026124bd028e2061765d1d5d5bc849bdbcea14dd5b2e3c1e2f4c4b3e439778a3f0aa930a50adf8e9b02a35d7e12b7362d4e4a88dcf07f695c55d174f9c8289ea583351e4b3356c891ca5e8c1711f4029c632165440030a845644d89b9529276debd3fa3261896d63e90cf78394d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde5717f42379ce34e777014ad663345f2b894a918350301a9afa670ffcd0a85604299f20616b56ad232654e486d28f63c277db2fdcf5943478b47ddd60e6645b675fb9a6e2496fdb373986678c681ff0e23bead7bdb607d933c1b99bf9dade38a523b5ffefacbb2cd6c341d82f78e678e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81ceb336520d758c9a9579390c2d88a889162a67bf03badad1c529d07cdca988ea46e055b05dcdba153973e055b36ac1c0657f881fac1189672a3e88b83793919820332074bbd750be7b9faa51f29c312d9b38d2cd18c3896212027e1661132b50a8ca50b9eb9efc7b21f51aab4aa3c19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4593212668d908c581fa3f24b847d552363c2f7f4e01fe4ec861df1fb7c632dddfc01984aead0f055c6a9a4cd918a3cde6810007120d37c2d7d74e3c027c120ea3edc1d7b5d33b9d3c752d6973ef6b0db409a7bb3e3e1d27dc7234b7505f3b3e169e1da003570fdaf3eb90631ed1c72e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9cd6b4b5e736564b0df4804b945d435c2f9dc3fa54383ae829ae61dba7a5897cc852a055bbaa20d2a98310df36293254d680dfa18dd35404d2661fa43589a47bf1d8f9de27cbb7f8c6273d2cba8ff9e9a8cb9f6be476244615f4de6a19e900ac6c1b297b88cdd1adeebb370150db67f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0835590b244ae8d5982a65e0b8f9f6802e2791a85f52a5affeb80f1c1fb341f37ded8b158d385fc4cd080cb1d22fd929d451e62f31da0181cbaa8461699a0268d71afd1e44e1c8bc89f8d0dd7a8f08398d8fefca9d3f1e401a307dbadd3fc70e4b36f3763de86f467d4804bd48be2807;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfad849aff0424c3fe6bc18854c5492157f651ef51b2039383503e695863de17e7bf40e0f7943723ded90673c3d81d47a3804be30e85836aa1fe4b66e11a5b5acb61b96e404cd30289b00662a97603ad0787b055ec7d3b647e50bba1afc4ec98f2ce3c5048ff80597d315f3f013007e6c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e8d81b6977b10d5a38db28f1e05ad8ae6b5d19ca5b627a051655a589439a5e779463851cab95cb6ee5aa349d27f78aaa0cdc1ea9d1b20c578739c46023edd1471a77500fc4e498ddbc454571ebb42cc960a79f3b165585e9fb8f74193f464e252e3a96d7656917c51f5007b138cb9290;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he313e72cba1d554b78bd0d2306227d718d3e34651c78ca0cedddfb9be35d1d1c6f41813cc0e3ac0b7a4448ae792910031be6ff4fd342b09401302feac92701ba2f165eef95e20372c2fc01e7cb99e9e1232804037f446456bd817c6a2e229d9d68e89dcf72436a8c41ae29b3c9568025e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecae2e223027e11fb9ce824ef725f12f5a0cc022b87e66012b0b75af037d02557a9e5efd4a7536287b255c1c2fe1dd8d83a8d3bf4ef3a01800ad4b280f967e9231ad2524b26b22fd325c9fe8519b1b67aaf5728b2aac536e5084743feffaf33be75c1de93ea4358831725d7760582fd6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h425e6537876be7c969a81b73f4d46017509652c5267742825a179bdc64c70f4003672a0b5d0a1e5a78441e895b92f0b9a9703346c6e2ae76be45ef71e38996c65d26a548de4c60e9de1097049f96895a72033c830d73a576942b8de4359b2f93bc71360a503ecc28924b6b0d75df256b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h421d779a1ba953583804bf636637161f873f52958968f07f3787d138c41a2c602597a4e80bb60f4f4445bc8a7276ccab0b349416ef1332c310d578575777bf2b34513acbfdb6e50b0b5bf7e6776260b67bf33d333856812553145d094d04313eda5dd2d1fd189d703b1cd4e5328d42d70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0b61242ea4228ef77e19c64533b52c155ef45c77dbd45d405d7cc1ef33f49c3c306f97ead5b43b4c0ae744c23f9ccf19524d51ecf3d3dbe3e5fecf35f0335285ffed9397ebda432ab770b4eddd9b0ef45949e34a301de7957c229aa27823200323b58de818e3a33dde97fa46d02fcaf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd08ba33df352baf236a27bc04b4fa338bf888d0670192b496d5c76ea2bb1d4cf2f2c21d451e114cf9326595323b8c5beeacdd3eced0d90d81b3df37c8af18e8d62957e053340aaebfda96a813b80cd688f9d37fcb8959b77f22c162773a69c5b4171ad30b1789a3e4cb48712bf9a7c0fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbff1159a1ac554263ecb125804b9823e5f9ed3b4ec7e3f3c6ef6e674bb81ba49449f58e6566b26b1796181c7f64be1d9f188a6a757a9b5acdac80246f062c9fbcd823933be587041b9999cd1acc86c9ea0bb7361d95531b1c62f9af5428a8fba7e951a313f1fe86d5d5eb2f18c8ff15bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40fd87caf2ef3269d3a3c5e3e5ac8d29ba701438045d6401ff6796f5a9e7f83303046e01e861e17378b52bf9b5c069c656186f294e84775eeb29fe3f418b53dd9bd5c8af36b846e66f9e65f6f56067347d72e335aef7923a4ea3ca537fd20094a9d068b16fa575c6dff596ccebbcab4be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53553493d5af98aa8323846ba196d8de177cb58ea4ea7b6d44907c55c885b649f82bf4709a3e8b41b6f24ee9a95ba86c20ffe011c77b4441ba34a548210274379ec8eed3120a5170e5f4eca2c72c942afcbdc13278c8e254a87d5fa9b7a37992f99cbfa79b02727063af9e398d1d8305f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd30bf6b9da4f6dd24e2f2ba1532111e08b48637fc435b8a8a8aeac607ca1c93a676e1aa2411cef161cddee326a34ce51c234a87550d2c4d3fdb91cee00197216db4cb99afb5378af0609c4a0a3fec0851640518c7b466e398245944ca4370350424433e8c72391dad0b0f4011cc4cb14f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18ae54a94b7c7740d358020afd5dd1c1ff082e17de7618e4d33854b5c5b3f8adbf188b255a0d791634b8ccf8c02660d0f99ec1edecbaf8cb765c3ca413dd684bfe14de1c715d5d927930af76dcb57d5cca7942a74321bd418da6698e839487f54e728e8392b006e59515378a8f7994d16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d39bd48095dc54e2f498aef73051ab3c869aa9053facb4050027910c61d49df38fdd3e8acead85f479ccb0359083ed79b1d44278919fe7391ab0f5babdef439f2a88acef55f10c366919ad643645c0b3755bf0cfcf37200b0f651bf4d168471439067d5bc02154da9d76d7f2991de15e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde89f6717abfea2ff272a5019ea8729d1ee39835d518b6aedd728fabc8954f6b119ac57d43a5e3e4fdf9a401757a762c1ff0afd287dcb15f38737985eac98369d60dac4a35b49ae0e118fbf85f5ddc3a80f54a7f528937cb0c816e60dac59b59d266f6a27b3be8db10bb0d518794d5d18;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5929f26bfcc926a0929442bc2b22ed544d09440d76f4d0e37ef45ed2075e826516a005820e22dc558083cdf96eb25f26de21a0288266c974573f0fc377438f3a33709ea05b16adac017eb1557a5b8d9f67f661f4f12c3e09696256ceb427eec0392238e0bb137f3d6521451739f676ac9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49416a632a1832a87f53363eb79449d8cfd8c418cf1e7914e7d595449e923100701d7642a5b589a02d97088c65a8222eff37d41caa84e35d8c8e0f3ed08d2250fa07c6424855b47ad0e237a515b132c91f5d5236e081b227ea9865a698e6ac17fe7d547a23a9f4fe18ed63c5deac85202;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac7a23e701326d9262a6cd097c67e8076a250b319411c5cb8480194b0d874ce0c7cef366c59976ec0a4a5e3f6d19ae122594966fb9a740a81766f2386f0da51b3fcbb52489dd2dadf8dabe946847ef972ef7b74e0f06b4a0e3d64cfbe9f256c072855eb3fe655189323604fc1206f3e3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cb91ba4f62646e0e6a68dc0d0d1eccfd567107117fe42d8c21d22add4b4e076f43173dfb21cfd0ccbaac1bbfba9bb4cb0cf2791cc5def58db8fc7489ad678b2d631c425b06acc458d3beea0967e76f6e533973ee81be6be5672a5044c44b761625e1cd623d6f75ea08bf663dc1acab8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ffcca42f60f28a959c66b71055f7f8529b8d94b986e5c948bd01ebb4c9f7a85f9ae269f0314a8047e9fc0c8edaf09537f15be604402e1f0c001a9b38d8b9ba1d93e66feb3133cf766ba28f2d7c5c7a06e42736ca15dff1b3c9e81f5110b64ff97efb43c4788265e3f32f4e21253a0dca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f4f2d261fbf06b74c409603d099941dfb144f710285793c0d1a9135b3eeb6aafb68aa615e999f8bfdac381e69e1dbc6e585af9de7fcb08a305663f6a4fff4e2227e6f370f596567c5ae852859b8ef3b146a5f748d290bb5e57bd2f8658cbe46e0927ee57a542f313ce235724471b29a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84274fda380fa8182b9690a605473462f83d4a93942eac50832a9528fc6b68083f62ee79860447762e3314ec386c27a3d13cf071deb4e2455dfc5abf183c7aeaf7a8284fad127196b150ca7f15fc59d828931e361f6838d91b2bece20e13c5573c50984a75a75f3508c866e179e7f7c16;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93f44acb4624357f4deb035402b3f1c0b5528e25307a9899d91e9ad4d358e0efe45f05ecb88e3a100c73658aa25fc8e03d9263586784d969ab0ac4264f5846dca2f81152fedddb68d4f0343c81289097a0da3145ad202026170d097d21b82c3d6de80b9fd571281da79b885e5cde43f66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c8677b60bd683b3c7bab805f17823ae8e62e4cb47bf5666c1b1e16c75fc38f004a8bef2afb2e49c0f39f910bcb1d23fa7872253eb3f5f67bb0d2ed4dac2665565ca8c0f40078319f8732c4cc494294583ca9d6702086db5911e648e5979b2c47bee4e80686332f906ced54d61ff46d79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4de7861fd4e91d987adbb04d3730205927045f95b31dc3c39004465791d73bc81b4390da91ffaa4f553c68c20dbe59e6897f457d4fa96dc258da0f11f94297bb0c4495a4fac57f82e898e4daa361a9cbe0b7fc9584f96c4faa63235431bcbb2fae23f5868d1b59e7416bea02b69799211;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61d8b4c5df97fc072ba1364847c57f1dc84662d39caff66e36d96bbe3e77c3bab38b8b5e8895190abab59900d2cf4b1dac3eaf4eb7ec031d6bef7448559b3e79ccf73e2719f7b50a3c16b15e69fe6d9375f0b74c214a4362b869949867f78cef4cdbbe1cf96b106b5b4a3a836f196b9f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82412ca1551d9d0895cd0bfdd6eaa0ca5ccb433f99b26b85776d439abfe230c26b19fdc799088f12f1d8d3843eeb26c3e718b7e468f643ba1b2e276a7033809d749f205830aa8b4e5190bf3c674fc850b8a5b89dd6b0226568fdc017d0363a67ac2016f4465cfb6b0e697c125a989b8b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b000f90b1925070fef633c7f6a00cd0278ddd8a36b28dab6412e21e6c6ac81c41c5511652209f3ba91b15c35dcc4597521331a8ee3a627e9aa3bfbb6cfaa1fcfb4c65b6a258687e6e118627d48bacdbd1518c04d032e2cc1a109607933cc00ff951ec395e6dfd2fab068a8790f57f1cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacdf9ded66b5050042a370db93ba8ef6fdfcba323666f3905bbaa2492a32a90df9511f0259764e6c7cee70d7a6dabdfd093d1b2fe4ecd48d9f24a4cc5e050a5c892fcf0c16adf6c2fccd25dd9c1126c348b6bf6552685db6126677bec03183dc9bc5c8a952e020fa3c07154ce163ed59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf979825922d25e33c8fb39c499ff7a83d66c9f496254e1582bc86e84a85a070b0f46515f9b27b87fd79c845625fb112caf3386063b5bd0d6ccfd35512a782262aa3bd895b6394942ff6e004fd8cd4472139317e0063f7d3208e6ab4a892928a9afcc2840ca8fc08d9e3ee05419606308d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e20d18db08e4e4d4f737ab6459adc832967096a2b90bd7f9500349d960013eb6bd8e88668dc34b333fa54c2726924ee68ea72d9426d0f240e08a903afcd427319306144ac8c272a10fcd8eb78c622266a186a7998d7ffa277bdb2a7d48baafe2d8cad3aa68c2fd8df1467a1eb4b59a21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98a424c8ff65987ed93f9d7f6c05dfed87042aa7ca932288338dd592aad9e183f828a63ca46d583aaaad10d4c29db9f21d068b6f2f0b162a8a71a069cc01bd58c01a960dc2279cc1cd362d58f849e78e893f8fabe7804b8f71c31130232c039ceecc5981fc928065ef29ae8a43b20c52f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d4c79310a3049f80365080b0a78eefe49ce0a955c67aa905a758ba1148f4a2817a47fcc8b5a402141192ee7ec4e64b582e3e14e24d7e8bde131bae4b706b019c9594412c96df8812837cddf54325f4e42d52b92637785c91a95fa69368235b0fe4593e780c88b26fa866f2646713dd98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4751d81a6fb56bd7c5d4c5f34e4e57cf37941975415e5de72ab3eb902bf793a898f4d3e2de330e2233322e38c0941e59df20a9aa3a61b25c9c48f12cd3f1c27b50ebe5ea71855ce73c1586015bcffcff99e08770dec652e4f82b577ae6153737401351cf733c033b58aa92f53bca31bbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc77e9cb179d430f0ba0ca4099bd80d4c64a2779e2bf08f1fc2f5b9a298f13cc6b5fcdd1c3ae9ffd24dbc9f57c8ab65d6b246d4f05b2256296d10f7eca2503b0568a0cec56293cf6eeda912556ab41369d0fea210aafcaf90c37bbe7993a790a8789543f51ed44fb71e3fc3e390dfd2f4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc500a58424ff3feb257a5dbb1b92feb72ada7b39da83c78e690f20a206dc39b3c0d234766aa6eacc1ad1a198468b9d5cc2691383d4b67bc762b28e13d674778a1466f1d63ef15793c44302c75e9cb39a1a653bbb6623e24fb861614e4e4e39c5de8b401f74d7753c953ea30c145dd9e74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d4cf1c0be8cbb91bdd4c9b843e3ab3d2bb67fa1d57a07e9c397d7b491f43dba7c5c755c18cb39643a41f748f050f175f0aa67a74009296b219965edd0ba0387349c042e7425443cca1650fd614eb4f942c2f7c428a248406eaa0b213c54631f4c0df0a957309ac691e52ccdbc90b0694;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96594a1435d861776940e2717843c8651dafa063f45f59ed9a7e71c33aad55e34bfaddad8f3de503b1eb9ba178d614bfe8045ead8f887037990c2ca8047a2444ffc86f7d98b212eb722f831241a251605f985d926d4cf87a2ebce6e58628e7a9ebb0014605006f5dede0c38fb23fa8ebb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h999b49744e6440e6087b66d45694de3b592f7a042c00104ae12c285cd2aa6d2acf4ce14c5b116c8f8fbcef053fe5c869bad8d63d8364f80257c5146e38f7a0fbd9258090faf67347709c9c828d1c84d1d0f0530dabd10b20204adec0aeae33928bbe3e7a47ea9a6e52557a14ea3b0c362;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb06386e0e97a2fe8a147557fe31d98cc223b56c74b880161458176b718969beb81b832b705c21cdc3efb29f59d74b6d056bec2c4a543ad9f0bb2355f1e8d315ccae0c2d1be65c4bd55691d9a2f57769383b4e758b9c53e5d03a76c5c1c6af75eb7b9b650dfda9c4c0eba7cd8e872ee6f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1794b90811749061bae1cde3e0de6151895addc1c84ec192d0f11d501ed51caab3223772dceb8c6a838171bc6a604ae4456c3131d95f3015ae544d843ca0d72c76e1c10f83bbde1feebfbfb9cf445c0706fb12bdc1c01f0c75e95918bc70121d89ae8992af044299031235dd451398f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf86a7ce97d810d757430ec95bf9745a38064b412a11145db429a846624549ec89c3385da111114e7e5a4d8ac58b5f12bf0725ad7a777b075f2a1eb825de32af76c2a4aba0251fb05f234908af43b462cafa979e37ecce7faa74e8a99ffeffa41eb3994223865d8b98332f0f0610a93ad8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h485c04600e614a2d597ee298b2f0028a9c353e5b7e1e66268526a8efe4e9230ddf9af64c76cafa8a690e5b524eae652956e064c5fcf0732faf0d799a763ee6f78c8db4e4db473d3e0ecb682330faf59024ba0c3812fb2d07bed95e0e93deaa6c5f09aae24bbd91a9c0483439f3acf84d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ad262a1f6ebfce4ed1771facba01e46af5585b1da4ff196f70d327df3b0fbc6b8aa6ca3b4e3c0ce814149c6d908cfa3e1ebf61c9cfde5c42656dff1ba1bc29cab1f3fd505d4e0bac881d382928db8df974db91d5bbbcbd255d7fc73f15614b3646cfc4bcfb79152a4c55e1066ec83e6b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7beef63892e00047682da4c6e8b34cd19902bb6ffe42588d3f21f9e82c1a4344f7466892e2b411efcf5c66288ba0d3e2402dd8a5aa4892d13fcf5fe35aa339687c665c2c345f27b596aac56f9801bdfe828195f1a12b21da7cb2fe022402d25c794509118d8916646fb1941798521f7ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3de085808a504b944577ac13e774dbcb31a0ebeeb56b8a75c6bae1e27cc14893980755b503715e6583dbcf390c91be785ffdea0df9f16cb516d35c3c836f09b667fad7b235b3f5a68e62ac96fbd4bde3c71d8d4d50c82115973f0afa1926ad938fc5bbc0f72a7e0562fd89be150cd2925;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17efe1f11e1ab311926ad6bb85d49c2371a25e090dfcae1dd11f46cb0117a6eef4cb6c832ce9678a477268d4195d9b321fc2c72bef872a606f252beee6b9e7de10772cf1deb2e99eac9cabf79c0c229adffc9ef8543d64696cf78ff9858ced322387116c5d63731dbf4a0a988486cd048;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h418b3a9109c8eceb948d1eb46f89649f781ab74e9d3871f815ac1fa1f404c8a15fe6b7594a47c530f4cbb8fc011e42acadd0e71c319d8b34cbc01f8f689556b670b050d68ca200311409bacc1e21c1933d2fc47bd2d22e18f89953aa34288b0ab35bb0996d3eb263f19029f22471ee4f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd180c4f7d7431749fe90f2ac97e9f741df41f987a8bb823d8d7e1f4c11a70fb1ee20545d23190c1dda1db714b05cdbfd2c92ebe3ee4ada3b14529504e0e66bd8eb264872092207e7b385d75f133bc27dad4d88345b50cbc198e8354011a5026ebba4c42dd2e760739d804eba8f5839ec6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59083b8fc598869a6fdefd66ee9dfd380b92bde3e630edc1c352e560f40c9cd378136c0196ae87f8e0a75538869f748ceead9539a4438f89401d3c127c64871082b52b5435dc118a02e7d906a93d1d340b1003f6eb15e9e683575914d4a397c1403a5b7eb79f2b58e67b6218b6acde8dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4bbe2adc64115be81a4318ea267c90d075959af6fa6fc323fd620fba4d1b01d3d66ba4536f2674a3327816650ac0f444791de23d16f2e3659ed11dfd62666c2a6a55d63059c7253c7d4db975bde2ffdc2d3a0bac4a5e07c98eef59cab8c7f76a312c0d952b5644ec9357660640689556;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b31c3442b51ee5d5faaa52c88142bfef9e8ef74c3a0138947d0c91eb8a21a4ef2cc43785c19b545546bac3c4c96ae603d5494e40c89a33c9470deb4a3c9173e67906e3020af58599f0a411c4c9cffbefcf6253c03942ba73d2b959e1ec3974ee7afed106d4733ae96554bb7b106104c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31f3a9acca6e05657bdb774ab63b4184c6ebb5d15734ca83d8e4531ad12e2de0534d925c1de0833d172d6511c037498c34043ceaccfacacf0e222e22c48850e15c66defaa9284662b3fa3bcfd6743036f332b3e63fa0edb4f3eed516bd8bec9d872c7ef2a5b31221b4e66b1c490a5c9cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3904088c6febba8af760169ff2daaf9e72af1d32daf36f1c10a0802bdffa7ff018813791008d015692e183acc877f75b3e0d5928d9767769571637d9e7faea34bab5c06870d578174dcdffd97ba0865708980fae906b097eb51d803c7de5af042a7aa7dc1832a0ca0f701b11c61a4121c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8ec8df6add7a06e1e2a3a40ebf75fde1951331c4a68b72245a233532002859d7ba2016054c526b7cf495172dd2720ac3392238c81eafd14d9ff43c04f243493dee3b1c5a3f14fb732949e7f98e589583fa4defd1160c3a6bcd35aa2da89ac3771ba3aa98da7bedd7e7ee79d82fa47e48;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98a4afb78fafc8e4459e899a3832a07dcd7e6872c41e66881d77138f3f63bacae148b165beeb4f25dc2ac4f3ecd37ea19899d089f978e316edfe2ed7a7a67ec3b310cf28e46b63b8d0cabfc0fdd326e057177060fb8e2ddf7b398a77196d38b85ca7a7767d1fe2007f97867bcf5fb2fe3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b46a9c1c4dc577e8b857bdfeb6a288b58b338952fdf4240885f1b11dd63c020c0cbbf2bbc00348149cda1d97ba558c187d86e28a8e9714d82410aed74f800b629fb30d42cc5624115cee55d51bc6dfb037e148ad1ee61cbd2f0c6d54303eefd3ee0e574fae9cd8f3e56796db2063fc7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fe2888a8e1d0407a40254b2b4cc543368b02db1bba77586ee2bbb4cb286918e949a8dd6b5485601b8c80d159d9212bcbf93bab3eeff83608cfb3db54de0b21ea160d64b70150aa7a793ce37084fd96a6db752fed4f6a674f2f4b18497a3751ad2626644d68e478c9bb3c228fea1f6224;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h219a91e8f2cdc29bf5c16c2b8de19d940ddcc36be0319cb58499e447520704b109239dd0a213079a94e897c3ad0b7ca9c52d429ab0b24c9164b701571901c225961d811a25e9ac32588400acce9c49a7958e63028ea0b47b3511cd6ced6e4e64bc4bf84a7fc2270c263ecace4e9e85e23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8041447529bf9b793b68528c46eef208d324545d19c40f32427b876c6fcd304fc58dcfec7c6e4722ea2b5171f8a712f950c73444f22b3c2bd34c243d4ff7cb503fec998d41da13d99bf405f1e9ff7dea6019bdb50f0bc19e814413767eb0bc6c501a43bef444c0be5309aa1ea4cd9dff7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c5f115f890658d5379cd29708d14ba7d6a58bdc1c1a2dca02d10e07bb91452a3eb1185ee694d40294291d1cee156f1ba7174b1140e6739dc62bc9b920200e071bcc8e9f312ca5b616c050555809b7b586bb469375c0631ca077f68c9072284ce70a382b700761ab8f97cf65f512e2109;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb959a1fb817c8f7b20d5049b0159f3d60d1bea20755730df7ceeb554687a4dc579f0a45df1bb4b3acf4ef08c1381867a1b9c020252865e6ea8f332459dccd07712eb6c2b48a8ba86370b69280dbcf46f0cfb1d9b7c23731d7b2fb4a1df54566f3811a40078df1ced93c7ee74924205496;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27e8b92ec4bcf4e25515ba2481c9a17b5d53ca1180e17bead00de1a8bbd5be5f9981c2bca8075e3d00185ea4148734760c251ee7b2fc60d5eb9223f473c89afacff35d7357d758b370feb51e6932597dff8adc183cd80b43e4588c29933a208611bcc6e8e9afda9ea52b081c3f86eb1b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26aa52db3c28afd5326b86b67b3de02104348b0c3ac721ea372bcd369a0a31e69b775fa2cfb4f62a6698dff137c84e3d39d8a4f5c1b129c6aacd80706911cb29011ac83a6236e88bcda3ed8af423dcdeb2c195e9f556fb32904b3dd2059aa9eed198f20f7fd1c6e85d602f994c1242da4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb24a8bff8d95ca213b31deaa659ea7ce3f5f00e61efe329284d4b637af2d44b01f5f8c12fed73adec52a1eb00a0268d9bee878db7e05791840ebfd892cfbc3c84c9cf72459f94f30bb6690fa5bd4ce6be8152ed1d048086b72989bc9943622dfba1296b6d90c9eeb963d17b490326054a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2be28a8fbfc2df24e0a6a49d195aa8056717703ff9fd76bfd2f19d2b6b31a694470b0c65462d197c331261f90c94cdaf54f46ef08e39be2d56e5dfa64f5ab244b7f1796e363644e68e801025aa32ada40d3054a3a175cac42633468a48ec7dbf6000d10ed131106ab771f6560028d90bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb419692390329e53a0f0701ca80ca9a8d7af7dab1f6fb141ee1d10613833d6c1feb895ea7093f02537fce7f1d4c0deab542309f8217addc0f02a67bde00fd6b19b1b295689f0f04ace9fd7447b92b6ec63324b79c50ea90d1165ee86e9bd3d794208832145609597d2ea7c6ffec24e04;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h851d7f3825c513086d3a2fad4103ff0b215441759cce9e70db38ac97926e5100d6ec599f3869ca31a349567917f1ede8718c43ff020d13d83516941e137b75437318d67911865f62431746eae21e193b845bda316452ce7a39e5bedb863ad07967398121290654cc015f92b0e49c09fce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6e8610d35e55800c3f0c176ac985af863531e041abe3c873b66819839fd1ac0db9938b1b36caa21504a4c810593d19db68b89dd058a8665f85adfaca9c6574cb5dfe95048f50195c4056f2bd08b68695aba30570e9624503e8a2b772553fc6ac7f40bc5ade552a29a6d6e9b88358d0cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8708eed836385f608ae1f62b1cb42b1b3a615e7a5b434bd41533f9eba38dc2eebaedc0a8c5c1b4bbcac0fc0f3a6a348ae806f9918a61342816d2e71bfae813edb2a0196190aa83d447d2f98d8800743fd556117412d99dd51e34cf6bef4bfdd8a5f08109247b6c4c0d81e1e6490179a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a24cbc19f5da957803c8f4f0d1f7da02c37358c4a856c7afe4de552b5c01a5c5c9668dc01232d1cd8542a0629744640e70a8ebb2c6d9f377d6d9e704e4671b6fdb4dbe2482f37716ed92c5ede0f8d4dce039f28a203a508e30fcbec5089f420f60c03771a2231f345b8e5795819e68c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18cfd09b70e0e7d525eada90d30be5eb208b6017e2fc365f0b8e78246767abba66d2825be6b94b3768dfeb4fcb4b144c95303ee833d2d76812c49e58efbf1dabd689bd7c1e575f19eb090ddb0f6ce823da7d7d9ec1dbcf96df8ebed4a65770fcb893ea6fe6fd7f1a6eba86afb0e3359b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc51b03bbd2ed6d9039a74982aa74c96fa6ef74a8ad771d710fbafdcecfeb5e1dbebe27e9e9fc41fa578984a9b4e1ebd8c32640eb4fa1a92fabf9f7bb4bf8e77a9a7625250aeaaef182ae3d1979a76a06d676ce2b11b43a570609f7d680b3391f436886f4096806f3116c6254cec4f5e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0d4a2faa234a8402931ae17cd49cec5bc0e65827e28e2804825432c6dbca2117ead90c2817275f32dc21081740c2a24f38ea549efd81cbf469ca9dc516c5af31ee84ce8c77f7272e9ecdd4a4081cf403ce2a49e261c3ae8fb839386d02defa5ebf774726c25fb26f967b6e94a2cd15a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf35f9d32db13e34411c6d88bc7ca57f797dc68189c7fec78e04ea47b8c40cdff1bf8afbd242f2e86e87b3af5549aff35fda20320e6a4027f6da3bc2872a7bc9c252db1bcb3d7ff3011a70c8d40dad7b7bb4594cbd240a74e2c88d891e2428756ca24ca19e0056e2c811097e35cd87772c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3906043bbf4f6953000c9d20e4bdd8bc6edd580e8391850be3ed10c6c081eb9f06be8e2d34910a5e8e04e735f8fce24bdc27142c1e58b427ff2b5b1d2698db8f7aa441b6009a0efd1b9fe13ba6a8f132011576c0ce359f8d7c4656a54239f7eca0924633332a5d3a11904ce70ed1c09bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34dadd609ba5c4e25f2994af159f1c7d65f64b5fe7ffcedda6a0c088f61bef4e89162643e2398765c79c78629496290ba3acc189c1f06a325ce363061dc364cf7f4dc6c351246f49fead99fef0927ed14858172e0ca5354dd0f1038871a57bf520b2f19963641ab8a53c6a251f43ca177;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dbc2104982bd7baabb8d244fba3be3893bc3c08c6be9c1ab466c55346e95cee4b792b0dd57d9b4a71c20dc6133a90732b082c0d6f1d788341373e48f02ee0945f8805e691e66577e8be9bfb06bfe8a209002ba3a798173138441a0a53c9ebfd717f9ab06b448a37a45983c740176a77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5a88cbb02ed1336489dce293460e9c6f81ae44819ba143ae5a59fd54f6852c229c858015b88901eb150ec27772606c8d53cebb47350a853ec15d4231a01addcdc9f3240159d1ada5aacae0ca78063645086a069de6ca00c2b6ade5664eedd91b58e622376634e07c2035454de6c5ce2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfced0ab171e4de41ad8cad6469e210c75afa14c3fe89b37c5422083f1263e4e71c2508dd8b7014d543b9d111d70637d56c9ffa7a1734fc06b3fe82115fdaeb2174bbd90f3d38508656dcb496bbe12f7fc77f3b66fb27c9eae2b29b902975a544d9fac6cc9b808a2e193d7a38039fcd74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b6e36ccd7134f0d2fe68a86cc67f89e5486fdf71a84192a97bc39f6933deb713b04ba9676e0d4926e371c488e22b69993c73f1fac9995ab6df0b19625a4b051afc1e5b63d144becae48c65f6690c878e730bf8e6b1d81369d2a30304f44292f343942df3f13513be824fe61c7f0cfac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ce5770a3f625f49dc7b84284b48e940499bd6f9c12045a5b0d4ba7a2232672de41dba421cbb338df40115088ba371f16f7a4ac55d10679752b4f3897742d8a238e751f97f6a2aacba73a07f3730cf77f1e9ff64b4b61e9f94512234eedfb2d33a96819184a0d0e84c2f2b70e9d7d2a18;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf41dc67ca28c83e03ebc091a3121c522a629fd120fcd0f5bb308ebc500b37a65ab793156c1e72fee40029e7f2a41053f109909195e2bc72abd20c0b684e81b73ce2916d132e0379850b050a89cad3b2b841a5790ccba89346009a0ae0840483fb4e1c59a8bd3722245f1432b835c1de48;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50a0696688ae4d25e33045d426ac827e5506546d3efdc0080fe2c2369b7d3a9f4eeace5695e9abff8e2042885147879fb5a31486d60ecb24ab60bfe9194515d7ed28874ad4e5016472de76ed0d42504a92ae65e6edaeef086c34a557a8b8fbedce5c9d83d0b208bc035a8e905eae03d85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19a4eaf9825e8820438df5b438ff410e3f7805f4f2316224b9f7e938655cdf96c92b891f07da1938888ad7ae13658f6d8c3094e3aa00107512d63eab9efe1790a38e5852a7e456187d2f9e2c72713164b35ef8ac0d119aa8498ab52909557c382b0c464cdcea71c56710b049c0dbb2e06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc05bb28c703cd91a781b5916b8cc316011520a90a6c0835752beeeeb3f61f081d39ff0786666da2928a8e8cf6e5622ccfbae5d455010ef23bc1e90832c4fc1c9db6abd928fb587e2691759ac506b7673dc6dd9263cbdd8eff86d8400749441422a0907e83dc79da76d258cbcc35e883eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h422dbd34c26afe073c93f4c9444748f3f9162e20cc9fe9c94dc884e5021cbc756c358bc9de63569b634c39f16bdd4d3a777837f2e09f0b20f5b2b29baeea4c29881637f953cdf67a1ce6587dbcb0fcf65c81400a1dc551d976a5e8d4654e9c26fa43f4724c63587573435faae83fe3e1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc6fc7d4fc2d5f8c0d4096c2597ad8e187e160f60b2e8d9e9b6bf05170f612beff2c6077dcd7f77fb16d837d7ca5d8020ef4cec14be3c90720674ac10f50baddca2344b4d174e3c480c49065f56acfb7e632ccbe80df674b01d219bbca65322d3e8185e57639a5723b631d7d3fc7f972f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b95858057f41382b40763af363ffeef17e3b9bd9c7a4c82b7b8e597dc356c16b26191cd818c3b26b2425e9b0047510a4e4882f510c17613b5330489628b94d174b76635ba2504a7f5e291cf2bb8631e37d91e3fc29148e84c50e93e8ec3205b3f266ca22339a1a738fde46eb28f194c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef965b3bca18ec9aa20766096bbb6a20f53ee4cda1cab6a659ab2ea5a37e0eb2681a73d709b57a703b7ca28a6d4cc71c14e9730c7ee3ac081c3a41cc5c195a7dea11e0ac3606584fd523e68422fdf3e4eaf046c5b6b84051672513912b8cbe942a4aff4bf3bd51c645294cb1485ac0c06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1600d4fbcaa06db6dfa3eb79ac12746a4883dc229480fdd00fab796f7a15f744efeca34260f92bdba8410ad090d1d78e9c40d2c839bb45eba9c93612676861c38c9e8f4408062125f53e352440681eda965d6c592deb7d5162167f600f11a1ac9f3465ee57c5de7b26599d693abf7381;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d5b9f352deba8e306e7f47811b0d732ef693f560bf69307e2a535dc892db7db985e32a7be3f575997944bd1673bd1819c5aea6f6ebcc2faa200d03e9d542a8e7565048b70753800965abaf7f05025653dcebeabd603bbc4c6fb2c36cb44f71ea2c72aa8fb3842f98670b598f99369ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39239aab3cbabe5c5af72b0505a1b5d7088a03bad81561d4255eebefe503beb43628c1035c9f615de804456ac5f82259ea95618c6e51ec8397368debde8c1a207fb71a19885a104f5fd94afc586cec180fe0ef2f1ccfa96153d9cf12297bf7efc94e0c23e7da378512d34ec9a220e2d24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30e7e1cac1a4adcaaf574fb851df8b544f26fd206d88288bf024d6da3e9aa0b63b787eb5d2bb372f2d2076cc9d44c77d253f20506f7dfd857375f240f47b063f54890b29c141031eac7200a91758556b190d869654909aa207a9ad8d77a0d43f963287c0ae1001b6cea571ab8ba23aa22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0c74acfef3eb648fe8122e20d71de9bb1687ae3a54abe03753b7a483a5c04a385631a54be221700101708d891d31bd443da933431e68dc5f76bf207082cab614835c87ac1678b7b2688eb03465cc40e03515803b58406bae40317d66d2cbe48e77dcfa8f102f39e57d4e03526238034b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceff2a55f4e01ea4b3cdca04f43da8907fbc8ecc705bc6562a4a8868374de9e38b879b1be44eaeeee8b1ea2d7225cca2b532731cc566be99065d2754ec2bd63b9883cf6a59552495e4e4bd1a7d30469cd576cbe07e9cfd7031c5d0485487b7f8c5ddc9102d2af544100986b42decb4b93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0f9a9dfe61f1d15b209a45634cdae37d20faa438d3af209e7965133a26f0c010e4542b769ac9f8e1dc26a8ca5e86b22ec5d66cff3cbbd507f04bd3c7fe514a9a08a46507c26dccc37a3532df88d980b6052649252be844ae258a35374f032a71ca42be9024ccf5a8f494a9b67b86cd6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29866a2418406258cc7dd9389f30f184a3342477d2e60e4ae4d4f86917eeee86a251e464d494fa2ff3da612cc15b3740453da15a09210115c7234d0c61211fa5107d548d44d73d6f69b3e875d6e7e46f7771691edb7dc42bd14d43dea7fc481c9ed1b44e8088c24522612cb36362608d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h317e779aaafc3bf599a6fc6c88634009eeadf7a9c1beffbe19098fe30e8416f1d4b4aca5a72cf3b1afecf5db4227235a08d5c10a82f9cef0599eccd431a83eff6929f6a7cd642fda91eaab7223dc0c86e52a11c9726017cb51b0343d6ec56d568ae38c3086ac81f66d9a526d002759d56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5fd49821589cf76c95786c1d2613e4876bf13d0a77eb4040ca15987c2366015ae069d895facda6934a0ab4c821c71ece62264682559a4b4ff4cecc1aeacc406dd43ead1afa13f3792a1d2fe57abffce8d288a9ea38b1dbd02a270906a960d5f7a54a276770c7e1a1972f62ff5741487e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he44f3e65fb78b21966046453a4b38b0e32e914f62681fa78f65d9ba6580ce7b732d0166bdd1bc8dd100ba5d8e0f9c9072dedb0d5ecfdf3fdb2a052ebd289577b341f165d4a9a64ad364d9b066745afae0dd6028ed1db86c6db3eee44fcc02589ea9283dfc17c47f5888ecff0cab88a117;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84293c70e77632f1faccb6d76f8e4f55667a08de7f1d536270b98767f34271a46aa45cd6071eb518f53544484f76c9e6eca4ecf903386a3289dc34170d8af14bcdba87295f94ee29e7c3065aadc62c723343eed7712ccdd2d300ddf709c061ce4c6bf3dbdb9967b46ae4569524785f3f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b1659f86f96b00542cc4fc5296b0f9f232b6ea02715da3e8284c2bcac59c53051c659350789e05544c90f155044dcbca118739938b5d72a7a0aca0705aed0f96c9300e512a32822fc39a5f87c1b9634cc17cc29402c03f29119ef9213373d677375bcf32969c72843c771dcf1852fb8c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29c0fcb92a5e1e71dc46045347f02c78d16846e5069f5220f63db3d4a0e3a65ff3a376a3964b4c08c0e71497e3a9fc8c02e748f4a3e0592eddf58b472bf94e675ea6a2b310dd3eff9f2ba01c22914aa5548c57f5741ecfad9d5f9f56dde7929e832daf816c8e293324fcf16e285e631c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f237c51f9d3bdd3cf19beda76a72b54fc201927e0d7634dc48e4fb6e63495140dd7a1ffdba984c07a61de62b4ed0b73d4591d8e15cb3ae0fc30764c49c7f9d101fc7f35a85fb25f2f16c4be9d427cbc29e4cab06dbd4660865f04b5759094d2f6dee6518d0be3700bac0f39153dd0f44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h806a7b935cd13300037eddc78df74795df4314b5131fdfb8bd64646add3583fe9a4b41e095cb93f18e53b47db67afb69348b6ea9c60636868e37976a830b65d2c9dbee2c815d156acb0f088ddd12e09acb79112a7afe2bd823de9cca88dc0acc507ada5c65102069caefcea2b0f501fb3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefb82f39672487f75529ec621323302efe6f116f5a1814a57a2de9199b1bdcaf48fc6759ecc71f2c7b87e4689b7c554be6a26c1bd2c3ba0dbe079b5cb67499ddd564eafa6a3fa8be2a03ab777b1b6ee598cd7d329367fb80381527965b2a67cf4d13af8b18dfe4d8ea921b51a90b91d76;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb54ab748bf767e4ff656bb5e81c0937dcd529f8e9a02e8a8cba5aaf04f59a57050795331dcf5027cad930ac7af83a2ed3a029d2f952245c225b731ceaa21cad11696e9acfa313fdda866156a73cce0af67e0c2a0e8345a5071dce71a45e9ac64eac452e1087f4b9b650bd212a9b54ae0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd90afae36036e4e611efa375e0ee3a9deda8740973c8831121f4fcdeb4104c0544d67fa31abe29a86f9de09837f8fd1278b4b4055a5bee125f641faa91476eeee65676310e53afb8ccf140a144f6bf299990e98571d310718958e7c9e7bf833cb9f801482983044cb893e7767aeedf2e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b01ad225216eb1821a3d47ffa56fbfce9dda8b4d2f73de6fe76de35d4532cbbd9943da5045a14c6a397a169fb6b0751827d54ae6c4cf01bdf6709b8f544ae4c11742943feb1902315c11613a62244263d647adcbbc80f036d6fe55d3a02361fee38bf3b492d66aeb8832cf7ac4d657ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d1a355985e153d4e931d1e4d30cfd203b4cf8d5e88b7e5a95fe7e8ceedb93f7365a84d535cbef897ab24f0c89e7e6f7e40fa2dcdd1817614e381ae4aaa6a2a77b56a29726177be11fde594a7be76f931ba710014e48f3c781e35593a8de4cdbc07627beb5b47b173b36b96bb39916985;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5e9d75f6d90680b0c4d00f2772aa2c841ce7764249119fbcd9e19f357e8fd78d97bb2d5a89aac09baf824743f1ec2e803a7e2b6c79190a89900ec382904bde870d7a2a3af5e354b36a370ae4b01255452e75dccbb1eb0a9a17b839be115ab5c169e7f88d3aaaef9fd45d8781db241a05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h371a7694ba06c7902b764b80a9b1eaf1cf264a1a407e5112ef22cc36cbc91bd38f2d74bbee3f4dae8dcd0c3c8994c537ab0a48c7e7c201ea2255d277c3c5131b02aed604f10cfd0243b19eb5161b672fd87afddcad3be23ffb826411bc92e4d24d371e0af364f0ae72f777e85a4fa6b3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45acfd7afb5aba2aa2e2d52efefc9d3ef7d8d44e5ae851202cf93a775875e81e43c961b9e301478ff09fb50414ce4bffa745ff7dc0804df5abdffd927ed7cbfef9d66dea3ff2718dce2ac73428f3928badc450ac45816d43717a2558901c68e6a41032c132d95b1021cb9f1aec504cbca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h561381a55f221a7d4bb76ccbe39ea59546a5300b8ab290ae2366648f8855ddb8a27303893ca2f414ecde6ed12d15ff0d74739b75b6ba875758e75d0fa5d5ecfb35652a6ee7a9f696b9d28623f6112b353ed3b850c83ec1cfbed64575fc8cac66e11acf8ffe0fe35b35768ac81d691b11f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h267c6a5cc635e8ca1dd453dd3b7d7e1f4439e8b09b8a4752d5f31582705e67bebf01e75014a7cd7b3542f936da9a061db3bc1add6b26a268bfd3f1565d1840205db92c0200a3c29eceff5395529f3e4189dba7a5c94c6c0a7211f22d4044424a71ad6ff943616b7f577ea0f7ccd3b9fbf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h402d394f067629059e29fbb2ff6a8d28a8984a0ff234c7d120246843ba241a75ecfa8a2eb7eca070c9eba9ba2a4e682b28cbe4fec8f9f88e6de69b44457b7f2a6932a9a4baa499ca07e266d1663681170c615e26dd0c332d5dc263c1d0ae1148703df44735b4e51d0f3d39d8f2b8ede4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38ffb6b4cd5eb35fc861d27e088ccb7f130431e833faa0b1efc1598336a14bee2a1f4918bebd33036da858c66bd1b8d9a71968de3c0ad7c7ec6e89ccf91438d1f2c42177fbad6af861ba9f7ec0463747838d6e3b1803a5193dd7ab1add5fa617af66d70a7a5740767c89d87d6c5d7285d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he75a5f6d766114c27f9ff3bc25b15f34e6841d393740a10b014aa24a42c48b0ca22197950d04952e1a1925c7a2ad13a5c4595ec4ef7dd8d9bc60f8535565ccce4ac4de5aaddec9f75fe3873a1ec4ba48340fdbae1ec8be494e038d96046a24dfa78ba70bff4f3876528ef8b591bc1b65d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c0998830d9dfdd995d4ea81894462041ad15b7b4437560b28125962a903e8ea8101f51f6ae00ef40b9465db5d252b774f47532980107285a2a62625284b48de318ee67b09198f5267810fb1501b8ec2ea77384fec85012d085e59d05f429193990b5a16f95307a294b1ef4af5d86f81e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f7979c2e6aa47406076a2db25c883a6e0a212ea1563b2ece266383faa52f0db8c4a730297b3729e92ccfe94b59a0c36fa3a3535bf182a0761fc71cfbc7b9b74992c3878f3c26fbc4f15bbe1c50a692357c6c97ade4abeeafcc1e54b3eac1c2e2b875cda555ca0e26568f46a7d81bd57d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68925d7a8cdaf08dbce79142fe7de09a80135cb0a4287c3ad5e18889fb3abe38e96348bd156e04111a081bd50b94a2282b0c8931b50408cf85529b2e367f026dc7b3b807eee6a299364ffe69eaa23042e06b4bd107a16ddca2f943fa76f811a13d60a604d1a4c60815c49078ac714e786;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50108beeff55f2f70d320ad75e0a82418ca41c35bd7ad94fab7c4d609bd609ba9764cbb9275312e7249c19d5c1b16c51d2b2e4f5617b699800598b8bbc9ade93b9ce65969800ad943b4afd323b791baedae8e8259eb4ecdd3a76013b8b53aaf646eb9659e32e07a98a600cb1c65ab43f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc916bb61b84e565cab4124e753993856a8ab04817ee4b6e704a23c96931dd4040c1ca0177e49c51420a1aebe5f18aa569d86b62344eb44898e1e782755e5363eebdb4d3af9219d1bc166aed481c0a6143f52251d3fb5e8346842a1241228daacca287ef4d61418b0776f6d0574c3cca1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96cf50ad984c7acd72b97b2435cd4f8541ab495ee22d6700a3b0ca744940620ce6b60ef487d99bcd94933363879e3346332521689cffcabb13981242629c41a186f9a822d2bcaba213f5456a72b5de74a33b9c2abf7116d81e34b001122f851b16a71c8ca4509de8a460594d0a9a6fd7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he61f8fcaf008ee80dd00db8a7991f5dab0ae7c276591e10b50083e9dbeb5d0da14c780a202f5eb4880e7ea96f84d2bbd08cc993d5b619fd835dd999b7d3c4d146dc058c31275a9604d11ca8a88b8c4909724f22ebc87e62a7b239425e6858e32a8edadea4438428839826a3e7c269e17d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h800ea923f8f1e3d546514f3e47ecc493130322cba82ae62f8f0a5adbd1f8567c70be2f6bc695c8c516ea5be88a5906d905a14c207be215ac6f16ea0d353c18b5899af3ad4d98621cb3ba7a993cda78eea9009539cad05d75ef53bf38b14a983c7fe9db37a8c0638f6f1374ede54d45d29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49a3f2da5a9ce24acdaf103f4bb348c5e4424b5e70d32d093c441b6625f3ad40521edfea8d495bebb829f64eb30fc327d8fe9127953c2738de239d0e689656b66f0893dfc1d693dae32ba0d974ce5801234cc309a50a2b5bfcdfb0a565f1ce7f81419870cd97c042353862f32d886241e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6876d440298f2064c5dfcd097eedba14b22a7167580ac55dc5c6dfba2a6cb354fd2b270c037e4f77127df073135f661a761b8a3cde8005d70784bbf5e84c2836dc48c8ce2ef6b77f094ab61817fc5f3a6361ced4599de6b40ec3d90e04147a92007c4e7d0c3da6b2ee740e269d1a9b3ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he102bd1b4f3e5745d8e624071ab46ecdb3225501071dcabe7029537aef853bd5ae6b3ee3360e1fe3832097f0523239523c29f1679b928ee0a8437eb48786e920cb4f5382855b2c1dfaa7883d81843e2b2d0a5bc2030169c72632771782a3e4ab5aab1325d4b7506f339ac4857440e933d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8bb7b53662077c6b2a6230e35b6de5a61033f515b87c0579e736b6b03f48a2adb8656e26c1c8519ae1a5c6969ee3f2a1038fd44585dfb3b6eaf97b9504c7e6fc0529986f2f3ab8b315a4cd01b4dff816f9d0d1541b32637eec20d70d5eff62b59c69b7ed09e6a3034e7465ce6d629d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd049467c0ec368698552b17938436a55064ba825f9c6ed591ef12d19ffa5cec347f1e0e01a143801c53fdc238b7fd0b93a1fbf499b11fb6e13164142af298f5196e1bbdc3181c80a4ee0296471d123334dcd492d5ffec61a20bef4d3a86f4b7d8a81bddccb2e86fc77cf584e0c039e38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9298f152fce8e187c938c82d9c8cce3b6de11ff16d9b38b19e04bb638b304fa699ee371592b1d2d9e492d10f4d0fa7507c1deb78f7c421a92454020436630f9cd64d0077847a60916338fc5f0e50a5a9e5391ae4fff1b4850528c4bab5189f55de525cea5f16b7f59a6f525cf22c51e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc836344caf70115cd1b1bf2283d32def934793cd04e3c4e4761a6169f3b8dd5318b10c1bf64e5a1f9581e8219e8292ca39d96e2521f2f7c1c30e43d51790aede0679d6fd211a82c800bf050538f3d57de8c6eb7e5fc2ef7af54c14f3a29ab63ac08513424fae18ec494386b73e7977404;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb82a1ab216039cb0f0a9dcfaf5bb2822baadc2112f403f88116b4cce41aaa813718d48c57b01437d5a2808ceb19a40584eb0b71cfad2d256375397e258020d964257dcbb9c8d00fe01dec77989cb4252f9c0135b5adc93a925cb6c8c825fa0091590cedb7829e839be55f8a5fe575cd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfbf7105384bd617cde2b89ab165f18da6d225cf25cdeafc1cbd00bef9696fcfceed3940a78b177fcb6927b11c288dbb697babc2bda8b2ecefba01d823852789fea024511e4e50482290cecce2f554394051b821d36d87ab32d8b93185b98acae7da367117133de9a0d6525d71da6481d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26f457c0bf61bbd8e65a09e794a21c6899c7389dd7a2178f23e17075a5626a3c1a8cb4f8be249a415ae4121a516820ea67d9111af7cc8205700f7856f5c2527f9ee74572046759a708136864dd67474503e760cb62eeb4d010cacaa050c1af21fdea0881f11a30440ab639b69a403f4d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb07e3080520108e140ee83daf8bbb3487239b5ed077d090049e8aa40b16878f64277adc522ac4c8de6cce6f07aa7755eadf848e8d613659a02f3a60180146d0b3cdc356e8bf4e7edf7d9634db31f8703976d320f22da61f0714ef76ce70cf02a8f09ec8722458724f0da4979920af97e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29b5c3e27a152b3b85579230ee3239581a276182b1aa479598bfdb0c9bf4414cebe2a19adadf81df233963eda9310e922f0cd39c398f05394854359b70057ad3016b9c14e36ad4649d5fe1d6b5466abc191e6d55f1c57b64fe2f90c1197ada3fa530c8bc506f690a7efb91fcb5b7167d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he84e96227f3ebbfe61dc27cef1429014e6f53f49d1ab5de5abbd006808230f449403ba5e81eeb1ed5222a1d26a2e9ffe3d481cba73f023772f7f818cc52563eda4049657102ff2a1b4e59b582a5422b9ed5756a579bb7e381acc0dd7ab5dece13ee688632dd7ea00621a1ac342b6a2a7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6560ff42dfb1723489c9da29315433f27f8cf909d28e4ff56b7ba4f8856a19839632358331000ba57e63ae434500ae32ea5459e80ce60a5e05fa64b75b88c28326bdee19ac272abe667c5262c3086f64384ba377a8fe029bf12694890b67e005ab15fb9d0afc7ac574dd8eb02a5ca1d65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32313a4df676c6d8f6202d1c431ab2587d94fe308bae09d3ce260eb6049cfcf900ef6a1dbe4aaf0073f92e9fc10eccf2691863641cca68314135aad67ad7e4f4fdf0057fc81d5b9667c716f4a1a4682b4820196fd2d9a6ebcaf4551c4e0efe51001ee5ad0721b0a5eded74fdf07ec32b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5a015dd915b6f10c53c04073a3b8fe874dd8c4a7fa9cea9c0855b7c57f67eeb1b07546d114d543bb2009dd9502f4d6c996d05e04a5e0ab6ee54bdaafa1dd2cd417c6b6fe5dac3253f54793f1591b4a69aba063ab3b8f5f7e1fba7f3b7f8857606d82756834667641651c2d3ea6a6c275;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a5a51302aee1ae9b72037481fe286b73fff396bff8b2b80f1d6d9b117503e8d25a2c944949133fc67749d382025931d49ca95ee3221eac2064f214931be3a9fa5b12846db05e8804ed2a2f33f7349cf85fab79dd4dae7dca8866aedb489f536136ec8eb17ac6392f8ddfb0c2cdeb749;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cfa2ddb82aefb8b384954f6bc32e01f24f902a728af24868dbb9d30f14085b00323cb14e01acc9798bd7db50e93ed70a1b20c202cc980da6417eb89966745e5ce2c714fba3dd4c510458f7dc6da1fa94229b515e16ea5d48b507d6b665a459ba875fa14dbc5da4ce648e9d83b1b864ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfb67c52c5cb4a86d31407b3afa08f9abb72a127cc116d75fad8e28c85c9e93315999920eae713ba4da5bc74336aace2559dcd1ea2d1882d99feb3dab20442cba7a8fb7a0e2706f4d014155a85e15e979ab5e8aecc85824db4c80314fb0d0d81c3ba499ff6aaaf002ba7e60c53bb1664f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf99229a6e34952610fd3251991c3caea733c2532b348d13adca4b6b1a8a612d4001667f012bc17aee524cae84cb47e4249089597463241251c337945615f3b32b716f7f69660b748c99e481f51e0e0d19afe171bfffeab60eea2c86dafb344859d3ec51fd4142169cdcb3e5a51e0ba545;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h875b4d7249c83c2c994454486b2f350c5c0ca59d56ab0e166b67ff9ae0ff31e9c6df24386338bd05220db9d4bbd2a2e9a1f3796e882ed3ac2a9c5cdbed22238c230426b322bcf8738e4c7ca3374f4a9885c5c2b236392492a0c1d9dc7759dc794481d7ff7f4f08febe1dcb1ad770c21bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8faa4eadfe91ba1df547360587380e8f58f30b7cb36d147716ed731732cdeea7b9d1d681b085c597de2926006813d99ca246ea1cb864cbfb46944f9572f85fd2f301073da505f103c671d3c652a504709317c3fd1190a3afc153f884863c8770e0e82725174b6848e893a104e1e1483c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had24079feb6c1e08a95dd183eff6269247375b543667d5cca4f49358518da97a33b16a54a86dcd4bb43a4573d489fb827fae431f6d75c83799ae9c1bbdf95015d4a0f110873a729f5a0b7bebbd058e9670c00881644fcfcda0fc31f05d40f4b2eaa7a1be153f6c9d5dc4db09450b574ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b19768ea5cb96d1339f005b786f85469ac7730c7808511a38d0ccbb9832b13e5fea360bb539b50251d4635f8873c75c8c8fa3ee18e6122b2abd96da5a485709f508a75193283edc1eb62b2bf8ff8a27450296f138e142e12d99361ccacf761d083097e9e795bbd4a3e5a12c0cf320486;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6096cddf9497635262502c148230d8f2946b220bd6f26bad2a429ffd419fbf4cd53c9258829c83089bdb5f132ea5184802542b085a492ec3184bc43655982cf034d95087ad8fbdd886104778ae6eef5eaa23927b3ff467040cd0ee9499caa68957d8bc13c8f8f1d8af0265f510124c468;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f125344f5ba7d0927c28154ddeceed6200e8795e1dd289cbb69809693bd34f3c675267560fb75af0e2b159451ae7c25ef914352ffca49bc7d994ec8bf279460f109234ca12f2deaeeed9df96bdc3976c9487f19a61f85bbbc8d69751ffda624608243f01f668828298de45270cad1684;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1ffae908cdc63684dafbad4d47bdbd76222b3beb529b661fbb2db0406489247ce32e50c2a61afe2a001db5386be50523d9efea95b947a66ad6f195cf3245472f5a251288c3fecae96cb2f04f071d108666cc70dbdb39d1444b6260a41ced5b0b147541f6ebe6df3b2be8b824aa16b1ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h381c6c2b2674dd33351c588cd46fab533468496e2c97968d037c551bd0568ddcdfbd9c9924d5508cf90b967eb65e3c937abd0d55698a214554a759adf0e19f7171eeff04092ed872515ea642299e1795346c8c1c30135ef8ad6574279dbbf9a3e935635ba7a7dd64564c8bff1d2dfac83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39feb245ef21531e2c04e943eddf1715d348d14c6941a49a3bfe73916ba4c394edda96493ea242d18d0bb8c6ffb87398883a6f893a33096b2aba7ded47f651c1c1d1dda6b033b3eb9bd53884d4f99675e9129698dfc128aca600e9befb9528e75f66b98803d8cb340cefd0bf4020b0d74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25fa9ac671278f629884622f877fd84b5a54c7810f738fc31283d5183953c1599bf9b0d15628f74614b5a263be15e8f53047e2a0aab023f8eca70c05c1e7c2de6cb717b3eaf323f12634abcab89cf53bac4a4b884aee7b5abdf079e406b757fd6292df60b2514322605f06b5603ff6fcd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4bb331608f9dfc95723f4e87eae94f1858c310511ad990e244d70cccd2021513cdfa976044466ed5535e2a1d9b1ca4d577bab2e356edc44fa90148a1abb2443a9d80dd0845fcbe8e4ab732f9605505a2719ec951fd4251c64806326795a10787a2e3a683de88f99e63535fc0a7325aaf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacdbd212d3db957f51fe524026d7ae72a4a55ea86256acbdc35571e795e371d73b1049e514f4c28a6ac7d1ef6885a3f9d21828fdc3b80b2a1d7c66660f71eea85d0dc2bca6ed121e18995372c80116dcd7442bdf86ae637f9b14b63f731bcd8477e2ce3e5452339ead99fbd6ca4b2cda7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42d317854ca3d8800c134fbadc9a65dd21d8fda42c48e55de394c1021da594c55ca538983434679fd30d8f790961f7ea2ae11b5a1b99777f1fc142d5533489e3d90de3c8ae8b1db94a01b9415b3d4c34d99c3a58670eee85ec0d630865d2ffd2399a161c5affc2f56f5bdcec79562b217;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6392bd3afb437021f8665a3fcaad208947571988bdaadb22e051ee6fe4d5bd4f39413dbe926b0af1fcebf70ec3fbabe7570c36e41b084e0c117441f8338ee28a501e747b2ffae72e318508bc360a0d61ad70931c8bdc3373f1d2616bb4bea1d8af7c4039a7de7eb62e1c25d98415cc315;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84762cb1438827914807493b7afbd3105d25eddff59e774fa1eef1391bc1c8a055aa8511bd598f3b4a6b7639f6d2f5b4bca50a2838ba4c30d34bfdc704331f639f531e5353cd2956c784365623b2a558bfd84f41c6cb759698184146f4175a550dd4d47278711728606e845a2ac298b21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb06a01771ca4575c80ad452046141ff5eefbb190bba788059e2e4ecb7735077e8bb276142e69f367433508ffd8d13d0d995b5a6ff8f7a394ed0801cd5f96144690fb2ac0597f5072c0fea89240e7ea04a9b8c393a5a408d61af13218acafb85e538482b8ba686b1583a9eee4711d2b79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc52021df97f110480b0afec00bba9eee770144942222d96fb763a1620b8703bc710ecff87cee2e57777c7a4652a547fb630fe90458c0c447fd1e37651748de153fddb2e60ba780467c22b836b1861d4cfcb1f67ffae882403ad8c67cd5c115a19b0d0e88c1c84591e2aab892365b570f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he829149a33b1e3d2ed4d77280383469cbed88a47709ea043b2c66207b964f74d70030a358005a749c8c580a3589f76a4e43ac24b20fecb775fd4ab0a07aaf424c52b07ce701ffc97d2f2cd644d35811ccf92452f33559f2ca2a6d71e5965fe850bede4c7ade0aeeba31c7dc3f3b163138;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he173f4a4aced580927114d093bbe2787b018711e3da85759ee7fe32297921358bb9dd3488012e1ec8511f422162ccff2d8dbb0471a1ffc4e9d273fad3c4987c08f648061fb66d9285564978d505ba828c84f663530fba3d00105b6611841796b6d6bb901a9f95b8bad25a5b6b26e1f74e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9850dfd8b2bfe6fa87afdb9f667c9890c9a6b3970c5be6e4d743e3c603e3ceb73710f9de667a8b2aa7d2157b32fcb93f4125200912773afb84932fe64ff536173df89b30ff2cbb6d9bc7ff0820de32defbe334652d0949a7b12ee1f40b3aeeffab327a9da1c28599a4db1db99ef711ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24ff2fb6c67b58f25e1925e5546175af6cfac8ab6aeda9f5a99f1e1640b85b266fac3ec3ac6f3667eb0b5a1a20e8fbb7f91c697554217ae867c725448fba4d39ccabfafcc0b68d9696e0afb4fcd78e76c7849466dfdcb15e50d27eedbfe43bef1680f493ad106f6d54c86b29f70901c47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fe39fde0ca65ebc9e4b78d312c8b55734877a234462b26d3d28b428c3871b71a3d64578688149b8663b217883a0a07c9edaab1b88258eeeb834d0ce6c84c973dd4c9fd76142c2d3fe1756501934827900b8967cba94dabc249c82e2bca69b66bc9f8bd24f562203809c60e91aee51d91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5890e134aae829351cdc73e91522d2681ed87beb1e05a1e8766665c09f1722549b75a6306bd102a8cc17891607896d7363b0c461b0afa9f690df0fb3f35e06257e51dcae24dac766ab846a8857ae727730e98453b4cc2e10d678622b377937643d2d72f22bc37cd07d00762c4342c588e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cb428dbddd356dc6195510e19183119fd2f5779a3ae47554e5e253e1012da7a5aecc043734d8b7f97c6bb63397ba9a1477b3f1a41138bab65f91fa2e755facad8d56c1fa138e5731555297cdaabe68802e8c0f870129be77c2dedb92861066b7dab3639fd37429d50682052d57de499c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36cd591d4e7f9c74993c9eacde382f0147a5a875a566e1bb5a6612f97ae547d77b22ccefd9ee24a554286adfd2b6c6b541071251082123e4ba77ab609b75d0a00963beee3e575a89954d0e7b1436a66ec40eac908afebc70b676dcebed14e89482ea2264137657d17ba7502c8ece3e43d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70376b733c97d46ed23227fd9181b80521b8de2e24faa528da34d59cc9e1cc1394fe80353e864bfc1a9b37eb68120632c34eead4b8e04859d8806d7360b3f5c83082d3022ed7e9f75ecbab86dd59e236018b64fe7e1dde5f12754daa4e9a32477362bf2699320f5c881cc027a769608aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37355bcbae31f203b06bbe04da938ef9e053b6739e2ce858d84ec47e2de1da29997f08a804d2b04e92fffabc2e5ceecda53db5ab56d0b853f4488842b4ec384935ba8ea88efb272f580feb6461e4e59c46f1a4b1e32a81db1dd309271d510266ec7680820ac85ea5b9a0a7d9107d7a021;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56a3cd70372f6ec343918d9e79bcba7c9833bb59757f65353db98ea6bedf23caacef7ccef8f35b6424c4fbc4771f464859a5f5ab87c40aed0b54da275247f1938539789c8afe5b7d183b96a903cfb2753990b6f0789ec465b859e64d44dd7c32036fb3b8b148d4dbd05d1b33f47961f80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3065e445ce04f0ba91ae5d0ed64a33984d0ee38ce1d35dde3149bc13ac4d2b0124143c44d335b3214fee326e6a55ef3b129badc1e7354d0858c830213783a80aedf7f92ab1d5576cfa24d79d6f798fb1280fd68ed9236546995eddf64382fb0d2e31d4c90b7c36d2aebadbc575545b3a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec34c62b4a7774c2079e0850683f6563fe180063570010a39c75fddc786fc296a9fb6b5b3cde6061b57547480c3f709130691bb89d9672eb0296a39f7b8bbc56e179559c01375f8b64f87e1a4c608eb162a3e2efccd48584560acd3b21cfdd2f14ef0f72dd1536131e8073686eb9596c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd1e44806fb3836253eda2ca57a718d8a911be4403c621178b4b4b80bcc42c06af0dea28d00193416a89b19f2e82ce9c2f0bab7200305cb903dbc1baffa8050b7ce56ee321c0fa4e98d40b4a6548955f490a5c2b5acc288061c50a43d34eeaeeb1640f235854c43788c9682520b68f0b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48dfe8ce29ea1e428984624c820d781d916b8571dec378ca829eaaadfd40a7269a9d07055443c329484aaf080dc59edacdad87b293a6721c481bd788f70f081cf1b853f91a36eee7f76761e618589a1ab3824515f9c0824709ad5afc94498170185349fe463793a8b742f99c1f9fbddfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e5df3967ba6ea6666ab05c0bf4e2cb4a074caa139b00111945ae49b250359d467dc0f046c3c2639321c61016eeeb986a2eb03fb6519de3b894be08c41acf046a8facce622c995cb09d1e0f024285fc26a269fafcd708ee27585c36bcff25b39621dc87b7b84daf00474175b915365092;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h407765c78b589f6ec700105a2d0350591e9419b50c3f8a08d8bad61f2c8cdf2e015d5dad7eb94e501355fb601f16d07fe37f79e1c8885b73d3a8411a0bcd1bdde5088550009061e362243d7466751e22a90f2abcabfda42dfdd25b41c084553df5c2f813816264867364345fa7150e4a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7facd568184de7439c1286d88dc7150a78673e9ce4ceb9c0275a3fb04ec0b60a5b4c6128d2454f8ec99162cb4df789d84bb7dc2c46edf0e6033680e91074e809a3ad6bf62c8750ef8ad87be2ae0540f8f31c7bfe0955d058850727f234453ef684953ce33c523461f2d3ea688b2043585;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb328e16a52adefcd79ee8e0cead4cec4c3a496d7084411992b99d4426f8c8fa03680e542409e0984da87d67491756b302775c04fd58df7d93d51bba066390467dac2fdf7fd55fb471587372757a8577bdd2fc31034b6dee0c5d6bc5d19186da7d7f05501c6e0b4ec3c4e89059c01e5e8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24c4c5aec2feda9739e63e5324e703cb8593cc879330601986bca85f0595391e9eaed7da507dbcec28c62ede1ddebb0540db60895eacb4d685b8af3d17833d609c95391368ed5e55c3e4b92561503df6050933d1c9e21c038b0d51c465ab0130f221def71fca2d1fa7d4467f98b470246;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb3135b50017d0632e3454462b650a10ea2da2ebf226b4e031024586e4834bfd765734cc510f74f58eee02913f3412af7613141b13e54884f732a2f6112e66600675c6a5cdb46da5e81e543afc405500d26982909015099a26862b0f8c8e07773fa8c7d6f34443e9cbd13b10b7cbfa4a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19668f7c6fec4be4601544911c864ec7a636ae967f056c38f1bdfda6fd48a298f486cf191b7422cdf9d5062f5ba065ed84ec3abbf9acd778bd70fd6127c25b1f0b7286ca1a492a1319437e3d19d9a6635cc2f330aabadd96c0721735c28e53611bf120f2e4f26b26727b6703748cf96c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b638d73fdbaee8a19e68d9bb5eeca8be5705fec42ba265908e4ecbd7cb6c8f859fd44c5293265ba46f4a5e8529cea73514a0c8acefa65b087abb50c91a8c5402195d8c8c50722fcc8e82751d504350a3b451ace1785dad50c065a3619d94f20d372435261db875c641328ab88595e098;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34ea732a4d6d4c7a668e51cdfcbe3cd00230ff421c0892a3b7d2e6b37f21eb4409dc062db7dcee346c647939467a6a1c07ca91dd454e536bb8a0eb947ccf9f61f0eb4da84d9e7f5549f130b042277cb681f0e575d51dac21e14b92b187c0aeadca34c25cd56b82c4b6f4c3a30a14bdfe1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd86ad3bd4460507534c2338997c4e6b926a328c6ff538659d035f6ad99034b8c7f8a195507abc9c3a1be3036b4e623ad500680015e70021dc39b79e6f466a6b75b50945a226b78505a2cd2e7e2f6d14b3add8e2ba186c3aae04849d939b0c18804850828abec3421a6951b27d1bf2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fea26945f34776c6488e74fc1c29a9b21f1a662cca3e4ecdac0f3285f4c53dfda6f51e093f87af5d062f4b195983c6efacb961ac6710097eb6063ed3f4c5950f16ac6456f03822f84e32738b064f6630230ad8f19f350076e3ef9fac11a6a92038b6f985f3a6a4e4fb84f8da4ea4c4a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde60764c98b3076a9fdc557b543a6e5b831dd24005211752b6a1ceb93f8f6f189fefbf99298e4ff33cd2fce8933c061592b377a385b54120ae0915fd616434f34c0bcfa777272750a172b4ebac74bb93814a5a230496fb7dab13c88d120c1e48320b6ea1e6961961bccfdffe09d993f41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c2f003c5bf95dbc270f594be63e7e4754bc1795877f5bf0a35309956e4efc4d3fed22a31b35c9e8f08fb9b7c0ee4cd20ef15ffddef4fffb8be01e7532262cc4d215d8410b9031bd87046814ff15888db5928bf40766c394de17c4b8cad050c2b52f9cb95787734e58910cfc51b00601b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0b6ebb30d7b081f2892689e1c20685b85f85f0dfc1e9c079056f3f2ef187497481b8d68680b01c0e426c1dd54dd1b1de83c265f40cbfef4399064cf6d588dcc00ea8b0b3068eda5fd39cf8270d08e40c172f9c2f88a0f5065091a176352b2a9de465c3baa6eb068be9234f8158e86fff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8d2d072ff7253bc2be92cad711c26e84cc03acf71d4129a7edd39638170c6378ddd3282d6e3d3c04e6d37837b713dcb8702b0520f7218ccee8024b45b11fde4c01a26ea961470cb20ac3385ebec9cc49e4161aa7bbc4a53a5b5139780579c6cedceea16d09b81e2c60e77e2f09a8a2b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7b4f0ae855cdfac9e5c68888fced779de20fcf1ac7a35cf9f56864ea64463b440c90528c6eed79dd1ac53c2c1783b71d65e917d3ca2ab464f82c928aae340f851b88dd3270e9873c6d9719f509ddacf4a18e0b4fca707da4883205c2f7ef7858ea1b077f6cc44f03f996000639d8eefd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71f87465b9f905233cf4c858f5037756a779a2e05cd24f1729f0adb2f047102d7668fec6fed7feed531872c9cfa0cc4ebce8936cd6f67508fd413b4fe33768d85384a836e5bae9fef2581e059a58287f9d07a8bde05f88339c03887d54fdde8f507f355f316bcf2bb71328c6892915797;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8617ab2eacbe4a46bd29f566543fa38fb69801b2bec6394a6f9444e3e6477a13995313aa55458ee0d287bfdb28e2838beca4cd758b7e8360a588ae1981ce730dde3aa034b00e5ab35c81a15f1893bcce781a1c55178410b6efad1ef6a4d047d2cb221acdd155773958ede7ebf64a2973a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha61200baa63015c0b2be20afb1626f0d27c01c48ec511dd7110eaaa159b2755a1b45fd969f83c9315614e57d4e532cb9e52fa5567fd04c8a7dc3dcbcbd38651ed511db8f24b28b1139ac9c1017f4fa867934d7f94eba8731538149a0c09cc87c1b216496d1a84d541c1a5cff640ef5621;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7534146bb1b102e71c59fa8cb3f26d34fe873a9b3026e0e140a90b2f20a0c9d5b7872b16b8a4c7c0aba91417d7f2beeeeb17f23308c4f466b4ab06ef64054ddc8b541add4f103382010455ee60dbab6bd4fcbb3dae69297b1220d06190db13e150f92ca6ad236859aa5de8c770c3ba4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29cad58f3389184df065a5a6c3caecd33cce72919f09abf2e9115d05223372dc6fdaeb5e8a0b6d3ff9f4300feae1978411f564c5e5caead110394b9f544c387df9cf53a5184b096ff5ad2c90378318f8102bb8f68ea9c93e7bc085c98ff53e6956fde0539ada5b3db9092cae40c8eb6d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbb4d6ed001b653c1b52cadbf00602b2d909d1857ee12a629db68b35dd1a91382ef7b76e58ccb33893090b20d13f0d6e6c822a2a9feabec79d75e4f9d174861b88634156442a4015bd7e419bee813ba72d1ffa8645b2687f6794b62185e92cf4854478ea09118f160c87a0575ea320bbf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee42fcee2d78ddb3a24c63e21d0d11ebb94f83b179103ca4338fe92dfc02c913848947b7829995bac994033dadac9d09cab2a31c79e53b47dcdb53a235706bd27a7c7693320615fa2d396fd058ba70abebd6de16a6296c425bdb50df9e5daf93f8c98fad9ab0622943c99b692130912b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9171be6d5634863db414f90c429a5d189f12682d7c578524dc85432126ae8f6a52b67107b3de15e44fb8e346f38d7cabb1a18d0a8afd3e5c21c8cefdcf61eb4287ea444bd383e3569220b0394888f367e0ca09b5879bd36232fc917af138d9a4c099fcda4852a6eb2f28af9238db50a53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf37acc5747c815701b72151385e5fc703adc86506f093272e9cbf55600729e530fd307b3919b946e23472de9f5dd6c7b0fdddecdca1604ecda67ef578ec8c224e62d445d596dafa074d651652471c0c3bb06108ca43a0779cc174238287291415a6f9b6fa73f98d46e929e9b1fc864b88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfbb7d993d72542770907a37076700e8db76d673ab61df4d4ad2af0045dc2f021df0f5c444fdbc4d874ef5d524417880bb56530ab426ad557445075bcb9654da9fc46e934fbe94996639a7b59c15f5cfe76bb8abd129b8340a31dcdb143c4c269246965668534ae35ec1500e2088f7049;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h587c56d4d07019092bc824bbe8fc06f37a489c50403b717b7e24c6a6b0e76f5c144895e3d015544882cce02113443a430c22d4d72243e3ff56414ae5609f9acca402766225b31e023aabb3fbcc4c75589cdb1619954bde5a5453dcb9d46462871e760eac18ef4ddce7177acb1c59f8cdf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4c8707383568f2e274bc609771b51abf45a9fa7c1c26e7877aad4f40107d4e516875eac0f1ac759bc035c90a9ce45909322507dd7c5f0926522a6a4ff79212c0945824f5e183da793044ac6acdb0fa3d4c0aa553ebd60fe69d6f46f518585394636ebde923452724df0342dbef084484;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7085055ff030f9672b53b4e2f4e781a5a819d24747c796e80952f8596aa15231e57a535f9df6b612c467d1ec63d534121acccf054a4bfa3b3b570f71178dece66555221bce808eb3b119adc787a9a4233402814d7af70b7e15c400ffcc61353f2cbc409d92bf0e2af547b4ddfda9382;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58dbad001568c049e7271b3d9246486051b2b0370a2b8f5ee1115ea2220e612430c89b92f364210919ed3def2c716f16010777b97d40695a77f7ea1816a1dd9b3e3ad44cff906d1222339da5dfd79d40e6fc143b7d0125a742a45a7b61b4e569448084744ddfd3134e8c954c5e592b1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc34800fb7a403ba64dc86596b1306b91289cea5a68711cc1fa39b23a63050b36a99384aa6b07867653f65f347234ce9217c08e023386b624b5554b56e9d531b38b31c65b0b40e6110cf5808769e356ef71c4d3ca770d27c1ad71db7fdd8310f86078e63c5dcf5f275710a32fca38a3026;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2891ddcfb3e9f0e28624daa4be12624c1f3ef87c41b6edbc111ee07814b65291d25528b63e65a8050fac313d748fc0a8367cd4f59932d4f34fe5a1c4dcfd716f6229942789ab725609a295b15a7c474722573c2c1fc7e8ab9b275fd06f1640ec4a18003d055a719ba19a96dd10a1ec10a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8af0ca5a8b77f43677104e2d7b3ee16256c0e8b52319a09f8647514b3eddfbc0dff660d7ad1949919e5ae2f0a3b3193953df32a2481c78997561a5b22f620b46baaa61616bd31fa866786828812cbe490b4e45152354dad32784ad640c15f3a51b9d11b185dcb32d322a640e7f5aca7a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he99b080044bbeec4b27fffd02a825fba51bdab01186e42ae37d35a102939a1984eb5a16663c4c5c6242e7e2c115cf2e9932438c153dab66f25c5336b80261cbfff2aec0115b375f23d203b05168e2972716ad41358beaafcf2d8d9a6af4d9201d39f1252a4d41b3d091ef71efa3bd06aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa97ebe2564e9e1b4f1a4ffc6bc7e2c413a805bfe4dd5cbcd53a0d9f1e2dd6604008e12a5ac53c796a362da687184a89846f629bfeeb8f43305754f2a40c3a0f61082f41715ab05b62949441e55d0e0c20a57e13e77f0afea59888461636c71181e11458274e559f4db404a930e5d27d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8133284c3bdabca42529f86bf0daf65d6bd9c8436076f9fdcd5e8b8e8dfb0bc22707382d6b8bc96c69e3831282e9e456aeef7019211c513b139a3087efc62781608df645d9976937ba984a72d5a1237c7d2e4edd61ab30122ce2f210ed056985c52bb9e323db8a47f34ec0d9dfbf9cd17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8301550e0d414e073c89f1103194e0b8e0d6acf5877e4825c3c99a176462973dc609bd18a017f37151b5e67d110c22df663b4bbabf11fe868cef6143703b706155944f83d1195b80ceb31c4e4bdee01c1450b0b6499feaf7211d08c50e384ccd6b8b8b9342928424aada4daa44f21fc61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ef939d30a5fe0da8f99d02aadb6b416e1867367d6b1ac4440985f4759fd5f37f2afe2f4e61cbdac1525f7bafaf139b89c1a75e73a74c7a0ca1675096831e3ac448effd68b0ccdda9e82e8c84ebca783abff2ad8aca622cc1d6f03d72f181fa2fef164d879b72a1b95d9aad73dc52bad3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2af2b1c344a643c0e2edf7db964f95e9cf83b6de0df85c18f2902397fe34a3cbebfabd7b85ddd99fdaec02c66fd41978f17f3c48ca9d1cbe5ce34ef9698ab280cd352c9c5e15edf7ee04d09fb44f896041bc34e36cefd7bd5780804fbc5ba6cec240d28d7fa97f7498d4fd7e975f229ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ebcef9022d7dc4bc7fd90bebc0d31ffc636e34c6ee73b88009fb76387d509231243ffe337ee4561b6ca3cc9679b97e413dd44c8f2db04aa44a41bf66f85b20750b3113b60a97b01846bf609056c8fc4b4c171219a4114e2da540a3bee292c050a4992201fac95fa150fcea0eafd5fbef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7bde8d9f0e6f042f98ae03d9db845d5fba3bfb0b39d30fe931f1796ef0ddd71920f76616f083f9e2049b42b2a10b8c59606b55d3169b948c8d2a2be940623b0a5931568c8c6bbad4a2977f697e31c7e0f197012a4f4b21e0558254cff712bbdff9050ca4d8a61243fba564d7636fd1d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bb43f05ba9426831c8783a16160b13c9552ef0d40dc6931399f0166684f3277add94dd33a4c55a5a5ae8d5df95df2c01ed9e4ea3aef1b34ca850c88b42132b25ef1d7d81693f7ed7fbbedf9e9d88bab4e0ec5a8bd5e8101a776a744453705ff55e442df20689e0031cfae019d6989881;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h590c1ff896cedb813a933b847198db3eb8bbd09eadf7408925d9e7a8b392f186ec326e399b3490aaf16cbd3101ae46854f7b397c6207125f5a560236354da97e7b2412f94145d6a18f4799661ea6d6e7d23627470c7707b83e8a7665114ce07ad941037e1fecd8f9384ce9994531d8f96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1efc3e77daf128560d730fc2c6a0dc8f4d0e2c274d07483dae8f4d714bdc5292832397a947c85c59427e2aa9edb917f53331d05eb2653d4594de174c37c47ccf94022929792cdf4ef11ccc2d3e1126989b5ec0d81919184e53606c160018cbe32c21308a56c1b9420681c4483b2ed478;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a5e168c0bd231d8c26f1b1afc6cbb08949619363c9f03195f5451123d5f83082f0c4067f45852e34b66663821508d7d7aead0f7d20090e4c4e3eb841958db81cf6e70a4c945f48ace7f974515532eb6937f8b51bd550d4ca3500f5f34736600c3f3061fc12e7083ff2d0dbd0c167ff77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a5eb1ae81cd0e8f80a7996bb48198b6bd02a1f2a4a60646bacf31a9507f3318a0aeaadfb58f0ee07ad8780720827fb53dfa7cfbc8f59b2148ec7cb4baf4acdef5d11b0c69d521a60adaf450749087ad01985749bf27867d1d6357f727cc93307badd44b86a93f40767a1f373ee1dfd80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccdde48736e7eb302dd3fc6e27ec5b9e87db18b6aee311dd7ee57e5a44dd9caf581d69ebfb49a625454ada7a4aa9018d25d7ba720a9198aef6d30d5be3c1dd92364f122a8a71b595f51e1bc1c00a695d7c11c33d0cac7ac23937b98e93527ee94624eedbaaa63f8575da2d79797923c63;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7d0c0d09b11cb807bc1dbf5350e8f394045d7e257e5431cbf4b6fedaa6efd3eee81eed547d423e04f9b942f9ef2f4f934b85d18477f90b100b4b48bfcb8899931abec205cf692eb85d05e230b31c2de0ab2d2cc20bafcc6b143764805741a8e61bfb05eaae5786df8859b8d8dddc2078;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6f8e35f3fed7bfb23cd591603b12a8437ece4e46f48ad8cc6f65caf6a54c520a0ae718b43842376e810d0a5d60891e97c87265df7b451c3089de84d3dad722ac3ad22287d7a7e21895a08eedbe7c5a57f32ee8ee6186b59910bd1c8284165457903bd3f27dddb973d87bfee1fdb10d97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf399497253ee4ecc8a5f8207ef5d4ef23073acef59c3d330d86d103d3f48075d3aea526303e579f690090a6cecb391c9546689d2eaacc703f71fe080c78b216e3771b00b8b9dd2ca0dcc50238845e540d051b78989af7ae269a2052d708c672153069bf1adf721f5b9e548c99e022ce1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b7a7ac6b0fe63c5230c172ffa682b1485492b568a47e13e9b5927caaab82b429768453b1b69313ec894be05f65960edbbc28534ec51fdfd08bdd7aaa2c7f019ddc7d73700481b8f2a20cd4ff6c7bc75f9017909d322c03941099db791e02fe48386f795b0a21826b718743b4cfa39c7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a75e47cbb3624a6b18476ce58643b3ff80b64ce680e14f33f5bd7ab9945fe1e7f5cacbf146dfff36a7ffeeb39371f1d33a479728f1888c296a93241656217325b595adf7a9b1f89364e85c440d830b5dbf7e1b4f025bc9380215e9b39ddbbcb8276cff82dd32908d8d2f1e9346f39890;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb54594c5ecaec97326c74aea42dd991b9c11d095d8bc4e6da628ecbfed30b056d45336437eed26ee4c93189b987285b9c082b482cda78773c8568d5695d6b6c6fb1c5acef2ab1defe77e246db34d198c795c2fb912ee7a28bb40e053ce1eeebbe9ea21a70edec70975abf7560c6bd17e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45fa767c4b3bc892e802197a13245898bed7349a274802a50be5b50170d70941b9339cb5a4039fbb69d4f7718c4902843cbd77347f34521913d4680fda401d765a99bc5a03380a9f0bd0403d49e9d1cab0f291e5590fb4825c399184730daf09d76e3476f3e94ef25a232476cce0bf688;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc21e4ec3045efb896293dfbe854a22fdedd38866ce74fb5f922892a1a476d45af6c96afd8b8b8e64b5f6e6a0485ca4b4ab353959bb3774214e242507176924b30ccb08ed81dc804d1f83ab577e79517112c2480894803bce7b9dc64e2b6727d0c733d90ced852b37e181790df2c84d055;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d3722674a12e6d82f73936696f7c053e27517ab8ad221fbc6ab06def3686adf1707a12e22fc0491f4b784f227cb1ddd5b2d73bf2d1aa966409b6afadd528ef195ee5f73f91d70fea23686b65057954d260b132b94da001f4aad1e82dd6b8449834ee6f621a0ccb9fbb8fb2cd3bfad276;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b507c1f851f98ac9e75a998c6360089ca677bfbdf48c61206c61734e320fc6a389aebcab2b168869b11c273a360ee0a23e5c9fc6494a987f683e71402b9618d29ec8ec7065858df8e1cbc500f41b460da884373211369620cc077884eded8eb6bd3bf9abf5262c425b774eb72482d63c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89214e131155b2673ff4d34543182fd60657ea59811e493908df3498c57f9b60a79989d0a47d38db8287c5ffe678963962b6b65b8a5feca71da5ad3ceb13e70e29f22d87d553c4db413662f66619b257f38ef0eca6747274d33cd4ff17cac268fafeaf1bd370ec7c17b5d865606069db5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a345224df6881a583ce311a928f84f6ed555f924d6490e339af44fcb252cb39834b95f275b316acf8e6f932a4664b503452e03247f4c90b76b0207e1e8ceac29c99eb91ff328d1480e3fc6eba15ab303361b2f6b9c5646cb8d1c0dda025a4adf6e61f6537e16b8b29bb9289c0a353e38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd178c60df510fbf5eac7e42f5bf0f04606acf2d070a1322140edd08821e24fd8b0e6fc8ad9ca9f8e33fe6c1d3644b4f653c06d854945fb91c6960921bbb84b3e6419e46a3d42535a76ec6641d67c851fc5c58d04e8ad48bed049b0704f0afc549ec13b4bdaf39c0d6c6455881f63d9b70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10524a5eae00d365b199cac156a342604ba66d1cf4d7f3d796edababbac7e89d149167f3ebc5b5ec66d1d6f326dd3d9a71de2a6d61578ec1c46dba778159a2e74bbb2a1d96c7114aefe78965d00fbec507f9b84033684b00648057fdd665d6579c2a4b75f06645a95c3f4a18949454c77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd85ffe35d02a9201381fed81818b27054d0d98ad2cedfb58ddffa2ffa42e6a0d43088e25a29d887a4c27b1109df6bcfd75869e8c607a515eb0c4ef79e8adbba3ded5c022aca40435ef0a9a2cc3ec6eb4609f948f621e0ce29d4733a3ab13d5c7085af1a5317744f498b45a9ddcd4d4090;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2dc55468cecc4b1f37829138ee75da8337bcdecc4fcedaa8a106d5ffa1d222bba8331f81184f3565b4e7d6a58eb7ea19506dbd022fe21498db5d1d278cd3892ee87db40553d169845ced8243beeb7e28960b6e3cdcd857c8ebbcd83d6544ce632b1a2b0d01cb97cc8f9a00f1de6c47b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef7a9f53732c7b47a15dc69a8103a92395e942e4cf876bfc270841ac6a5befc9ac7f358907b51cd2fafbd87c0c8f39c4b2f67bc0d9256361f20b912043899478006f9b885b0edf327e3340ea551723f7adc9fe710abaf4c7511bf6a2eebaa5d216ea433203abec86449f89f02545ad7ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f704f11a0a7a4569227a02f6d01d9c0b9dcba773c9e56379eef810bfc64946ce2f683d0e4118a8abd27a71b3b35ab7f69d18e5821d1a710231aa99f9d4ebce3ee95f3a8801a43ab6e1d414f7ba3295a294b67b5bc4945469c3a9edde654c9f03478c2a325c60fa69b9ac9d496014f812;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha27622747e31bb1ab79984743aadaf45005c9223b371ba14d15361b323d14a65cf176d557a6e43fe86215701906bd778109ccc219123ef10c014bf27165fed6d07ba7b4c357f96314949018bdefb14ebcfbe8c97c58ec9a5d17b3a221c482a292b5b18c7296e63c27f3c6a0991e5de0a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc824c6143b007dbc6becb865498b1e835b6f5aac1c3d57c610851668fda43087f5bf1c4f3c2aa93765e72a624b7ac585ceebb6df660ee8a43ae4892581a48886dde0803fcfbe44a65ef1ac05098450107860fa3a6643daf1dd47069b0266bdb3f3ff2d3999e7f6e9488a0f2083f2e2f1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96130c97a41f4794c85cab88a09c5dc76afd2baa4732f3ba14c1eea37484abc975717401c004e6b449eee4d5614ad6f4a41fe0579a702e63f94a86619d868ce3dcddb37be2c2a894d19e7b77ff2550917f5dc361c40e03c58576a77235ffaabfff1b84091aead18a60bca09325580df9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c88de46d9e97f42bef4ef15c0505fedfc4608254d9922f616eb86266d585d648b3f21be16ed8fdefc46b4080479d44249c6c10ee78e7b897deb059bc0fa01c54b0c5f174692f447fcdbd8e66486eada32a976f32658b287b15425f68b4994bd916b3726a0daa0f2f92366121a281ccc3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha72d61be8531d98c6ce5a2dec26da5e6f75c81875564cdd53c69c3fff66ad6d6dd625c6d367139642d4a53b037d88c6e3ec768b2537244114f0c2d2dce31d571eb8bbb6230d5e1a2f428fc0ae8cd2fd5268590149226e00c68fe0bb8a16678ddc6330fd7b0b0f5a83645ac5bd2f62cc32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5ed8f6da6c64bddc87a2bf048fa37d73ed7be0d13a74031ea4f65c8941f1776839a1a6f0f5f308bb89e50d0c1173984d9f9249bc967eaa7ec55fcd44f3bc718a327e741748d16d04b12db09aa2c899bf2d0f339f029b33bf73e9d56ed55b835470c48e9009c3827452cfa58c1d0b1a3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8d8cb0441cc758db63c6fbea8d88bf18710599d55dfe923305d608707e5a2b3ba18f0744d49ece3b318d9f8a98666a4ba5339ce41fa04dbc88b6951bc5f8bb0cf7920e65e979f75024e9428bc192098d46f8b1383e91f053b3df681ec0edc23bd3af22f6ad71b6f016a404941bbdc1a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2912cd3450b5b6bc112a1c2251cdae54c3193d1425825859646984a661b6c111b23674d05af54d12a14b1adac6cc11692a706a66cf60ab4f1222885c3399f7b04146d604265b22f0128db486632ebfeee08d80c5d6aab208cf4a9ff435a3eb91fde62ac785eadc3b62668b445d5305601;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h348836179b96e49d3a928e2305a3ac1198fd6b8d2040214018dbbcf83495f1bbc33aef6cc7f5e20ce8a058b325245d863c6f64136096a643f69e02836a43c475e19a3b2aa4d18096ebb216f51721b0f0769c0c53681793bd695e23de4036109eb77a00c66ce64421a8773e3db122fbd5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dfad986c4aba87c2cbe95b11544d832cb1f3e13bf93875756555c2a2bf22fefc035ecf8a1ba9d648da78600fe4a3f2f0db49e62f72e9dc9f25b0c16d53dd3a22c077bd4cc2c8c2a30f3fb8719cdffb82774ac6a2a97e7bf4be6b7f7825175f5e856c19076af031687692efdcb1bc1524;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbdb63779aebf0a81d47974c5709f068dfa46df94f59616def4bc5deccd8abf77f0f41aafbb0c1c88db163f9f417e83779a44097b0c7fcd224726fc11275abb530b85cdf3fee1cdc4959dd034e91def0fbd873ca5eaa96b513c7b891ba3351283a1a12056438f5ebffd756524eba68e42;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c88df353e9934b0f98d3d3f35463331d9928c5b5f9780629a7bfd68cc3e06ff6c52f4e2de7c641188c8d8848cab1996e64f585b3f3871360d14198d8b5f65d69fc12d63db7a00332d0a709f5c762ef18519bc94f20de3984d165ad377efb07a21d478d0148b19296f510066bdf5fa3a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7b8627f2be507210473df21a7d696d3285e4bb8a6f533a4f85352bab1926286ffb36f32226c09ec42880bdc2b9d402d41b1b766ccc4e98aec6e7bcb1d89ecfa47f9446895ff29e15edf88cfe34a2e236307267c0305f210c8409bd60867bfef8c79331ea23e41909932d0e47e457f601;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc632688e71e47c957d420dd150ddd127672f52b240e25cb46a2197a7c82a554d172bc65d161840ad48f96686c2c8990fab4cf50f0cdb647e1bf7e102f8fadd11fb832ab8a4f3f6e95f783c079bdde2d2a5cb5e07e4357de5982369422fefbae784ef0522a6b1db24a8c19f25c8444fb9b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h843535f03bfaba664dc4887de97529345951543a30e80fd219009f227b3b744b3f8a0059ea777666726b93d3f39fa59df18af14a1494b2b78e566b32319f32a3df31d227ecea8f9f5f061e9af92f40084be0d56332fa3212b114fa02d16a20e57336a4cb0274b3620f0fde0b413d21cbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a14e7fde528fe5978d78ab84d28b492f402eee655172bcb2d775199a45b585ca02a91dbf1635b337fa86643d4d016b39ccfea58e0cd97c7f435ed2ece66a624aada47d590fa1c85b819146f03e83523dd9799c89165dfef72be980ae985fee41420895a10432cc68aba44be95076611f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c44659ff2db147c1ecf1dd41e0de8f3409aa57f0271a9d17ce63b4394218ccf90363931a37c2c8ef61915f0e5f5718037d672a217bae93fb6ca8b6694be9bbce19fa183abc8427cfd8bcc1a4a7e5feca5641d4270d52938812c9b4e0b9f012d16b1ea363e7b697945b2ed4957a8c6d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68cc65ca7ddd49a2e13065b1d24fdaf034592cd9a9147f6ded1af20484de2e3239a26338e33ef67dbbfdde3395c8fdbddcbb8e17f3ca5cb6b335c9b86b17f4edd0a9c6b38aaf0bc364bda45e6d6a0c36a3e733e284479b414154c6917ffe6153684c92b65d17367414f83b0db55e2c54b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22b8c7e8b1c751780bb7b6ccde793efca26aab8f8ba98d31dc4feb17cfaec0bd0edc62e92a892cb94f01cab39af16738d96d1a8363548bccf63b89f1b92771714ae350480c7470ee099f109769129819b910f9c1315f8120057bdbb0a29fde693d2ae0590d38ef50c3237741d15277bd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebce1d3b9f305c7c5ae8996c1b9a020de1d2c1a6526c7579ba336213fe66d42ccaa12b49e08f838e44361ca771fd8fca5aef0b62daa6ca6277e90a75e73a28140e8b60b8dad94d046c45bf502cf951a9bd4f6c596a4b43ad4d48365fbc83638b9d38ab8131f1744466c507a2360f9f001;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb01f6d3b67d0942e3931a6373faf59cc1036875b2bb795a21d489530bc2fee4a8f7637628157148560a609b3d106d09f41b11d6901f0b8ab6fa336ca71a4d804cb6978ccb2529be9fa364f245d3dce70edbd0e170908a52b3a8d382cd769f4cfa1dcaa64361a337db7add310aff260fa1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6df07bf0a71188e9af7c3ba021e105f3a6e99133c7f70c5d53b1d3ede2696e45b733c3d8e444235637f9a4574626540990a6921fdeae446dafca9eb2849bd5221c80eff9d917ef2bf5b921a4fa0469160ef35bbe0967fda2f9c2d2b7abbf29fd3e2e4d386bac4ceee792bd3ec7f0c3698;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17a610602225b73caccc90a5f30757f741d20a6afb580202922de61a5f4fab26afb3edd74269b2d6974b92fd196271e181c3fac7dfd745f95ba25ece07bce2d454a62d20e69e905f6a5f290a18fb22e5ac436a15dc444ad192491eb1033683a29c609281d4da871afd7dc63af51e9c607;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac88b20143e7f2633f4985d6a18815b5ceb5181548e6ad625c3bb1b61541acb8ab5241e42ac607ee8014a03f55a3c3b389f39a3c2a83cc872f47a3abe3a43f933c0a3a5910f78b67822e6fecf7db0b72e322d1d6366193234a7c3a8d837df4a6d520c5889751a71e6c833bf1fef6231a3;
        #1
        $finish();
    end
endmodule
