module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    reg [31:0] src32;
    reg [31:0] src33;
    reg [31:0] src34;
    reg [31:0] src35;
    reg [31:0] src36;
    reg [31:0] src37;
    reg [31:0] src38;
    reg [31:0] src39;
    reg [31:0] src40;
    reg [31:0] src41;
    reg [31:0] src42;
    reg [31:0] src43;
    reg [31:0] src44;
    reg [31:0] src45;
    reg [31:0] src46;
    reg [31:0] src47;
    reg [31:0] src48;
    reg [31:0] src49;
    reg [31:0] src50;
    reg [31:0] src51;
    reg [31:0] src52;
    reg [31:0] src53;
    reg [31:0] src54;
    reg [31:0] src55;
    reg [31:0] src56;
    reg [31:0] src57;
    reg [31:0] src58;
    reg [31:0] src59;
    reg [31:0] src60;
    reg [31:0] src61;
    reg [31:0] src62;
    reg [31:0] src63;
    compressor_CLA32_64 compressor_CLA32_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
        src16 <= 32'h0;
        src17 <= 32'h0;
        src18 <= 32'h0;
        src19 <= 32'h0;
        src20 <= 32'h0;
        src21 <= 32'h0;
        src22 <= 32'h0;
        src23 <= 32'h0;
        src24 <= 32'h0;
        src25 <= 32'h0;
        src26 <= 32'h0;
        src27 <= 32'h0;
        src28 <= 32'h0;
        src29 <= 32'h0;
        src30 <= 32'h0;
        src31 <= 32'h0;
        src32 <= 32'h0;
        src33 <= 32'h0;
        src34 <= 32'h0;
        src35 <= 32'h0;
        src36 <= 32'h0;
        src37 <= 32'h0;
        src38 <= 32'h0;
        src39 <= 32'h0;
        src40 <= 32'h0;
        src41 <= 32'h0;
        src42 <= 32'h0;
        src43 <= 32'h0;
        src44 <= 32'h0;
        src45 <= 32'h0;
        src46 <= 32'h0;
        src47 <= 32'h0;
        src48 <= 32'h0;
        src49 <= 32'h0;
        src50 <= 32'h0;
        src51 <= 32'h0;
        src52 <= 32'h0;
        src53 <= 32'h0;
        src54 <= 32'h0;
        src55 <= 32'h0;
        src56 <= 32'h0;
        src57 <= 32'h0;
        src58 <= 32'h0;
        src59 <= 32'h0;
        src60 <= 32'h0;
        src61 <= 32'h0;
        src62 <= 32'h0;
        src63 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA32_64(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    input [31:0]src16,
    input [31:0]src17,
    input [31:0]src18,
    input [31:0]src19,
    input [31:0]src20,
    input [31:0]src21,
    input [31:0]src22,
    input [31:0]src23,
    input [31:0]src24,
    input [31:0]src25,
    input [31:0]src26,
    input [31:0]src27,
    input [31:0]src28,
    input [31:0]src29,
    input [31:0]src30,
    input [31:0]src31,
    input [31:0]src32,
    input [31:0]src33,
    input [31:0]src34,
    input [31:0]src35,
    input [31:0]src36,
    input [31:0]src37,
    input [31:0]src38,
    input [31:0]src39,
    input [31:0]src40,
    input [31:0]src41,
    input [31:0]src42,
    input [31:0]src43,
    input [31:0]src44,
    input [31:0]src45,
    input [31:0]src46,
    input [31:0]src47,
    input [31:0]src48,
    input [31:0]src49,
    input [31:0]src50,
    input [31:0]src51,
    input [31:0]src52,
    input [31:0]src53,
    input [31:0]src54,
    input [31:0]src55,
    input [31:0]src56,
    input [31:0]src57,
    input [31:0]src58,
    input [31:0]src59,
    input [31:0]src60,
    input [31:0]src61,
    input [31:0]src62,
    input [31:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [0:0] comp_out68;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      input wire [31:0] src32,
      input wire [31:0] src33,
      input wire [31:0] src34,
      input wire [31:0] src35,
      input wire [31:0] src36,
      input wire [31:0] src37,
      input wire [31:0] src38,
      input wire [31:0] src39,
      input wire [31:0] src40,
      input wire [31:0] src41,
      input wire [31:0] src42,
      input wire [31:0] src43,
      input wire [31:0] src44,
      input wire [31:0] src45,
      input wire [31:0] src46,
      input wire [31:0] src47,
      input wire [31:0] src48,
      input wire [31:0] src49,
      input wire [31:0] src50,
      input wire [31:0] src51,
      input wire [31:0] src52,
      input wire [31:0] src53,
      input wire [31:0] src54,
      input wire [31:0] src55,
      input wire [31:0] src56,
      input wire [31:0] src57,
      input wire [31:0] src58,
      input wire [31:0] src59,
      input wire [31:0] src60,
      input wire [31:0] src61,
      input wire [31:0] src62,
      input wire [31:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [0:0] dst68);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [31:0] stage0_16;
   wire [31:0] stage0_17;
   wire [31:0] stage0_18;
   wire [31:0] stage0_19;
   wire [31:0] stage0_20;
   wire [31:0] stage0_21;
   wire [31:0] stage0_22;
   wire [31:0] stage0_23;
   wire [31:0] stage0_24;
   wire [31:0] stage0_25;
   wire [31:0] stage0_26;
   wire [31:0] stage0_27;
   wire [31:0] stage0_28;
   wire [31:0] stage0_29;
   wire [31:0] stage0_30;
   wire [31:0] stage0_31;
   wire [31:0] stage0_32;
   wire [31:0] stage0_33;
   wire [31:0] stage0_34;
   wire [31:0] stage0_35;
   wire [31:0] stage0_36;
   wire [31:0] stage0_37;
   wire [31:0] stage0_38;
   wire [31:0] stage0_39;
   wire [31:0] stage0_40;
   wire [31:0] stage0_41;
   wire [31:0] stage0_42;
   wire [31:0] stage0_43;
   wire [31:0] stage0_44;
   wire [31:0] stage0_45;
   wire [31:0] stage0_46;
   wire [31:0] stage0_47;
   wire [31:0] stage0_48;
   wire [31:0] stage0_49;
   wire [31:0] stage0_50;
   wire [31:0] stage0_51;
   wire [31:0] stage0_52;
   wire [31:0] stage0_53;
   wire [31:0] stage0_54;
   wire [31:0] stage0_55;
   wire [31:0] stage0_56;
   wire [31:0] stage0_57;
   wire [31:0] stage0_58;
   wire [31:0] stage0_59;
   wire [31:0] stage0_60;
   wire [31:0] stage0_61;
   wire [31:0] stage0_62;
   wire [31:0] stage0_63;
   wire [10:0] stage1_0;
   wire [7:0] stage1_1;
   wire [24:0] stage1_2;
   wire [16:0] stage1_3;
   wire [29:0] stage1_4;
   wire [13:0] stage1_5;
   wire [28:0] stage1_6;
   wire [8:0] stage1_7;
   wire [18:0] stage1_8;
   wire [15:0] stage1_9;
   wire [17:0] stage1_10;
   wire [16:0] stage1_11;
   wire [18:0] stage1_12;
   wire [13:0] stage1_13;
   wire [16:0] stage1_14;
   wire [12:0] stage1_15;
   wire [30:0] stage1_16;
   wire [21:0] stage1_17;
   wire [10:0] stage1_18;
   wire [18:0] stage1_19;
   wire [11:0] stage1_20;
   wire [17:0] stage1_21;
   wire [13:0] stage1_22;
   wire [17:0] stage1_23;
   wire [11:0] stage1_24;
   wire [17:0] stage1_25;
   wire [16:0] stage1_26;
   wire [10:0] stage1_27;
   wire [15:0] stage1_28;
   wire [17:0] stage1_29;
   wire [10:0] stage1_30;
   wire [16:0] stage1_31;
   wire [24:0] stage1_32;
   wire [18:0] stage1_33;
   wire [20:0] stage1_34;
   wire [12:0] stage1_35;
   wire [12:0] stage1_36;
   wire [13:0] stage1_37;
   wire [17:0] stage1_38;
   wire [14:0] stage1_39;
   wire [15:0] stage1_40;
   wire [19:0] stage1_41;
   wire [12:0] stage1_42;
   wire [13:0] stage1_43;
   wire [13:0] stage1_44;
   wire [24:0] stage1_45;
   wire [11:0] stage1_46;
   wire [17:0] stage1_47;
   wire [19:0] stage1_48;
   wire [19:0] stage1_49;
   wire [11:0] stage1_50;
   wire [20:0] stage1_51;
   wire [11:0] stage1_52;
   wire [22:0] stage1_53;
   wire [9:0] stage1_54;
   wire [29:0] stage1_55;
   wire [14:0] stage1_56;
   wire [16:0] stage1_57;
   wire [13:0] stage1_58;
   wire [23:0] stage1_59;
   wire [12:0] stage1_60;
   wire [12:0] stage1_61;
   wire [16:0] stage1_62;
   wire [10:0] stage1_63;
   wire [8:0] stage1_64;
   wire [4:0] stage1_65;
   wire [10:0] stage2_0;
   wire [2:0] stage2_1;
   wire [8:0] stage2_2;
   wire [8:0] stage2_3;
   wire [6:0] stage2_4;
   wire [9:0] stage2_5;
   wire [17:0] stage2_6;
   wire [5:0] stage2_7;
   wire [5:0] stage2_8;
   wire [9:0] stage2_9;
   wire [7:0] stage2_10;
   wire [5:0] stage2_11;
   wire [5:0] stage2_12;
   wire [8:0] stage2_13;
   wire [11:0] stage2_14;
   wire [4:0] stage2_15;
   wire [11:0] stage2_16;
   wire [11:0] stage2_17;
   wire [7:0] stage2_18;
   wire [5:0] stage2_19;
   wire [7:0] stage2_20;
   wire [6:0] stage2_21;
   wire [9:0] stage2_22;
   wire [5:0] stage2_23;
   wire [7:0] stage2_24;
   wire [5:0] stage2_25;
   wire [5:0] stage2_26;
   wire [6:0] stage2_27;
   wire [8:0] stage2_28;
   wire [5:0] stage2_29;
   wire [5:0] stage2_30;
   wire [8:0] stage2_31;
   wire [7:0] stage2_32;
   wire [16:0] stage2_33;
   wire [6:0] stage2_34;
   wire [5:0] stage2_35;
   wire [7:0] stage2_36;
   wire [13:0] stage2_37;
   wire [4:0] stage2_38;
   wire [6:0] stage2_39;
   wire [5:0] stage2_40;
   wire [6:0] stage2_41;
   wire [10:0] stage2_42;
   wire [6:0] stage2_43;
   wire [17:0] stage2_44;
   wire [4:0] stage2_45;
   wire [7:0] stage2_46;
   wire [9:0] stage2_47;
   wire [6:0] stage2_48;
   wire [11:0] stage2_49;
   wire [6:0] stage2_50;
   wire [5:0] stage2_51;
   wire [5:0] stage2_52;
   wire [10:0] stage2_53;
   wire [6:0] stage2_54;
   wire [6:0] stage2_55;
   wire [9:0] stage2_56;
   wire [8:0] stage2_57;
   wire [5:0] stage2_58;
   wire [11:0] stage2_59;
   wire [6:0] stage2_60;
   wire [6:0] stage2_61;
   wire [5:0] stage2_62;
   wire [9:0] stage2_63;
   wire [4:0] stage2_64;
   wire [7:0] stage2_65;
   wire [0:0] stage2_66;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [3:0] stage3_2;
   wire [4:0] stage3_3;
   wire [4:0] stage3_4;
   wire [2:0] stage3_5;
   wire [5:0] stage3_6;
   wire [4:0] stage3_7;
   wire [2:0] stage3_8;
   wire [3:0] stage3_9;
   wire [5:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [4:0] stage3_13;
   wire [3:0] stage3_14;
   wire [3:0] stage3_15;
   wire [2:0] stage3_16;
   wire [3:0] stage3_17;
   wire [5:0] stage3_18;
   wire [2:0] stage3_19;
   wire [4:0] stage3_20;
   wire [2:0] stage3_21;
   wire [4:0] stage3_22;
   wire [2:0] stage3_23;
   wire [4:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [4:0] stage3_27;
   wire [4:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [3:0] stage3_31;
   wire [3:0] stage3_32;
   wire [3:0] stage3_33;
   wire [3:0] stage3_34;
   wire [3:0] stage3_35;
   wire [3:0] stage3_36;
   wire [3:0] stage3_37;
   wire [3:0] stage3_38;
   wire [3:0] stage3_39;
   wire [1:0] stage3_40;
   wire [2:0] stage3_41;
   wire [4:0] stage3_42;
   wire [3:0] stage3_43;
   wire [3:0] stage3_44;
   wire [3:0] stage3_45;
   wire [5:0] stage3_46;
   wire [4:0] stage3_47;
   wire [2:0] stage3_48;
   wire [2:0] stage3_49;
   wire [5:0] stage3_50;
   wire [3:0] stage3_51;
   wire [2:0] stage3_52;
   wire [2:0] stage3_53;
   wire [5:0] stage3_54;
   wire [2:0] stage3_55;
   wire [5:0] stage3_56;
   wire [2:0] stage3_57;
   wire [3:0] stage3_58;
   wire [5:0] stage3_59;
   wire [3:0] stage3_60;
   wire [2:0] stage3_61;
   wire [5:0] stage3_62;
   wire [2:0] stage3_63;
   wire [5:0] stage3_64;
   wire [3:0] stage3_65;
   wire [1:0] stage3_66;
   wire [0:0] stage3_67;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [1:0] stage4_33;
   wire [1:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage4_38;
   wire [1:0] stage4_39;
   wire [1:0] stage4_40;
   wire [1:0] stage4_41;
   wire [1:0] stage4_42;
   wire [1:0] stage4_43;
   wire [1:0] stage4_44;
   wire [1:0] stage4_45;
   wire [1:0] stage4_46;
   wire [1:0] stage4_47;
   wire [1:0] stage4_48;
   wire [1:0] stage4_49;
   wire [1:0] stage4_50;
   wire [1:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [1:0] stage4_54;
   wire [1:0] stage4_55;
   wire [1:0] stage4_56;
   wire [1:0] stage4_57;
   wire [1:0] stage4_58;
   wire [1:0] stage4_59;
   wire [1:0] stage4_60;
   wire [1:0] stage4_61;
   wire [1:0] stage4_62;
   wire [1:0] stage4_63;
   wire [1:0] stage4_64;
   wire [1:0] stage4_65;
   wire [1:0] stage4_66;
   wire [1:0] stage4_67;
   wire [0:0] stage4_68;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;
   assign dst37 = stage4_37;
   assign dst38 = stage4_38;
   assign dst39 = stage4_39;
   assign dst40 = stage4_40;
   assign dst41 = stage4_41;
   assign dst42 = stage4_42;
   assign dst43 = stage4_43;
   assign dst44 = stage4_44;
   assign dst45 = stage4_45;
   assign dst46 = stage4_46;
   assign dst47 = stage4_47;
   assign dst48 = stage4_48;
   assign dst49 = stage4_49;
   assign dst50 = stage4_50;
   assign dst51 = stage4_51;
   assign dst52 = stage4_52;
   assign dst53 = stage4_53;
   assign dst54 = stage4_54;
   assign dst55 = stage4_55;
   assign dst56 = stage4_56;
   assign dst57 = stage4_57;
   assign dst58 = stage4_58;
   assign dst59 = stage4_59;
   assign dst60 = stage4_60;
   assign dst61 = stage4_61;
   assign dst62 = stage4_62;
   assign dst63 = stage4_63;
   assign dst64 = stage4_64;
   assign dst65 = stage4_65;
   assign dst66 = stage4_66;
   assign dst67 = stage4_67;
   assign dst68 = stage4_68;

   gpc2116_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2116_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[0],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[1],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc615_5 gpc8 (
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15]},
      {stage0_3[19]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[9],stage1_3[9]}
   );
   gpc606_5 gpc10 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[10]}
   );
   gpc1343_5 gpc11 (
      {stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9]},
      {stage0_7[0], stage0_7[1], stage0_7[2]},
      {stage0_8[0]},
      {stage1_9[0],stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc12 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[1],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc606_5 gpc13 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[2],stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[7]}
   );
   gpc606_5 gpc14 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[3],stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[8]}
   );
   gpc615_5 gpc15 (
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25]},
      {stage0_8[1]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[4],stage1_8[5],stage1_7[6]}
   );
   gpc615_5 gpc16 (
      {stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30]},
      {stage0_8[2]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[1],stage1_9[5],stage1_8[6],stage1_7[7]}
   );
   gpc2135_5 gpc17 (
      {stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7]},
      {stage0_9[12], stage0_9[13], stage0_9[14]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[2],stage1_10[2],stage1_9[6],stage1_8[7]}
   );
   gpc606_5 gpc18 (
      {stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[1],stage1_11[3],stage1_10[3],stage1_9[7],stage1_8[8]}
   );
   gpc615_5 gpc19 (
      {stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_9[15]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[2],stage1_11[4],stage1_10[4],stage1_9[8],stage1_8[9]}
   );
   gpc615_5 gpc20 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[16]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[3],stage1_11[5],stage1_10[5],stage1_9[9],stage1_8[10]}
   );
   gpc606_5 gpc21 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[0],stage1_12[4],stage1_11[6],stage1_10[6],stage1_9[10]}
   );
   gpc623_5 gpc22 (
      {stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_10[19], stage0_10[20]},
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13]},
      {stage1_13[1],stage1_12[5],stage1_11[7],stage1_10[7],stage1_9[11]}
   );
   gpc623_5 gpc23 (
      {stage0_9[26], stage0_9[27], stage0_9[28]},
      {stage0_10[21], stage0_10[22]},
      {stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18], stage0_11[19]},
      {stage1_13[2],stage1_12[6],stage1_11[8],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc24 (
      {stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[3],stage1_12[7],stage1_11[9]}
   );
   gpc606_5 gpc25 (
      {stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[4],stage1_12[8]}
   );
   gpc606_5 gpc26 (
      {stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[5],stage1_12[9]}
   );
   gpc606_5 gpc27 (
      {stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc28 (
      {stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc29 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[8]}
   );
   gpc606_5 gpc30 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[9]}
   );
   gpc606_5 gpc31 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[10]}
   );
   gpc606_5 gpc32 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[11]}
   );
   gpc615_5 gpc33 (
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28]},
      {stage0_16[0]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[0],stage1_17[4],stage1_16[8],stage1_15[9]}
   );
   gpc606_5 gpc34 (
      {stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5], stage0_16[6]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[1],stage1_18[1],stage1_17[5],stage1_16[9]}
   );
   gpc615_5 gpc35 (
      {stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage0_17[6]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[2],stage1_18[2],stage1_17[6],stage1_16[10]}
   );
   gpc606_5 gpc36 (
      {stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11], stage0_17[12]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[2],stage1_19[3],stage1_18[3],stage1_17[7]}
   );
   gpc606_5 gpc37 (
      {stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17], stage0_17[18]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[3],stage1_19[4],stage1_18[4],stage1_17[8]}
   );
   gpc1406_5 gpc38 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3]},
      {stage0_21[0]},
      {stage1_22[0],stage1_21[2],stage1_20[4],stage1_19[5],stage1_18[5]}
   );
   gpc1406_5 gpc39 (
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage0_20[4], stage0_20[5], stage0_20[6], stage0_20[7]},
      {stage0_21[1]},
      {stage1_22[1],stage1_21[3],stage1_20[5],stage1_19[6],stage1_18[6]}
   );
   gpc615_5 gpc40 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28]},
      {stage0_19[12]},
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13]},
      {stage1_22[2],stage1_21[4],stage1_20[6],stage1_19[7],stage1_18[7]}
   );
   gpc615_5 gpc41 (
      {stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage0_20[14]},
      {stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7]},
      {stage1_23[0],stage1_22[3],stage1_21[5],stage1_20[7],stage1_19[8]}
   );
   gpc615_5 gpc42 (
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22]},
      {stage0_20[15]},
      {stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13]},
      {stage1_23[1],stage1_22[4],stage1_21[6],stage1_20[8],stage1_19[9]}
   );
   gpc606_5 gpc43 (
      {stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[5],stage1_21[7],stage1_20[9]}
   );
   gpc606_5 gpc44 (
      {stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[6],stage1_21[8],stage1_20[10]}
   );
   gpc606_5 gpc45 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], 1'b0, 1'b0},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[7],stage1_21[9],stage1_20[11]}
   );
   gpc606_5 gpc46 (
      {stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[3],stage1_23[5],stage1_22[8],stage1_21[10]}
   );
   gpc606_5 gpc47 (
      {stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[4],stage1_23[6],stage1_22[9],stage1_21[11]}
   );
   gpc1163_5 gpc48 (
      {stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage0_24[0]},
      {stage0_25[0]},
      {stage1_26[0],stage1_25[2],stage1_24[5],stage1_23[7],stage1_22[10]}
   );
   gpc615_5 gpc49 (
      {stage0_22[21], stage0_22[22], stage0_22[23], stage0_22[24], stage0_22[25]},
      {stage0_23[18]},
      {stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6]},
      {stage1_26[1],stage1_25[3],stage1_24[6],stage1_23[8],stage1_22[11]}
   );
   gpc615_5 gpc50 (
      {stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30]},
      {stage0_23[19]},
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage1_26[2],stage1_25[4],stage1_24[7],stage1_23[9],stage1_22[12]}
   );
   gpc615_5 gpc51 (
      {stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24]},
      {stage0_24[13]},
      {stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5], stage0_25[6]},
      {stage1_27[0],stage1_26[3],stage1_25[5],stage1_24[8],stage1_23[10]}
   );
   gpc606_5 gpc52 (
      {stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18], stage0_24[19]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[4],stage1_25[6],stage1_24[9]}
   );
   gpc606_5 gpc53 (
      {stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24], stage0_24[25]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[5],stage1_25[7],stage1_24[10]}
   );
   gpc606_5 gpc54 (
      {stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[3],stage1_26[6],stage1_25[8],stage1_24[11]}
   );
   gpc615_5 gpc55 (
      {stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage0_26[18]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[3],stage1_27[4],stage1_26[7],stage1_25[9]}
   );
   gpc615_5 gpc56 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16]},
      {stage0_26[19]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[4],stage1_27[5],stage1_26[8],stage1_25[10]}
   );
   gpc615_5 gpc57 (
      {stage0_25[17], stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21]},
      {stage0_26[20]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[5],stage1_27[6],stage1_26[9],stage1_25[11]}
   );
   gpc615_5 gpc58 (
      {stage0_25[22], stage0_25[23], stage0_25[24], stage0_25[25], stage0_25[26]},
      {stage0_26[21]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[6],stage1_27[7],stage1_26[10],stage1_25[12]}
   );
   gpc615_5 gpc59 (
      {stage0_26[22], stage0_26[23], stage0_26[24], stage0_26[25], stage0_26[26]},
      {stage0_27[24]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[4],stage1_28[7],stage1_27[8],stage1_26[11]}
   );
   gpc606_5 gpc60 (
      {stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29], stage0_27[30]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[5],stage1_28[8],stage1_27[9]}
   );
   gpc606_5 gpc61 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[1],stage1_30[2],stage1_29[6],stage1_28[9]}
   );
   gpc606_5 gpc62 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[2],stage1_30[3],stage1_29[7],stage1_28[10]}
   );
   gpc606_5 gpc63 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[3],stage1_30[4],stage1_29[8],stage1_28[11]}
   );
   gpc615_5 gpc64 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28]},
      {stage0_29[6]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[4],stage1_30[5],stage1_29[9],stage1_28[12]}
   );
   gpc606_5 gpc65 (
      {stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[4],stage1_31[5],stage1_30[6],stage1_29[10]}
   );
   gpc615_5 gpc66 (
      {stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_30[24]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[5],stage1_31[6],stage1_30[7],stage1_29[11]}
   );
   gpc615_5 gpc67 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22]},
      {stage0_30[25]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[6],stage1_31[7],stage1_30[8],stage1_29[12]}
   );
   gpc615_5 gpc68 (
      {stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27]},
      {stage0_30[26]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[7],stage1_31[8],stage1_30[9],stage1_29[13]}
   );
   gpc615_5 gpc69 (
      {stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30], stage0_30[31]},
      {stage0_31[24]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[4],stage1_32[8],stage1_31[9],stage1_30[10]}
   );
   gpc606_5 gpc70 (
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[0],stage1_34[1],stage1_33[5],stage1_32[9]}
   );
   gpc606_5 gpc71 (
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[1],stage1_34[2],stage1_33[6],stage1_32[10]}
   );
   gpc606_5 gpc72 (
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[2],stage1_35[2],stage1_34[3],stage1_33[7]}
   );
   gpc606_5 gpc73 (
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[3],stage1_35[3],stage1_34[4],stage1_33[8]}
   );
   gpc606_5 gpc74 (
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[4],stage1_35[4],stage1_34[5],stage1_33[9]}
   );
   gpc606_5 gpc75 (
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[5],stage1_35[5],stage1_34[6],stage1_33[10]}
   );
   gpc615_5 gpc76 (
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16]},
      {stage0_35[24]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[4],stage1_36[6],stage1_35[6],stage1_34[7]}
   );
   gpc623_5 gpc77 (
      {stage0_34[17], stage0_34[18], stage0_34[19]},
      {stage0_35[25], stage0_35[26]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[5],stage1_36[7],stage1_35[7],stage1_34[8]}
   );
   gpc606_5 gpc78 (
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[0],stage1_38[2],stage1_37[6],stage1_36[8]}
   );
   gpc606_5 gpc79 (
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[1],stage1_38[3],stage1_37[7],stage1_36[9]}
   );
   gpc606_5 gpc80 (
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[2],stage1_38[4],stage1_37[8],stage1_36[10]}
   );
   gpc117_4 gpc81 (
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5], stage0_37[6]},
      {stage0_38[18]},
      {stage0_39[0]},
      {stage1_40[3],stage1_39[3],stage1_38[5],stage1_37[9]}
   );
   gpc117_4 gpc82 (
      {stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12], stage0_37[13]},
      {stage0_38[19]},
      {stage0_39[1]},
      {stage1_40[4],stage1_39[4],stage1_38[6],stage1_37[10]}
   );
   gpc606_5 gpc83 (
      {stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17], stage0_37[18], stage0_37[19]},
      {stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5], stage0_39[6], stage0_39[7]},
      {stage1_41[0],stage1_40[5],stage1_39[5],stage1_38[7],stage1_37[11]}
   );
   gpc606_5 gpc84 (
      {stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23], stage0_37[24], stage0_37[25]},
      {stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11], stage0_39[12], stage0_39[13]},
      {stage1_41[1],stage1_40[6],stage1_39[6],stage1_38[8],stage1_37[12]}
   );
   gpc606_5 gpc85 (
      {stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29], stage0_37[30], stage0_37[31]},
      {stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17], stage0_39[18], stage0_39[19]},
      {stage1_41[2],stage1_40[7],stage1_39[7],stage1_38[9],stage1_37[13]}
   );
   gpc615_5 gpc86 (
      {stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23], stage0_38[24]},
      {stage0_39[20]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[3],stage1_40[8],stage1_39[8],stage1_38[10]}
   );
   gpc606_5 gpc87 (
      {stage0_39[21], stage0_39[22], stage0_39[23], stage0_39[24], stage0_39[25], stage0_39[26]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[4],stage1_40[9],stage1_39[9]}
   );
   gpc606_5 gpc88 (
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[1],stage1_42[2],stage1_41[5],stage1_40[10]}
   );
   gpc606_5 gpc89 (
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[2],stage1_42[3],stage1_41[6],stage1_40[11]}
   );
   gpc606_5 gpc90 (
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[3],stage1_42[4],stage1_41[7],stage1_40[12]}
   );
   gpc606_5 gpc91 (
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[4],stage1_42[5],stage1_41[8],stage1_40[13]}
   );
   gpc606_5 gpc92 (
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[4],stage1_43[5],stage1_42[6],stage1_41[9]}
   );
   gpc606_5 gpc93 (
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[5],stage1_43[6],stage1_42[7],stage1_41[10]}
   );
   gpc606_5 gpc94 (
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[6],stage1_43[7],stage1_42[8],stage1_41[11]}
   );
   gpc615_5 gpc95 (
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28]},
      {stage0_43[18]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[3],stage1_44[7],stage1_43[8],stage1_42[9]}
   );
   gpc615_5 gpc96 (
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage0_44[6]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[1],stage1_45[4],stage1_44[8],stage1_43[9]}
   );
   gpc615_5 gpc97 (
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28]},
      {stage0_44[7]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[2],stage1_45[5],stage1_44[9],stage1_43[10]}
   );
   gpc606_5 gpc98 (
      {stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11], stage0_44[12], stage0_44[13]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[2],stage1_46[3],stage1_45[6],stage1_44[10]}
   );
   gpc606_5 gpc99 (
      {stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17], stage0_44[18], stage0_44[19]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[3],stage1_46[4],stage1_45[7],stage1_44[11]}
   );
   gpc606_5 gpc100 (
      {stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23], stage0_44[24], stage0_44[25]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[4],stage1_46[5],stage1_45[8],stage1_44[12]}
   );
   gpc606_5 gpc101 (
      {stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29], stage0_44[30], stage0_44[31]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[5],stage1_46[6],stage1_45[9],stage1_44[13]}
   );
   gpc606_5 gpc102 (
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[4],stage1_47[6],stage1_46[7],stage1_45[10]}
   );
   gpc615_5 gpc103 (
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28]},
      {stage0_47[6]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[1],stage1_48[5],stage1_47[7],stage1_46[8]}
   );
   gpc606_5 gpc104 (
      {stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11], stage0_47[12]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[1],stage1_49[2],stage1_48[6],stage1_47[8]}
   );
   gpc606_5 gpc105 (
      {stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17], stage0_47[18]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[2],stage1_49[3],stage1_48[7],stage1_47[9]}
   );
   gpc606_5 gpc106 (
      {stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[3],stage1_49[4],stage1_48[8],stage1_47[10]}
   );
   gpc606_5 gpc107 (
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[3],stage1_50[4],stage1_49[5],stage1_48[9]}
   );
   gpc606_5 gpc108 (
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[4],stage1_50[5],stage1_49[6],stage1_48[10]}
   );
   gpc606_5 gpc109 (
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[5],stage1_50[6],stage1_49[7],stage1_48[11]}
   );
   gpc623_5 gpc110 (
      {stage0_49[18], stage0_49[19], stage0_49[20]},
      {stage0_50[18], stage0_50[19]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[3],stage1_51[6],stage1_50[7],stage1_49[8]}
   );
   gpc615_5 gpc111 (
      {stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23], stage0_50[24]},
      {stage0_51[6]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[1],stage1_52[4],stage1_51[7],stage1_50[8]}
   );
   gpc615_5 gpc112 (
      {stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage0_51[7]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[2],stage1_52[5],stage1_51[8],stage1_50[9]}
   );
   gpc615_5 gpc113 (
      {stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11], stage0_51[12]},
      {stage0_52[12]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[2],stage1_53[3],stage1_52[6],stage1_51[9]}
   );
   gpc615_5 gpc114 (
      {stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage0_52[13]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[3],stage1_53[4],stage1_52[7],stage1_51[10]}
   );
   gpc615_5 gpc115 (
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22]},
      {stage0_52[14]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[4],stage1_53[5],stage1_52[8],stage1_51[11]}
   );
   gpc606_5 gpc116 (
      {stage0_52[15], stage0_52[16], stage0_52[17], stage0_52[18], stage0_52[19], stage0_52[20]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[3],stage1_54[5],stage1_53[6],stage1_52[9]}
   );
   gpc606_5 gpc117 (
      {stage0_52[21], stage0_52[22], stage0_52[23], stage0_52[24], stage0_52[25], stage0_52[26]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[4],stage1_54[6],stage1_53[7],stage1_52[10]}
   );
   gpc606_5 gpc118 (
      {stage0_52[27], stage0_52[28], stage0_52[29], stage0_52[30], stage0_52[31], 1'b0},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[5],stage1_54[7],stage1_53[8],stage1_52[11]}
   );
   gpc207_4 gpc119 (
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23], stage0_54[24]},
      {stage0_56[0], stage0_56[1]},
      {stage1_57[0],stage1_56[3],stage1_55[6],stage1_54[8]}
   );
   gpc207_4 gpc120 (
      {stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29], stage0_54[30], stage0_54[31]},
      {stage0_56[2], stage0_56[3]},
      {stage1_57[1],stage1_56[4],stage1_55[7],stage1_54[9]}
   );
   gpc1163_5 gpc121 (
      {stage0_55[0], stage0_55[1], stage0_55[2]},
      {stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9]},
      {stage0_57[0]},
      {stage0_58[0]},
      {stage1_59[0],stage1_58[0],stage1_57[2],stage1_56[5],stage1_55[8]}
   );
   gpc615_5 gpc122 (
      {stage0_55[3], stage0_55[4], stage0_55[5], stage0_55[6], stage0_55[7]},
      {stage0_56[10]},
      {stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6]},
      {stage1_59[1],stage1_58[1],stage1_57[3],stage1_56[6],stage1_55[9]}
   );
   gpc615_5 gpc123 (
      {stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11], stage0_55[12]},
      {stage0_56[11]},
      {stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11], stage0_57[12]},
      {stage1_59[2],stage1_58[2],stage1_57[4],stage1_56[7],stage1_55[10]}
   );
   gpc606_5 gpc124 (
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5], stage0_58[6]},
      {stage1_60[0],stage1_59[3],stage1_58[3],stage1_57[5],stage1_56[8]}
   );
   gpc615_5 gpc125 (
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22]},
      {stage0_57[13]},
      {stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11], stage0_58[12]},
      {stage1_60[1],stage1_59[4],stage1_58[4],stage1_57[6],stage1_56[9]}
   );
   gpc615_5 gpc126 (
      {stage0_56[23], stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27]},
      {stage0_57[14]},
      {stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17], stage0_58[18]},
      {stage1_60[2],stage1_59[5],stage1_58[5],stage1_57[7],stage1_56[10]}
   );
   gpc615_5 gpc127 (
      {stage0_57[15], stage0_57[16], stage0_57[17], stage0_57[18], stage0_57[19]},
      {stage0_58[19]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[3],stage1_59[6],stage1_58[6],stage1_57[8]}
   );
   gpc615_5 gpc128 (
      {stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23], stage0_57[24]},
      {stage0_58[20]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[4],stage1_59[7],stage1_58[7],stage1_57[9]}
   );
   gpc606_5 gpc129 (
      {stage0_58[21], stage0_58[22], stage0_58[23], stage0_58[24], stage0_58[25], stage0_58[26]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[2],stage1_60[5],stage1_59[8],stage1_58[8]}
   );
   gpc606_5 gpc130 (
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[1],stage1_61[3],stage1_60[6],stage1_59[9]}
   );
   gpc1406_5 gpc131 (
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3]},
      {stage0_63[0]},
      {stage1_64[0],stage1_63[1],stage1_62[2],stage1_61[4],stage1_60[7]}
   );
   gpc606_5 gpc132 (
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage0_62[4], stage0_62[5], stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9]},
      {stage1_64[1],stage1_63[2],stage1_62[3],stage1_61[5],stage1_60[8]}
   );
   gpc606_5 gpc133 (
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage0_62[10], stage0_62[11], stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15]},
      {stage1_64[2],stage1_63[3],stage1_62[4],stage1_61[6],stage1_60[9]}
   );
   gpc606_5 gpc134 (
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage0_62[16], stage0_62[17], stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21]},
      {stage1_64[3],stage1_63[4],stage1_62[5],stage1_61[7],stage1_60[10]}
   );
   gpc606_5 gpc135 (
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5], stage0_63[6]},
      {stage1_65[0],stage1_64[4],stage1_63[5],stage1_62[6],stage1_61[8]}
   );
   gpc615_5 gpc136 (
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16]},
      {stage0_62[22]},
      {stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11], stage0_63[12]},
      {stage1_65[1],stage1_64[5],stage1_63[6],stage1_62[7],stage1_61[9]}
   );
   gpc615_5 gpc137 (
      {stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21]},
      {stage0_62[23]},
      {stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17], stage0_63[18]},
      {stage1_65[2],stage1_64[6],stage1_63[7],stage1_62[8],stage1_61[10]}
   );
   gpc615_5 gpc138 (
      {stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26]},
      {stage0_62[24]},
      {stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23], stage0_63[24]},
      {stage1_65[3],stage1_64[7],stage1_63[8],stage1_62[9],stage1_61[11]}
   );
   gpc615_5 gpc139 (
      {stage0_61[27], stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31]},
      {stage0_62[25]},
      {stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29], stage0_63[30]},
      {stage1_65[4],stage1_64[8],stage1_63[9],stage1_62[10],stage1_61[12]}
   );
   gpc1_1 gpc140 (
      {stage0_0[27]},
      {stage1_0[6]}
   );
   gpc1_1 gpc141 (
      {stage0_0[28]},
      {stage1_0[7]}
   );
   gpc1_1 gpc142 (
      {stage0_0[29]},
      {stage1_0[8]}
   );
   gpc1_1 gpc143 (
      {stage0_0[30]},
      {stage1_0[9]}
   );
   gpc1_1 gpc144 (
      {stage0_0[31]},
      {stage1_0[10]}
   );
   gpc1_1 gpc145 (
      {stage0_2[16]},
      {stage1_2[9]}
   );
   gpc1_1 gpc146 (
      {stage0_2[17]},
      {stage1_2[10]}
   );
   gpc1_1 gpc147 (
      {stage0_2[18]},
      {stage1_2[11]}
   );
   gpc1_1 gpc148 (
      {stage0_2[19]},
      {stage1_2[12]}
   );
   gpc1_1 gpc149 (
      {stage0_2[20]},
      {stage1_2[13]}
   );
   gpc1_1 gpc150 (
      {stage0_2[21]},
      {stage1_2[14]}
   );
   gpc1_1 gpc151 (
      {stage0_2[22]},
      {stage1_2[15]}
   );
   gpc1_1 gpc152 (
      {stage0_2[23]},
      {stage1_2[16]}
   );
   gpc1_1 gpc153 (
      {stage0_2[24]},
      {stage1_2[17]}
   );
   gpc1_1 gpc154 (
      {stage0_2[25]},
      {stage1_2[18]}
   );
   gpc1_1 gpc155 (
      {stage0_2[26]},
      {stage1_2[19]}
   );
   gpc1_1 gpc156 (
      {stage0_2[27]},
      {stage1_2[20]}
   );
   gpc1_1 gpc157 (
      {stage0_2[28]},
      {stage1_2[21]}
   );
   gpc1_1 gpc158 (
      {stage0_2[29]},
      {stage1_2[22]}
   );
   gpc1_1 gpc159 (
      {stage0_2[30]},
      {stage1_2[23]}
   );
   gpc1_1 gpc160 (
      {stage0_2[31]},
      {stage1_2[24]}
   );
   gpc1_1 gpc161 (
      {stage0_3[25]},
      {stage1_3[10]}
   );
   gpc1_1 gpc162 (
      {stage0_3[26]},
      {stage1_3[11]}
   );
   gpc1_1 gpc163 (
      {stage0_3[27]},
      {stage1_3[12]}
   );
   gpc1_1 gpc164 (
      {stage0_3[28]},
      {stage1_3[13]}
   );
   gpc1_1 gpc165 (
      {stage0_3[29]},
      {stage1_3[14]}
   );
   gpc1_1 gpc166 (
      {stage0_3[30]},
      {stage1_3[15]}
   );
   gpc1_1 gpc167 (
      {stage0_3[31]},
      {stage1_3[16]}
   );
   gpc1_1 gpc168 (
      {stage0_4[13]},
      {stage1_4[11]}
   );
   gpc1_1 gpc169 (
      {stage0_4[14]},
      {stage1_4[12]}
   );
   gpc1_1 gpc170 (
      {stage0_4[15]},
      {stage1_4[13]}
   );
   gpc1_1 gpc171 (
      {stage0_4[16]},
      {stage1_4[14]}
   );
   gpc1_1 gpc172 (
      {stage0_4[17]},
      {stage1_4[15]}
   );
   gpc1_1 gpc173 (
      {stage0_4[18]},
      {stage1_4[16]}
   );
   gpc1_1 gpc174 (
      {stage0_4[19]},
      {stage1_4[17]}
   );
   gpc1_1 gpc175 (
      {stage0_4[20]},
      {stage1_4[18]}
   );
   gpc1_1 gpc176 (
      {stage0_4[21]},
      {stage1_4[19]}
   );
   gpc1_1 gpc177 (
      {stage0_4[22]},
      {stage1_4[20]}
   );
   gpc1_1 gpc178 (
      {stage0_4[23]},
      {stage1_4[21]}
   );
   gpc1_1 gpc179 (
      {stage0_4[24]},
      {stage1_4[22]}
   );
   gpc1_1 gpc180 (
      {stage0_4[25]},
      {stage1_4[23]}
   );
   gpc1_1 gpc181 (
      {stage0_4[26]},
      {stage1_4[24]}
   );
   gpc1_1 gpc182 (
      {stage0_4[27]},
      {stage1_4[25]}
   );
   gpc1_1 gpc183 (
      {stage0_4[28]},
      {stage1_4[26]}
   );
   gpc1_1 gpc184 (
      {stage0_4[29]},
      {stage1_4[27]}
   );
   gpc1_1 gpc185 (
      {stage0_4[30]},
      {stage1_4[28]}
   );
   gpc1_1 gpc186 (
      {stage0_4[31]},
      {stage1_4[29]}
   );
   gpc1_1 gpc187 (
      {stage0_5[27]},
      {stage1_5[9]}
   );
   gpc1_1 gpc188 (
      {stage0_5[28]},
      {stage1_5[10]}
   );
   gpc1_1 gpc189 (
      {stage0_5[29]},
      {stage1_5[11]}
   );
   gpc1_1 gpc190 (
      {stage0_5[30]},
      {stage1_5[12]}
   );
   gpc1_1 gpc191 (
      {stage0_5[31]},
      {stage1_5[13]}
   );
   gpc1_1 gpc192 (
      {stage0_6[10]},
      {stage1_6[7]}
   );
   gpc1_1 gpc193 (
      {stage0_6[11]},
      {stage1_6[8]}
   );
   gpc1_1 gpc194 (
      {stage0_6[12]},
      {stage1_6[9]}
   );
   gpc1_1 gpc195 (
      {stage0_6[13]},
      {stage1_6[10]}
   );
   gpc1_1 gpc196 (
      {stage0_6[14]},
      {stage1_6[11]}
   );
   gpc1_1 gpc197 (
      {stage0_6[15]},
      {stage1_6[12]}
   );
   gpc1_1 gpc198 (
      {stage0_6[16]},
      {stage1_6[13]}
   );
   gpc1_1 gpc199 (
      {stage0_6[17]},
      {stage1_6[14]}
   );
   gpc1_1 gpc200 (
      {stage0_6[18]},
      {stage1_6[15]}
   );
   gpc1_1 gpc201 (
      {stage0_6[19]},
      {stage1_6[16]}
   );
   gpc1_1 gpc202 (
      {stage0_6[20]},
      {stage1_6[17]}
   );
   gpc1_1 gpc203 (
      {stage0_6[21]},
      {stage1_6[18]}
   );
   gpc1_1 gpc204 (
      {stage0_6[22]},
      {stage1_6[19]}
   );
   gpc1_1 gpc205 (
      {stage0_6[23]},
      {stage1_6[20]}
   );
   gpc1_1 gpc206 (
      {stage0_6[24]},
      {stage1_6[21]}
   );
   gpc1_1 gpc207 (
      {stage0_6[25]},
      {stage1_6[22]}
   );
   gpc1_1 gpc208 (
      {stage0_6[26]},
      {stage1_6[23]}
   );
   gpc1_1 gpc209 (
      {stage0_6[27]},
      {stage1_6[24]}
   );
   gpc1_1 gpc210 (
      {stage0_6[28]},
      {stage1_6[25]}
   );
   gpc1_1 gpc211 (
      {stage0_6[29]},
      {stage1_6[26]}
   );
   gpc1_1 gpc212 (
      {stage0_6[30]},
      {stage1_6[27]}
   );
   gpc1_1 gpc213 (
      {stage0_6[31]},
      {stage1_6[28]}
   );
   gpc1_1 gpc214 (
      {stage0_7[31]},
      {stage1_7[8]}
   );
   gpc1_1 gpc215 (
      {stage0_8[24]},
      {stage1_8[11]}
   );
   gpc1_1 gpc216 (
      {stage0_8[25]},
      {stage1_8[12]}
   );
   gpc1_1 gpc217 (
      {stage0_8[26]},
      {stage1_8[13]}
   );
   gpc1_1 gpc218 (
      {stage0_8[27]},
      {stage1_8[14]}
   );
   gpc1_1 gpc219 (
      {stage0_8[28]},
      {stage1_8[15]}
   );
   gpc1_1 gpc220 (
      {stage0_8[29]},
      {stage1_8[16]}
   );
   gpc1_1 gpc221 (
      {stage0_8[30]},
      {stage1_8[17]}
   );
   gpc1_1 gpc222 (
      {stage0_8[31]},
      {stage1_8[18]}
   );
   gpc1_1 gpc223 (
      {stage0_9[29]},
      {stage1_9[13]}
   );
   gpc1_1 gpc224 (
      {stage0_9[30]},
      {stage1_9[14]}
   );
   gpc1_1 gpc225 (
      {stage0_9[31]},
      {stage1_9[15]}
   );
   gpc1_1 gpc226 (
      {stage0_10[23]},
      {stage1_10[9]}
   );
   gpc1_1 gpc227 (
      {stage0_10[24]},
      {stage1_10[10]}
   );
   gpc1_1 gpc228 (
      {stage0_10[25]},
      {stage1_10[11]}
   );
   gpc1_1 gpc229 (
      {stage0_10[26]},
      {stage1_10[12]}
   );
   gpc1_1 gpc230 (
      {stage0_10[27]},
      {stage1_10[13]}
   );
   gpc1_1 gpc231 (
      {stage0_10[28]},
      {stage1_10[14]}
   );
   gpc1_1 gpc232 (
      {stage0_10[29]},
      {stage1_10[15]}
   );
   gpc1_1 gpc233 (
      {stage0_10[30]},
      {stage1_10[16]}
   );
   gpc1_1 gpc234 (
      {stage0_10[31]},
      {stage1_10[17]}
   );
   gpc1_1 gpc235 (
      {stage0_11[25]},
      {stage1_11[10]}
   );
   gpc1_1 gpc236 (
      {stage0_11[26]},
      {stage1_11[11]}
   );
   gpc1_1 gpc237 (
      {stage0_11[27]},
      {stage1_11[12]}
   );
   gpc1_1 gpc238 (
      {stage0_11[28]},
      {stage1_11[13]}
   );
   gpc1_1 gpc239 (
      {stage0_11[29]},
      {stage1_11[14]}
   );
   gpc1_1 gpc240 (
      {stage0_11[30]},
      {stage1_11[15]}
   );
   gpc1_1 gpc241 (
      {stage0_11[31]},
      {stage1_11[16]}
   );
   gpc1_1 gpc242 (
      {stage0_12[25]},
      {stage1_12[12]}
   );
   gpc1_1 gpc243 (
      {stage0_12[26]},
      {stage1_12[13]}
   );
   gpc1_1 gpc244 (
      {stage0_12[27]},
      {stage1_12[14]}
   );
   gpc1_1 gpc245 (
      {stage0_12[28]},
      {stage1_12[15]}
   );
   gpc1_1 gpc246 (
      {stage0_12[29]},
      {stage1_12[16]}
   );
   gpc1_1 gpc247 (
      {stage0_12[30]},
      {stage1_12[17]}
   );
   gpc1_1 gpc248 (
      {stage0_12[31]},
      {stage1_12[18]}
   );
   gpc1_1 gpc249 (
      {stage0_13[30]},
      {stage1_13[12]}
   );
   gpc1_1 gpc250 (
      {stage0_13[31]},
      {stage1_13[13]}
   );
   gpc1_1 gpc251 (
      {stage0_14[24]},
      {stage1_14[9]}
   );
   gpc1_1 gpc252 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc253 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc254 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc255 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc256 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc257 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc258 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc259 (
      {stage0_15[29]},
      {stage1_15[10]}
   );
   gpc1_1 gpc260 (
      {stage0_15[30]},
      {stage1_15[11]}
   );
   gpc1_1 gpc261 (
      {stage0_15[31]},
      {stage1_15[12]}
   );
   gpc1_1 gpc262 (
      {stage0_16[12]},
      {stage1_16[11]}
   );
   gpc1_1 gpc263 (
      {stage0_16[13]},
      {stage1_16[12]}
   );
   gpc1_1 gpc264 (
      {stage0_16[14]},
      {stage1_16[13]}
   );
   gpc1_1 gpc265 (
      {stage0_16[15]},
      {stage1_16[14]}
   );
   gpc1_1 gpc266 (
      {stage0_16[16]},
      {stage1_16[15]}
   );
   gpc1_1 gpc267 (
      {stage0_16[17]},
      {stage1_16[16]}
   );
   gpc1_1 gpc268 (
      {stage0_16[18]},
      {stage1_16[17]}
   );
   gpc1_1 gpc269 (
      {stage0_16[19]},
      {stage1_16[18]}
   );
   gpc1_1 gpc270 (
      {stage0_16[20]},
      {stage1_16[19]}
   );
   gpc1_1 gpc271 (
      {stage0_16[21]},
      {stage1_16[20]}
   );
   gpc1_1 gpc272 (
      {stage0_16[22]},
      {stage1_16[21]}
   );
   gpc1_1 gpc273 (
      {stage0_16[23]},
      {stage1_16[22]}
   );
   gpc1_1 gpc274 (
      {stage0_16[24]},
      {stage1_16[23]}
   );
   gpc1_1 gpc275 (
      {stage0_16[25]},
      {stage1_16[24]}
   );
   gpc1_1 gpc276 (
      {stage0_16[26]},
      {stage1_16[25]}
   );
   gpc1_1 gpc277 (
      {stage0_16[27]},
      {stage1_16[26]}
   );
   gpc1_1 gpc278 (
      {stage0_16[28]},
      {stage1_16[27]}
   );
   gpc1_1 gpc279 (
      {stage0_16[29]},
      {stage1_16[28]}
   );
   gpc1_1 gpc280 (
      {stage0_16[30]},
      {stage1_16[29]}
   );
   gpc1_1 gpc281 (
      {stage0_16[31]},
      {stage1_16[30]}
   );
   gpc1_1 gpc282 (
      {stage0_17[19]},
      {stage1_17[9]}
   );
   gpc1_1 gpc283 (
      {stage0_17[20]},
      {stage1_17[10]}
   );
   gpc1_1 gpc284 (
      {stage0_17[21]},
      {stage1_17[11]}
   );
   gpc1_1 gpc285 (
      {stage0_17[22]},
      {stage1_17[12]}
   );
   gpc1_1 gpc286 (
      {stage0_17[23]},
      {stage1_17[13]}
   );
   gpc1_1 gpc287 (
      {stage0_17[24]},
      {stage1_17[14]}
   );
   gpc1_1 gpc288 (
      {stage0_17[25]},
      {stage1_17[15]}
   );
   gpc1_1 gpc289 (
      {stage0_17[26]},
      {stage1_17[16]}
   );
   gpc1_1 gpc290 (
      {stage0_17[27]},
      {stage1_17[17]}
   );
   gpc1_1 gpc291 (
      {stage0_17[28]},
      {stage1_17[18]}
   );
   gpc1_1 gpc292 (
      {stage0_17[29]},
      {stage1_17[19]}
   );
   gpc1_1 gpc293 (
      {stage0_17[30]},
      {stage1_17[20]}
   );
   gpc1_1 gpc294 (
      {stage0_17[31]},
      {stage1_17[21]}
   );
   gpc1_1 gpc295 (
      {stage0_18[29]},
      {stage1_18[8]}
   );
   gpc1_1 gpc296 (
      {stage0_18[30]},
      {stage1_18[9]}
   );
   gpc1_1 gpc297 (
      {stage0_18[31]},
      {stage1_18[10]}
   );
   gpc1_1 gpc298 (
      {stage0_19[23]},
      {stage1_19[10]}
   );
   gpc1_1 gpc299 (
      {stage0_19[24]},
      {stage1_19[11]}
   );
   gpc1_1 gpc300 (
      {stage0_19[25]},
      {stage1_19[12]}
   );
   gpc1_1 gpc301 (
      {stage0_19[26]},
      {stage1_19[13]}
   );
   gpc1_1 gpc302 (
      {stage0_19[27]},
      {stage1_19[14]}
   );
   gpc1_1 gpc303 (
      {stage0_19[28]},
      {stage1_19[15]}
   );
   gpc1_1 gpc304 (
      {stage0_19[29]},
      {stage1_19[16]}
   );
   gpc1_1 gpc305 (
      {stage0_19[30]},
      {stage1_19[17]}
   );
   gpc1_1 gpc306 (
      {stage0_19[31]},
      {stage1_19[18]}
   );
   gpc1_1 gpc307 (
      {stage0_21[26]},
      {stage1_21[12]}
   );
   gpc1_1 gpc308 (
      {stage0_21[27]},
      {stage1_21[13]}
   );
   gpc1_1 gpc309 (
      {stage0_21[28]},
      {stage1_21[14]}
   );
   gpc1_1 gpc310 (
      {stage0_21[29]},
      {stage1_21[15]}
   );
   gpc1_1 gpc311 (
      {stage0_21[30]},
      {stage1_21[16]}
   );
   gpc1_1 gpc312 (
      {stage0_21[31]},
      {stage1_21[17]}
   );
   gpc1_1 gpc313 (
      {stage0_22[31]},
      {stage1_22[13]}
   );
   gpc1_1 gpc314 (
      {stage0_23[25]},
      {stage1_23[11]}
   );
   gpc1_1 gpc315 (
      {stage0_23[26]},
      {stage1_23[12]}
   );
   gpc1_1 gpc316 (
      {stage0_23[27]},
      {stage1_23[13]}
   );
   gpc1_1 gpc317 (
      {stage0_23[28]},
      {stage1_23[14]}
   );
   gpc1_1 gpc318 (
      {stage0_23[29]},
      {stage1_23[15]}
   );
   gpc1_1 gpc319 (
      {stage0_23[30]},
      {stage1_23[16]}
   );
   gpc1_1 gpc320 (
      {stage0_23[31]},
      {stage1_23[17]}
   );
   gpc1_1 gpc321 (
      {stage0_25[27]},
      {stage1_25[13]}
   );
   gpc1_1 gpc322 (
      {stage0_25[28]},
      {stage1_25[14]}
   );
   gpc1_1 gpc323 (
      {stage0_25[29]},
      {stage1_25[15]}
   );
   gpc1_1 gpc324 (
      {stage0_25[30]},
      {stage1_25[16]}
   );
   gpc1_1 gpc325 (
      {stage0_25[31]},
      {stage1_25[17]}
   );
   gpc1_1 gpc326 (
      {stage0_26[27]},
      {stage1_26[12]}
   );
   gpc1_1 gpc327 (
      {stage0_26[28]},
      {stage1_26[13]}
   );
   gpc1_1 gpc328 (
      {stage0_26[29]},
      {stage1_26[14]}
   );
   gpc1_1 gpc329 (
      {stage0_26[30]},
      {stage1_26[15]}
   );
   gpc1_1 gpc330 (
      {stage0_26[31]},
      {stage1_26[16]}
   );
   gpc1_1 gpc331 (
      {stage0_27[31]},
      {stage1_27[10]}
   );
   gpc1_1 gpc332 (
      {stage0_28[29]},
      {stage1_28[13]}
   );
   gpc1_1 gpc333 (
      {stage0_28[30]},
      {stage1_28[14]}
   );
   gpc1_1 gpc334 (
      {stage0_28[31]},
      {stage1_28[15]}
   );
   gpc1_1 gpc335 (
      {stage0_29[28]},
      {stage1_29[14]}
   );
   gpc1_1 gpc336 (
      {stage0_29[29]},
      {stage1_29[15]}
   );
   gpc1_1 gpc337 (
      {stage0_29[30]},
      {stage1_29[16]}
   );
   gpc1_1 gpc338 (
      {stage0_29[31]},
      {stage1_29[17]}
   );
   gpc1_1 gpc339 (
      {stage0_31[25]},
      {stage1_31[10]}
   );
   gpc1_1 gpc340 (
      {stage0_31[26]},
      {stage1_31[11]}
   );
   gpc1_1 gpc341 (
      {stage0_31[27]},
      {stage1_31[12]}
   );
   gpc1_1 gpc342 (
      {stage0_31[28]},
      {stage1_31[13]}
   );
   gpc1_1 gpc343 (
      {stage0_31[29]},
      {stage1_31[14]}
   );
   gpc1_1 gpc344 (
      {stage0_31[30]},
      {stage1_31[15]}
   );
   gpc1_1 gpc345 (
      {stage0_31[31]},
      {stage1_31[16]}
   );
   gpc1_1 gpc346 (
      {stage0_32[18]},
      {stage1_32[11]}
   );
   gpc1_1 gpc347 (
      {stage0_32[19]},
      {stage1_32[12]}
   );
   gpc1_1 gpc348 (
      {stage0_32[20]},
      {stage1_32[13]}
   );
   gpc1_1 gpc349 (
      {stage0_32[21]},
      {stage1_32[14]}
   );
   gpc1_1 gpc350 (
      {stage0_32[22]},
      {stage1_32[15]}
   );
   gpc1_1 gpc351 (
      {stage0_32[23]},
      {stage1_32[16]}
   );
   gpc1_1 gpc352 (
      {stage0_32[24]},
      {stage1_32[17]}
   );
   gpc1_1 gpc353 (
      {stage0_32[25]},
      {stage1_32[18]}
   );
   gpc1_1 gpc354 (
      {stage0_32[26]},
      {stage1_32[19]}
   );
   gpc1_1 gpc355 (
      {stage0_32[27]},
      {stage1_32[20]}
   );
   gpc1_1 gpc356 (
      {stage0_32[28]},
      {stage1_32[21]}
   );
   gpc1_1 gpc357 (
      {stage0_32[29]},
      {stage1_32[22]}
   );
   gpc1_1 gpc358 (
      {stage0_32[30]},
      {stage1_32[23]}
   );
   gpc1_1 gpc359 (
      {stage0_32[31]},
      {stage1_32[24]}
   );
   gpc1_1 gpc360 (
      {stage0_33[24]},
      {stage1_33[11]}
   );
   gpc1_1 gpc361 (
      {stage0_33[25]},
      {stage1_33[12]}
   );
   gpc1_1 gpc362 (
      {stage0_33[26]},
      {stage1_33[13]}
   );
   gpc1_1 gpc363 (
      {stage0_33[27]},
      {stage1_33[14]}
   );
   gpc1_1 gpc364 (
      {stage0_33[28]},
      {stage1_33[15]}
   );
   gpc1_1 gpc365 (
      {stage0_33[29]},
      {stage1_33[16]}
   );
   gpc1_1 gpc366 (
      {stage0_33[30]},
      {stage1_33[17]}
   );
   gpc1_1 gpc367 (
      {stage0_33[31]},
      {stage1_33[18]}
   );
   gpc1_1 gpc368 (
      {stage0_34[20]},
      {stage1_34[9]}
   );
   gpc1_1 gpc369 (
      {stage0_34[21]},
      {stage1_34[10]}
   );
   gpc1_1 gpc370 (
      {stage0_34[22]},
      {stage1_34[11]}
   );
   gpc1_1 gpc371 (
      {stage0_34[23]},
      {stage1_34[12]}
   );
   gpc1_1 gpc372 (
      {stage0_34[24]},
      {stage1_34[13]}
   );
   gpc1_1 gpc373 (
      {stage0_34[25]},
      {stage1_34[14]}
   );
   gpc1_1 gpc374 (
      {stage0_34[26]},
      {stage1_34[15]}
   );
   gpc1_1 gpc375 (
      {stage0_34[27]},
      {stage1_34[16]}
   );
   gpc1_1 gpc376 (
      {stage0_34[28]},
      {stage1_34[17]}
   );
   gpc1_1 gpc377 (
      {stage0_34[29]},
      {stage1_34[18]}
   );
   gpc1_1 gpc378 (
      {stage0_34[30]},
      {stage1_34[19]}
   );
   gpc1_1 gpc379 (
      {stage0_34[31]},
      {stage1_34[20]}
   );
   gpc1_1 gpc380 (
      {stage0_35[27]},
      {stage1_35[8]}
   );
   gpc1_1 gpc381 (
      {stage0_35[28]},
      {stage1_35[9]}
   );
   gpc1_1 gpc382 (
      {stage0_35[29]},
      {stage1_35[10]}
   );
   gpc1_1 gpc383 (
      {stage0_35[30]},
      {stage1_35[11]}
   );
   gpc1_1 gpc384 (
      {stage0_35[31]},
      {stage1_35[12]}
   );
   gpc1_1 gpc385 (
      {stage0_36[30]},
      {stage1_36[11]}
   );
   gpc1_1 gpc386 (
      {stage0_36[31]},
      {stage1_36[12]}
   );
   gpc1_1 gpc387 (
      {stage0_38[25]},
      {stage1_38[11]}
   );
   gpc1_1 gpc388 (
      {stage0_38[26]},
      {stage1_38[12]}
   );
   gpc1_1 gpc389 (
      {stage0_38[27]},
      {stage1_38[13]}
   );
   gpc1_1 gpc390 (
      {stage0_38[28]},
      {stage1_38[14]}
   );
   gpc1_1 gpc391 (
      {stage0_38[29]},
      {stage1_38[15]}
   );
   gpc1_1 gpc392 (
      {stage0_38[30]},
      {stage1_38[16]}
   );
   gpc1_1 gpc393 (
      {stage0_38[31]},
      {stage1_38[17]}
   );
   gpc1_1 gpc394 (
      {stage0_39[27]},
      {stage1_39[10]}
   );
   gpc1_1 gpc395 (
      {stage0_39[28]},
      {stage1_39[11]}
   );
   gpc1_1 gpc396 (
      {stage0_39[29]},
      {stage1_39[12]}
   );
   gpc1_1 gpc397 (
      {stage0_39[30]},
      {stage1_39[13]}
   );
   gpc1_1 gpc398 (
      {stage0_39[31]},
      {stage1_39[14]}
   );
   gpc1_1 gpc399 (
      {stage0_40[30]},
      {stage1_40[14]}
   );
   gpc1_1 gpc400 (
      {stage0_40[31]},
      {stage1_40[15]}
   );
   gpc1_1 gpc401 (
      {stage0_41[24]},
      {stage1_41[12]}
   );
   gpc1_1 gpc402 (
      {stage0_41[25]},
      {stage1_41[13]}
   );
   gpc1_1 gpc403 (
      {stage0_41[26]},
      {stage1_41[14]}
   );
   gpc1_1 gpc404 (
      {stage0_41[27]},
      {stage1_41[15]}
   );
   gpc1_1 gpc405 (
      {stage0_41[28]},
      {stage1_41[16]}
   );
   gpc1_1 gpc406 (
      {stage0_41[29]},
      {stage1_41[17]}
   );
   gpc1_1 gpc407 (
      {stage0_41[30]},
      {stage1_41[18]}
   );
   gpc1_1 gpc408 (
      {stage0_41[31]},
      {stage1_41[19]}
   );
   gpc1_1 gpc409 (
      {stage0_42[29]},
      {stage1_42[10]}
   );
   gpc1_1 gpc410 (
      {stage0_42[30]},
      {stage1_42[11]}
   );
   gpc1_1 gpc411 (
      {stage0_42[31]},
      {stage1_42[12]}
   );
   gpc1_1 gpc412 (
      {stage0_43[29]},
      {stage1_43[11]}
   );
   gpc1_1 gpc413 (
      {stage0_43[30]},
      {stage1_43[12]}
   );
   gpc1_1 gpc414 (
      {stage0_43[31]},
      {stage1_43[13]}
   );
   gpc1_1 gpc415 (
      {stage0_45[18]},
      {stage1_45[11]}
   );
   gpc1_1 gpc416 (
      {stage0_45[19]},
      {stage1_45[12]}
   );
   gpc1_1 gpc417 (
      {stage0_45[20]},
      {stage1_45[13]}
   );
   gpc1_1 gpc418 (
      {stage0_45[21]},
      {stage1_45[14]}
   );
   gpc1_1 gpc419 (
      {stage0_45[22]},
      {stage1_45[15]}
   );
   gpc1_1 gpc420 (
      {stage0_45[23]},
      {stage1_45[16]}
   );
   gpc1_1 gpc421 (
      {stage0_45[24]},
      {stage1_45[17]}
   );
   gpc1_1 gpc422 (
      {stage0_45[25]},
      {stage1_45[18]}
   );
   gpc1_1 gpc423 (
      {stage0_45[26]},
      {stage1_45[19]}
   );
   gpc1_1 gpc424 (
      {stage0_45[27]},
      {stage1_45[20]}
   );
   gpc1_1 gpc425 (
      {stage0_45[28]},
      {stage1_45[21]}
   );
   gpc1_1 gpc426 (
      {stage0_45[29]},
      {stage1_45[22]}
   );
   gpc1_1 gpc427 (
      {stage0_45[30]},
      {stage1_45[23]}
   );
   gpc1_1 gpc428 (
      {stage0_45[31]},
      {stage1_45[24]}
   );
   gpc1_1 gpc429 (
      {stage0_46[29]},
      {stage1_46[9]}
   );
   gpc1_1 gpc430 (
      {stage0_46[30]},
      {stage1_46[10]}
   );
   gpc1_1 gpc431 (
      {stage0_46[31]},
      {stage1_46[11]}
   );
   gpc1_1 gpc432 (
      {stage0_47[25]},
      {stage1_47[11]}
   );
   gpc1_1 gpc433 (
      {stage0_47[26]},
      {stage1_47[12]}
   );
   gpc1_1 gpc434 (
      {stage0_47[27]},
      {stage1_47[13]}
   );
   gpc1_1 gpc435 (
      {stage0_47[28]},
      {stage1_47[14]}
   );
   gpc1_1 gpc436 (
      {stage0_47[29]},
      {stage1_47[15]}
   );
   gpc1_1 gpc437 (
      {stage0_47[30]},
      {stage1_47[16]}
   );
   gpc1_1 gpc438 (
      {stage0_47[31]},
      {stage1_47[17]}
   );
   gpc1_1 gpc439 (
      {stage0_48[24]},
      {stage1_48[12]}
   );
   gpc1_1 gpc440 (
      {stage0_48[25]},
      {stage1_48[13]}
   );
   gpc1_1 gpc441 (
      {stage0_48[26]},
      {stage1_48[14]}
   );
   gpc1_1 gpc442 (
      {stage0_48[27]},
      {stage1_48[15]}
   );
   gpc1_1 gpc443 (
      {stage0_48[28]},
      {stage1_48[16]}
   );
   gpc1_1 gpc444 (
      {stage0_48[29]},
      {stage1_48[17]}
   );
   gpc1_1 gpc445 (
      {stage0_48[30]},
      {stage1_48[18]}
   );
   gpc1_1 gpc446 (
      {stage0_48[31]},
      {stage1_48[19]}
   );
   gpc1_1 gpc447 (
      {stage0_49[21]},
      {stage1_49[9]}
   );
   gpc1_1 gpc448 (
      {stage0_49[22]},
      {stage1_49[10]}
   );
   gpc1_1 gpc449 (
      {stage0_49[23]},
      {stage1_49[11]}
   );
   gpc1_1 gpc450 (
      {stage0_49[24]},
      {stage1_49[12]}
   );
   gpc1_1 gpc451 (
      {stage0_49[25]},
      {stage1_49[13]}
   );
   gpc1_1 gpc452 (
      {stage0_49[26]},
      {stage1_49[14]}
   );
   gpc1_1 gpc453 (
      {stage0_49[27]},
      {stage1_49[15]}
   );
   gpc1_1 gpc454 (
      {stage0_49[28]},
      {stage1_49[16]}
   );
   gpc1_1 gpc455 (
      {stage0_49[29]},
      {stage1_49[17]}
   );
   gpc1_1 gpc456 (
      {stage0_49[30]},
      {stage1_49[18]}
   );
   gpc1_1 gpc457 (
      {stage0_49[31]},
      {stage1_49[19]}
   );
   gpc1_1 gpc458 (
      {stage0_50[30]},
      {stage1_50[10]}
   );
   gpc1_1 gpc459 (
      {stage0_50[31]},
      {stage1_50[11]}
   );
   gpc1_1 gpc460 (
      {stage0_51[23]},
      {stage1_51[12]}
   );
   gpc1_1 gpc461 (
      {stage0_51[24]},
      {stage1_51[13]}
   );
   gpc1_1 gpc462 (
      {stage0_51[25]},
      {stage1_51[14]}
   );
   gpc1_1 gpc463 (
      {stage0_51[26]},
      {stage1_51[15]}
   );
   gpc1_1 gpc464 (
      {stage0_51[27]},
      {stage1_51[16]}
   );
   gpc1_1 gpc465 (
      {stage0_51[28]},
      {stage1_51[17]}
   );
   gpc1_1 gpc466 (
      {stage0_51[29]},
      {stage1_51[18]}
   );
   gpc1_1 gpc467 (
      {stage0_51[30]},
      {stage1_51[19]}
   );
   gpc1_1 gpc468 (
      {stage0_51[31]},
      {stage1_51[20]}
   );
   gpc1_1 gpc469 (
      {stage0_53[18]},
      {stage1_53[9]}
   );
   gpc1_1 gpc470 (
      {stage0_53[19]},
      {stage1_53[10]}
   );
   gpc1_1 gpc471 (
      {stage0_53[20]},
      {stage1_53[11]}
   );
   gpc1_1 gpc472 (
      {stage0_53[21]},
      {stage1_53[12]}
   );
   gpc1_1 gpc473 (
      {stage0_53[22]},
      {stage1_53[13]}
   );
   gpc1_1 gpc474 (
      {stage0_53[23]},
      {stage1_53[14]}
   );
   gpc1_1 gpc475 (
      {stage0_53[24]},
      {stage1_53[15]}
   );
   gpc1_1 gpc476 (
      {stage0_53[25]},
      {stage1_53[16]}
   );
   gpc1_1 gpc477 (
      {stage0_53[26]},
      {stage1_53[17]}
   );
   gpc1_1 gpc478 (
      {stage0_53[27]},
      {stage1_53[18]}
   );
   gpc1_1 gpc479 (
      {stage0_53[28]},
      {stage1_53[19]}
   );
   gpc1_1 gpc480 (
      {stage0_53[29]},
      {stage1_53[20]}
   );
   gpc1_1 gpc481 (
      {stage0_53[30]},
      {stage1_53[21]}
   );
   gpc1_1 gpc482 (
      {stage0_53[31]},
      {stage1_53[22]}
   );
   gpc1_1 gpc483 (
      {stage0_55[13]},
      {stage1_55[11]}
   );
   gpc1_1 gpc484 (
      {stage0_55[14]},
      {stage1_55[12]}
   );
   gpc1_1 gpc485 (
      {stage0_55[15]},
      {stage1_55[13]}
   );
   gpc1_1 gpc486 (
      {stage0_55[16]},
      {stage1_55[14]}
   );
   gpc1_1 gpc487 (
      {stage0_55[17]},
      {stage1_55[15]}
   );
   gpc1_1 gpc488 (
      {stage0_55[18]},
      {stage1_55[16]}
   );
   gpc1_1 gpc489 (
      {stage0_55[19]},
      {stage1_55[17]}
   );
   gpc1_1 gpc490 (
      {stage0_55[20]},
      {stage1_55[18]}
   );
   gpc1_1 gpc491 (
      {stage0_55[21]},
      {stage1_55[19]}
   );
   gpc1_1 gpc492 (
      {stage0_55[22]},
      {stage1_55[20]}
   );
   gpc1_1 gpc493 (
      {stage0_55[23]},
      {stage1_55[21]}
   );
   gpc1_1 gpc494 (
      {stage0_55[24]},
      {stage1_55[22]}
   );
   gpc1_1 gpc495 (
      {stage0_55[25]},
      {stage1_55[23]}
   );
   gpc1_1 gpc496 (
      {stage0_55[26]},
      {stage1_55[24]}
   );
   gpc1_1 gpc497 (
      {stage0_55[27]},
      {stage1_55[25]}
   );
   gpc1_1 gpc498 (
      {stage0_55[28]},
      {stage1_55[26]}
   );
   gpc1_1 gpc499 (
      {stage0_55[29]},
      {stage1_55[27]}
   );
   gpc1_1 gpc500 (
      {stage0_55[30]},
      {stage1_55[28]}
   );
   gpc1_1 gpc501 (
      {stage0_55[31]},
      {stage1_55[29]}
   );
   gpc1_1 gpc502 (
      {stage0_56[28]},
      {stage1_56[11]}
   );
   gpc1_1 gpc503 (
      {stage0_56[29]},
      {stage1_56[12]}
   );
   gpc1_1 gpc504 (
      {stage0_56[30]},
      {stage1_56[13]}
   );
   gpc1_1 gpc505 (
      {stage0_56[31]},
      {stage1_56[14]}
   );
   gpc1_1 gpc506 (
      {stage0_57[25]},
      {stage1_57[10]}
   );
   gpc1_1 gpc507 (
      {stage0_57[26]},
      {stage1_57[11]}
   );
   gpc1_1 gpc508 (
      {stage0_57[27]},
      {stage1_57[12]}
   );
   gpc1_1 gpc509 (
      {stage0_57[28]},
      {stage1_57[13]}
   );
   gpc1_1 gpc510 (
      {stage0_57[29]},
      {stage1_57[14]}
   );
   gpc1_1 gpc511 (
      {stage0_57[30]},
      {stage1_57[15]}
   );
   gpc1_1 gpc512 (
      {stage0_57[31]},
      {stage1_57[16]}
   );
   gpc1_1 gpc513 (
      {stage0_58[27]},
      {stage1_58[9]}
   );
   gpc1_1 gpc514 (
      {stage0_58[28]},
      {stage1_58[10]}
   );
   gpc1_1 gpc515 (
      {stage0_58[29]},
      {stage1_58[11]}
   );
   gpc1_1 gpc516 (
      {stage0_58[30]},
      {stage1_58[12]}
   );
   gpc1_1 gpc517 (
      {stage0_58[31]},
      {stage1_58[13]}
   );
   gpc1_1 gpc518 (
      {stage0_59[18]},
      {stage1_59[10]}
   );
   gpc1_1 gpc519 (
      {stage0_59[19]},
      {stage1_59[11]}
   );
   gpc1_1 gpc520 (
      {stage0_59[20]},
      {stage1_59[12]}
   );
   gpc1_1 gpc521 (
      {stage0_59[21]},
      {stage1_59[13]}
   );
   gpc1_1 gpc522 (
      {stage0_59[22]},
      {stage1_59[14]}
   );
   gpc1_1 gpc523 (
      {stage0_59[23]},
      {stage1_59[15]}
   );
   gpc1_1 gpc524 (
      {stage0_59[24]},
      {stage1_59[16]}
   );
   gpc1_1 gpc525 (
      {stage0_59[25]},
      {stage1_59[17]}
   );
   gpc1_1 gpc526 (
      {stage0_59[26]},
      {stage1_59[18]}
   );
   gpc1_1 gpc527 (
      {stage0_59[27]},
      {stage1_59[19]}
   );
   gpc1_1 gpc528 (
      {stage0_59[28]},
      {stage1_59[20]}
   );
   gpc1_1 gpc529 (
      {stage0_59[29]},
      {stage1_59[21]}
   );
   gpc1_1 gpc530 (
      {stage0_59[30]},
      {stage1_59[22]}
   );
   gpc1_1 gpc531 (
      {stage0_59[31]},
      {stage1_59[23]}
   );
   gpc1_1 gpc532 (
      {stage0_60[30]},
      {stage1_60[11]}
   );
   gpc1_1 gpc533 (
      {stage0_60[31]},
      {stage1_60[12]}
   );
   gpc1_1 gpc534 (
      {stage0_62[26]},
      {stage1_62[11]}
   );
   gpc1_1 gpc535 (
      {stage0_62[27]},
      {stage1_62[12]}
   );
   gpc1_1 gpc536 (
      {stage0_62[28]},
      {stage1_62[13]}
   );
   gpc1_1 gpc537 (
      {stage0_62[29]},
      {stage1_62[14]}
   );
   gpc1_1 gpc538 (
      {stage0_62[30]},
      {stage1_62[15]}
   );
   gpc1_1 gpc539 (
      {stage0_62[31]},
      {stage1_62[16]}
   );
   gpc1_1 gpc540 (
      {stage0_63[31]},
      {stage1_63[10]}
   );
   gpc606_5 gpc541 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0]}
   );
   gpc606_5 gpc542 (
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[1],stage2_4[1],stage2_3[1],stage2_2[1]}
   );
   gpc615_5 gpc543 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[2],stage2_4[2],stage2_3[2],stage2_2[2]}
   );
   gpc615_5 gpc544 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[3],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc545 (
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_3[8]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[4],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc546 (
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[5],stage2_4[5],stage2_3[5]}
   );
   gpc606_5 gpc547 (
      {stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29], 1'b0},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[5],stage2_5[6],stage2_4[6]}
   );
   gpc606_5 gpc548 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[2],stage2_6[6],stage2_5[7]}
   );
   gpc615_5 gpc549 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[3],stage2_6[7]}
   );
   gpc615_5 gpc550 (
      {stage1_6[11], stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[4],stage2_6[8]}
   );
   gpc615_5 gpc551 (
      {stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20]},
      {stage1_7[8]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[5],stage2_6[9]}
   );
   gpc606_5 gpc552 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc553 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[5]}
   );
   gpc606_5 gpc554 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[2],stage2_11[2],stage2_10[5]}
   );
   gpc606_5 gpc555 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[3],stage2_11[3],stage2_10[6]}
   );
   gpc606_5 gpc556 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[4],stage2_11[4],stage2_10[7]}
   );
   gpc615_5 gpc557 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[18]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[3],stage2_13[5],stage2_12[5],stage2_11[5]}
   );
   gpc606_5 gpc558 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[1],stage2_14[4],stage2_13[6]}
   );
   gpc1163_5 gpc559 (
      {stage1_14[0], stage1_14[1], stage1_14[2]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[2],stage2_14[5]}
   );
   gpc615_5 gpc560 (
      {stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage1_15[12]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[3],stage2_14[6]}
   );
   gpc615_5 gpc561 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {1'b0},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[4],stage2_14[7]}
   );
   gpc606_5 gpc562 (
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[3],stage2_17[4],stage2_16[4]}
   );
   gpc606_5 gpc563 (
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], 1'b0},
      {stage2_20[1],stage2_19[1],stage2_18[4],stage2_17[5],stage2_16[5]}
   );
   gpc606_5 gpc564 (
      {stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[5],stage2_17[6]}
   );
   gpc606_5 gpc565 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[6],stage2_17[7]}
   );
   gpc606_5 gpc566 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[7],stage2_17[8]}
   );
   gpc1163_5 gpc567 (
      {stage1_20[0], stage1_20[1], stage1_20[2]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_22[0]},
      {stage1_23[0]},
      {stage2_24[0],stage2_23[0],stage2_22[0],stage2_21[3],stage2_20[5]}
   );
   gpc1163_5 gpc568 (
      {stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage1_22[1]},
      {stage1_23[1]},
      {stage2_24[1],stage2_23[1],stage2_22[1],stage2_21[4],stage2_20[6]}
   );
   gpc606_5 gpc569 (
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5], stage1_22[6], stage1_22[7]},
      {stage2_24[2],stage2_23[2],stage2_22[2],stage2_21[5],stage2_20[7]}
   );
   gpc606_5 gpc570 (
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5], stage1_23[6], stage1_23[7]},
      {stage2_25[0],stage2_24[3],stage2_23[3],stage2_22[3],stage2_21[6]}
   );
   gpc615_5 gpc571 (
      {stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11], stage1_23[12]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[0],stage2_25[1],stage2_24[4],stage2_23[4]}
   );
   gpc615_5 gpc572 (
      {stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage1_24[1]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[1],stage2_25[2],stage2_24[5],stage2_23[5]}
   );
   gpc615_5 gpc573 (
      {stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage1_25[12]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[2],stage2_26[2],stage2_25[3],stage2_24[6]}
   );
   gpc615_5 gpc574 (
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage1_25[13]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[3],stage2_26[3],stage2_25[4],stage2_24[7]}
   );
   gpc606_5 gpc575 (
      {stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], 1'b0, 1'b0},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[4],stage2_26[4],stage2_25[5]}
   );
   gpc615_5 gpc576 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16]},
      {stage1_27[6]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[1],stage2_28[3],stage2_27[5],stage2_26[5]}
   );
   gpc615_5 gpc577 (
      {stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], 1'b0},
      {stage1_28[6]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[1],stage2_29[2],stage2_28[4],stage2_27[6]}
   );
   gpc606_5 gpc578 (
      {stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[2],stage2_29[3],stage2_28[5]}
   );
   gpc606_5 gpc579 (
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[2],stage2_30[3],stage2_29[4]}
   );
   gpc606_5 gpc580 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[3],stage2_30[4],stage2_29[5]}
   );
   gpc615_5 gpc581 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10]},
      {stage1_31[12]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[2],stage2_32[3],stage2_31[4],stage2_30[5]}
   );
   gpc1406_5 gpc582 (
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3]},
      {stage1_35[0]},
      {stage2_36[0],stage2_35[0],stage2_34[1],stage2_33[3],stage2_32[4]}
   );
   gpc1406_5 gpc583 (
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage1_34[4], stage1_34[5], stage1_34[6], stage1_34[7]},
      {stage1_35[1]},
      {stage2_36[1],stage2_35[1],stage2_34[2],stage2_33[4],stage2_32[5]}
   );
   gpc606_5 gpc584 (
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11], stage1_34[12], stage1_34[13]},
      {stage2_36[2],stage2_35[2],stage2_34[3],stage2_33[5],stage2_32[6]}
   );
   gpc615_5 gpc585 (
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4]},
      {stage1_34[14]},
      {stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6], stage1_35[7]},
      {stage2_37[0],stage2_36[3],stage2_35[3],stage2_34[4],stage2_33[6]}
   );
   gpc615_5 gpc586 (
      {stage1_33[5], stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9]},
      {stage1_34[15]},
      {stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11], stage1_35[12], 1'b0},
      {stage2_37[1],stage2_36[4],stage2_35[4],stage2_34[5],stage2_33[7]}
   );
   gpc615_5 gpc587 (
      {stage1_34[16], stage1_34[17], stage1_34[18], stage1_34[19], stage1_34[20]},
      {1'b0},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[2],stage2_36[5],stage2_35[5],stage2_34[6]}
   );
   gpc606_5 gpc588 (
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[0],stage2_38[1],stage2_37[3],stage2_36[6]}
   );
   gpc615_5 gpc589 (
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4]},
      {stage1_38[6]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[2],stage2_37[4]}
   );
   gpc606_5 gpc590 (
      {stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[3]}
   );
   gpc615_5 gpc591 (
      {stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17]},
      {stage1_39[6]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[4]}
   );
   gpc606_5 gpc592 (
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[2],stage2_41[3],stage2_40[4],stage2_39[4]}
   );
   gpc606_5 gpc593 (
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], 1'b0, 1'b0},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[1],stage2_42[3],stage2_41[4],stage2_40[5]}
   );
   gpc117_4 gpc594 (
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11], stage1_41[12]},
      {stage1_42[6]},
      {stage1_43[0]},
      {stage2_44[1],stage2_43[2],stage2_42[4],stage2_41[5]}
   );
   gpc117_4 gpc595 (
      {stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19]},
      {stage1_42[7]},
      {stage1_43[1]},
      {stage2_44[2],stage2_43[3],stage2_42[5],stage2_41[6]}
   );
   gpc606_5 gpc596 (
      {stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5], stage1_43[6], stage1_43[7]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[0],stage2_44[3],stage2_43[4]}
   );
   gpc615_5 gpc597 (
      {stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11], stage1_43[12]},
      {stage1_44[0]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[1],stage2_44[4],stage2_43[5]}
   );
   gpc606_5 gpc598 (
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[2],stage2_46[2],stage2_45[2]}
   );
   gpc606_5 gpc599 (
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[1],stage2_47[3],stage2_46[3],stage2_45[3]}
   );
   gpc615_5 gpc600 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4]},
      {stage1_47[12]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[2],stage2_48[2],stage2_47[4],stage2_46[4]}
   );
   gpc615_5 gpc601 (
      {stage1_46[5], stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9]},
      {stage1_47[13]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[3],stage2_48[3],stage2_47[5],stage2_46[5]}
   );
   gpc606_5 gpc602 (
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[0],stage2_50[2],stage2_49[4],stage2_48[4]}
   );
   gpc606_5 gpc603 (
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[1],stage2_51[1],stage2_50[3],stage2_49[5]}
   );
   gpc615_5 gpc604 (
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10]},
      {stage1_50[6]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[2],stage2_51[2],stage2_50[4],stage2_49[6]}
   );
   gpc615_5 gpc605 (
      {stage1_49[11], stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15]},
      {stage1_50[7]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[3],stage2_51[3],stage2_50[5],stage2_49[7]}
   );
   gpc615_5 gpc606 (
      {stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11], 1'b0},
      {stage1_51[18]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[3],stage2_52[4],stage2_51[4],stage2_50[6]}
   );
   gpc1163_5 gpc607 (
      {stage1_51[19], stage1_51[20], 1'b0},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage1_53[0]},
      {stage1_54[0]},
      {stage2_55[0],stage2_54[1],stage2_53[4],stage2_52[5],stage2_51[5]}
   );
   gpc615_5 gpc608 (
      {stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage1_54[1]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[0],stage2_55[1],stage2_54[2],stage2_53[5]}
   );
   gpc615_5 gpc609 (
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10]},
      {stage1_54[2]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[1],stage2_55[2],stage2_54[3],stage2_53[6]}
   );
   gpc615_5 gpc610 (
      {stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15]},
      {stage1_54[3]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[2],stage2_55[3],stage2_54[4],stage2_53[7]}
   );
   gpc615_5 gpc611 (
      {stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20]},
      {stage1_54[4]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[3],stage2_55[4],stage2_54[5],stage2_53[8]}
   );
   gpc615_5 gpc612 (
      {stage1_54[5], stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9]},
      {stage1_55[24]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[4],stage2_56[4],stage2_55[5],stage2_54[6]}
   );
   gpc615_5 gpc613 (
      {stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage1_56[6]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[1],stage2_57[5],stage2_56[5],stage2_55[6]}
   );
   gpc615_5 gpc614 (
      {stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage1_57[6]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[1],stage2_58[2],stage2_57[6],stage2_56[6]}
   );
   gpc615_5 gpc615 (
      {stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage1_58[6]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[1],stage2_59[2],stage2_58[3],stage2_57[7]}
   );
   gpc615_5 gpc616 (
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16]},
      {stage1_58[7]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[2],stage2_59[3],stage2_58[4],stage2_57[8]}
   );
   gpc606_5 gpc617 (
      {stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11], stage1_58[12], stage1_58[13]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[2],stage2_60[3],stage2_59[4],stage2_58[5]}
   );
   gpc606_5 gpc618 (
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[1],stage2_61[3],stage2_60[4],stage2_59[5]}
   );
   gpc606_5 gpc619 (
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[1],stage2_62[2],stage2_61[4],stage2_60[5]}
   );
   gpc606_5 gpc620 (
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[1],stage2_63[2],stage2_62[3],stage2_61[5]}
   );
   gpc207_4 gpc621 (
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11], stage1_62[12]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[1],stage2_64[2],stage2_63[3],stage2_62[4]}
   );
   gpc606_5 gpc622 (
      {stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], 1'b0, 1'b0},
      {stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7]},
      {stage2_66[0],stage2_65[2],stage2_64[3],stage2_63[4],stage2_62[5]}
   );
   gpc1_1 gpc623 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc624 (
      {stage1_0[1]},
      {stage2_0[1]}
   );
   gpc1_1 gpc625 (
      {stage1_0[2]},
      {stage2_0[2]}
   );
   gpc1_1 gpc626 (
      {stage1_0[3]},
      {stage2_0[3]}
   );
   gpc1_1 gpc627 (
      {stage1_0[4]},
      {stage2_0[4]}
   );
   gpc1_1 gpc628 (
      {stage1_0[5]},
      {stage2_0[5]}
   );
   gpc1_1 gpc629 (
      {stage1_0[6]},
      {stage2_0[6]}
   );
   gpc1_1 gpc630 (
      {stage1_0[7]},
      {stage2_0[7]}
   );
   gpc1_1 gpc631 (
      {stage1_0[8]},
      {stage2_0[8]}
   );
   gpc1_1 gpc632 (
      {stage1_0[9]},
      {stage2_0[9]}
   );
   gpc1_1 gpc633 (
      {stage1_0[10]},
      {stage2_0[10]}
   );
   gpc1_1 gpc634 (
      {stage1_1[6]},
      {stage2_1[1]}
   );
   gpc1_1 gpc635 (
      {stage1_1[7]},
      {stage2_1[2]}
   );
   gpc1_1 gpc636 (
      {stage1_2[21]},
      {stage2_2[5]}
   );
   gpc1_1 gpc637 (
      {stage1_2[22]},
      {stage2_2[6]}
   );
   gpc1_1 gpc638 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc639 (
      {stage1_2[24]},
      {stage2_2[8]}
   );
   gpc1_1 gpc640 (
      {stage1_3[14]},
      {stage2_3[6]}
   );
   gpc1_1 gpc641 (
      {stage1_3[15]},
      {stage2_3[7]}
   );
   gpc1_1 gpc642 (
      {stage1_3[16]},
      {stage2_3[8]}
   );
   gpc1_1 gpc643 (
      {stage1_5[12]},
      {stage2_5[8]}
   );
   gpc1_1 gpc644 (
      {stage1_5[13]},
      {stage2_5[9]}
   );
   gpc1_1 gpc645 (
      {stage1_6[21]},
      {stage2_6[10]}
   );
   gpc1_1 gpc646 (
      {stage1_6[22]},
      {stage2_6[11]}
   );
   gpc1_1 gpc647 (
      {stage1_6[23]},
      {stage2_6[12]}
   );
   gpc1_1 gpc648 (
      {stage1_6[24]},
      {stage2_6[13]}
   );
   gpc1_1 gpc649 (
      {stage1_6[25]},
      {stage2_6[14]}
   );
   gpc1_1 gpc650 (
      {stage1_6[26]},
      {stage2_6[15]}
   );
   gpc1_1 gpc651 (
      {stage1_6[27]},
      {stage2_6[16]}
   );
   gpc1_1 gpc652 (
      {stage1_6[28]},
      {stage2_6[17]}
   );
   gpc1_1 gpc653 (
      {stage1_8[18]},
      {stage2_8[5]}
   );
   gpc1_1 gpc654 (
      {stage1_9[12]},
      {stage2_9[6]}
   );
   gpc1_1 gpc655 (
      {stage1_9[13]},
      {stage2_9[7]}
   );
   gpc1_1 gpc656 (
      {stage1_9[14]},
      {stage2_9[8]}
   );
   gpc1_1 gpc657 (
      {stage1_9[15]},
      {stage2_9[9]}
   );
   gpc1_1 gpc658 (
      {stage1_13[12]},
      {stage2_13[7]}
   );
   gpc1_1 gpc659 (
      {stage1_13[13]},
      {stage2_13[8]}
   );
   gpc1_1 gpc660 (
      {stage1_14[13]},
      {stage2_14[8]}
   );
   gpc1_1 gpc661 (
      {stage1_14[14]},
      {stage2_14[9]}
   );
   gpc1_1 gpc662 (
      {stage1_14[15]},
      {stage2_14[10]}
   );
   gpc1_1 gpc663 (
      {stage1_14[16]},
      {stage2_14[11]}
   );
   gpc1_1 gpc664 (
      {stage1_16[25]},
      {stage2_16[6]}
   );
   gpc1_1 gpc665 (
      {stage1_16[26]},
      {stage2_16[7]}
   );
   gpc1_1 gpc666 (
      {stage1_16[27]},
      {stage2_16[8]}
   );
   gpc1_1 gpc667 (
      {stage1_16[28]},
      {stage2_16[9]}
   );
   gpc1_1 gpc668 (
      {stage1_16[29]},
      {stage2_16[10]}
   );
   gpc1_1 gpc669 (
      {stage1_16[30]},
      {stage2_16[11]}
   );
   gpc1_1 gpc670 (
      {stage1_17[19]},
      {stage2_17[9]}
   );
   gpc1_1 gpc671 (
      {stage1_17[20]},
      {stage2_17[10]}
   );
   gpc1_1 gpc672 (
      {stage1_17[21]},
      {stage2_17[11]}
   );
   gpc1_1 gpc673 (
      {stage1_19[18]},
      {stage2_19[5]}
   );
   gpc1_1 gpc674 (
      {stage1_22[8]},
      {stage2_22[4]}
   );
   gpc1_1 gpc675 (
      {stage1_22[9]},
      {stage2_22[5]}
   );
   gpc1_1 gpc676 (
      {stage1_22[10]},
      {stage2_22[6]}
   );
   gpc1_1 gpc677 (
      {stage1_22[11]},
      {stage2_22[7]}
   );
   gpc1_1 gpc678 (
      {stage1_22[12]},
      {stage2_22[8]}
   );
   gpc1_1 gpc679 (
      {stage1_22[13]},
      {stage2_22[9]}
   );
   gpc1_1 gpc680 (
      {stage1_28[13]},
      {stage2_28[6]}
   );
   gpc1_1 gpc681 (
      {stage1_28[14]},
      {stage2_28[7]}
   );
   gpc1_1 gpc682 (
      {stage1_28[15]},
      {stage2_28[8]}
   );
   gpc1_1 gpc683 (
      {stage1_31[13]},
      {stage2_31[5]}
   );
   gpc1_1 gpc684 (
      {stage1_31[14]},
      {stage2_31[6]}
   );
   gpc1_1 gpc685 (
      {stage1_31[15]},
      {stage2_31[7]}
   );
   gpc1_1 gpc686 (
      {stage1_31[16]},
      {stage2_31[8]}
   );
   gpc1_1 gpc687 (
      {stage1_32[24]},
      {stage2_32[7]}
   );
   gpc1_1 gpc688 (
      {stage1_33[10]},
      {stage2_33[8]}
   );
   gpc1_1 gpc689 (
      {stage1_33[11]},
      {stage2_33[9]}
   );
   gpc1_1 gpc690 (
      {stage1_33[12]},
      {stage2_33[10]}
   );
   gpc1_1 gpc691 (
      {stage1_33[13]},
      {stage2_33[11]}
   );
   gpc1_1 gpc692 (
      {stage1_33[14]},
      {stage2_33[12]}
   );
   gpc1_1 gpc693 (
      {stage1_33[15]},
      {stage2_33[13]}
   );
   gpc1_1 gpc694 (
      {stage1_33[16]},
      {stage2_33[14]}
   );
   gpc1_1 gpc695 (
      {stage1_33[17]},
      {stage2_33[15]}
   );
   gpc1_1 gpc696 (
      {stage1_33[18]},
      {stage2_33[16]}
   );
   gpc1_1 gpc697 (
      {stage1_36[12]},
      {stage2_36[7]}
   );
   gpc1_1 gpc698 (
      {stage1_37[5]},
      {stage2_37[5]}
   );
   gpc1_1 gpc699 (
      {stage1_37[6]},
      {stage2_37[6]}
   );
   gpc1_1 gpc700 (
      {stage1_37[7]},
      {stage2_37[7]}
   );
   gpc1_1 gpc701 (
      {stage1_37[8]},
      {stage2_37[8]}
   );
   gpc1_1 gpc702 (
      {stage1_37[9]},
      {stage2_37[9]}
   );
   gpc1_1 gpc703 (
      {stage1_37[10]},
      {stage2_37[10]}
   );
   gpc1_1 gpc704 (
      {stage1_37[11]},
      {stage2_37[11]}
   );
   gpc1_1 gpc705 (
      {stage1_37[12]},
      {stage2_37[12]}
   );
   gpc1_1 gpc706 (
      {stage1_37[13]},
      {stage2_37[13]}
   );
   gpc1_1 gpc707 (
      {stage1_39[13]},
      {stage2_39[5]}
   );
   gpc1_1 gpc708 (
      {stage1_39[14]},
      {stage2_39[6]}
   );
   gpc1_1 gpc709 (
      {stage1_42[8]},
      {stage2_42[6]}
   );
   gpc1_1 gpc710 (
      {stage1_42[9]},
      {stage2_42[7]}
   );
   gpc1_1 gpc711 (
      {stage1_42[10]},
      {stage2_42[8]}
   );
   gpc1_1 gpc712 (
      {stage1_42[11]},
      {stage2_42[9]}
   );
   gpc1_1 gpc713 (
      {stage1_42[12]},
      {stage2_42[10]}
   );
   gpc1_1 gpc714 (
      {stage1_43[13]},
      {stage2_43[6]}
   );
   gpc1_1 gpc715 (
      {stage1_44[1]},
      {stage2_44[5]}
   );
   gpc1_1 gpc716 (
      {stage1_44[2]},
      {stage2_44[6]}
   );
   gpc1_1 gpc717 (
      {stage1_44[3]},
      {stage2_44[7]}
   );
   gpc1_1 gpc718 (
      {stage1_44[4]},
      {stage2_44[8]}
   );
   gpc1_1 gpc719 (
      {stage1_44[5]},
      {stage2_44[9]}
   );
   gpc1_1 gpc720 (
      {stage1_44[6]},
      {stage2_44[10]}
   );
   gpc1_1 gpc721 (
      {stage1_44[7]},
      {stage2_44[11]}
   );
   gpc1_1 gpc722 (
      {stage1_44[8]},
      {stage2_44[12]}
   );
   gpc1_1 gpc723 (
      {stage1_44[9]},
      {stage2_44[13]}
   );
   gpc1_1 gpc724 (
      {stage1_44[10]},
      {stage2_44[14]}
   );
   gpc1_1 gpc725 (
      {stage1_44[11]},
      {stage2_44[15]}
   );
   gpc1_1 gpc726 (
      {stage1_44[12]},
      {stage2_44[16]}
   );
   gpc1_1 gpc727 (
      {stage1_44[13]},
      {stage2_44[17]}
   );
   gpc1_1 gpc728 (
      {stage1_45[24]},
      {stage2_45[4]}
   );
   gpc1_1 gpc729 (
      {stage1_46[10]},
      {stage2_46[6]}
   );
   gpc1_1 gpc730 (
      {stage1_46[11]},
      {stage2_46[7]}
   );
   gpc1_1 gpc731 (
      {stage1_47[14]},
      {stage2_47[6]}
   );
   gpc1_1 gpc732 (
      {stage1_47[15]},
      {stage2_47[7]}
   );
   gpc1_1 gpc733 (
      {stage1_47[16]},
      {stage2_47[8]}
   );
   gpc1_1 gpc734 (
      {stage1_47[17]},
      {stage2_47[9]}
   );
   gpc1_1 gpc735 (
      {stage1_48[18]},
      {stage2_48[5]}
   );
   gpc1_1 gpc736 (
      {stage1_48[19]},
      {stage2_48[6]}
   );
   gpc1_1 gpc737 (
      {stage1_49[16]},
      {stage2_49[8]}
   );
   gpc1_1 gpc738 (
      {stage1_49[17]},
      {stage2_49[9]}
   );
   gpc1_1 gpc739 (
      {stage1_49[18]},
      {stage2_49[10]}
   );
   gpc1_1 gpc740 (
      {stage1_49[19]},
      {stage2_49[11]}
   );
   gpc1_1 gpc741 (
      {stage1_53[21]},
      {stage2_53[9]}
   );
   gpc1_1 gpc742 (
      {stage1_53[22]},
      {stage2_53[10]}
   );
   gpc1_1 gpc743 (
      {stage1_56[12]},
      {stage2_56[7]}
   );
   gpc1_1 gpc744 (
      {stage1_56[13]},
      {stage2_56[8]}
   );
   gpc1_1 gpc745 (
      {stage1_56[14]},
      {stage2_56[9]}
   );
   gpc1_1 gpc746 (
      {stage1_59[18]},
      {stage2_59[6]}
   );
   gpc1_1 gpc747 (
      {stage1_59[19]},
      {stage2_59[7]}
   );
   gpc1_1 gpc748 (
      {stage1_59[20]},
      {stage2_59[8]}
   );
   gpc1_1 gpc749 (
      {stage1_59[21]},
      {stage2_59[9]}
   );
   gpc1_1 gpc750 (
      {stage1_59[22]},
      {stage2_59[10]}
   );
   gpc1_1 gpc751 (
      {stage1_59[23]},
      {stage2_59[11]}
   );
   gpc1_1 gpc752 (
      {stage1_60[12]},
      {stage2_60[6]}
   );
   gpc1_1 gpc753 (
      {stage1_61[12]},
      {stage2_61[6]}
   );
   gpc1_1 gpc754 (
      {stage1_63[6]},
      {stage2_63[5]}
   );
   gpc1_1 gpc755 (
      {stage1_63[7]},
      {stage2_63[6]}
   );
   gpc1_1 gpc756 (
      {stage1_63[8]},
      {stage2_63[7]}
   );
   gpc1_1 gpc757 (
      {stage1_63[9]},
      {stage2_63[8]}
   );
   gpc1_1 gpc758 (
      {stage1_63[10]},
      {stage2_63[9]}
   );
   gpc1_1 gpc759 (
      {stage1_64[8]},
      {stage2_64[4]}
   );
   gpc1_1 gpc760 (
      {stage1_65[0]},
      {stage2_65[3]}
   );
   gpc1_1 gpc761 (
      {stage1_65[1]},
      {stage2_65[4]}
   );
   gpc1_1 gpc762 (
      {stage1_65[2]},
      {stage2_65[5]}
   );
   gpc1_1 gpc763 (
      {stage1_65[3]},
      {stage2_65[6]}
   );
   gpc1_1 gpc764 (
      {stage1_65[4]},
      {stage2_65[7]}
   );
   gpc135_4 gpc765 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc766 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1343_5 gpc767 (
      {stage2_3[0], stage2_3[1], stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc768 (
      {stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_4[4]},
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2],stage3_3[3]}
   );
   gpc2135_5 gpc769 (
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[2]}
   );
   gpc2135_5 gpc770 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10]},
      {stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_8[1]},
      {stage2_9[2], stage2_9[3]},
      {stage3_10[1],stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[3]}
   );
   gpc1406_5 gpc771 (
      {stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[4]},
      {stage3_10[2],stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[4]}
   );
   gpc615_5 gpc772 (
      {stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9]},
      {stage2_10[0]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[3],stage3_9[3]}
   );
   gpc606_5 gpc773 (
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[1],stage3_11[1],stage3_10[4]}
   );
   gpc7_3 gpc774 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[0],stage3_14[1],stage3_13[2]}
   );
   gpc606_5 gpc775 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[0],stage3_15[1],stage3_14[2]}
   );
   gpc606_5 gpc776 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[1],stage3_15[2],stage3_14[3]}
   );
   gpc615_5 gpc777 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4]},
      {1'b0},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[2],stage3_15[3]}
   );
   gpc606_5 gpc778 (
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[3],stage3_17[3]}
   );
   gpc7_3 gpc779 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[1],stage3_19[2],stage3_18[4]}
   );
   gpc606_5 gpc780 (
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[2]}
   );
   gpc117_4 gpc781 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6]},
      {stage2_22[6]},
      {stage2_23[0]},
      {stage3_24[1],stage3_23[1],stage3_22[1],stage3_21[2]}
   );
   gpc615_5 gpc782 (
      {stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage2_24[0]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[2],stage3_23[2]}
   );
   gpc606_5 gpc783 (
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[3]}
   );
   gpc615_5 gpc784 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4]},
      {stage2_28[0]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[0],stage3_28[1],stage3_27[2]}
   );
   gpc606_5 gpc785 (
      {stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[1],stage3_29[1],stage3_28[2]}
   );
   gpc615_5 gpc786 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4]},
      {stage2_32[0]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[2]}
   );
   gpc615_5 gpc787 (
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], 1'b0},
      {stage2_32[1]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[1],stage3_32[2],stage3_31[3]}
   );
   gpc606_5 gpc788 (
      {stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5], stage2_32[6], stage2_32[7]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[2],stage3_34[2],stage3_33[2],stage3_32[3]}
   );
   gpc615_5 gpc789 (
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16]},
      {stage2_34[6]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[3],stage3_34[3],stage3_33[3]}
   );
   gpc7_3 gpc790 (
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5], stage2_36[6]},
      {stage3_38[0],stage3_37[1],stage3_36[2]}
   );
   gpc7_3 gpc791 (
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5], stage2_37[6]},
      {stage3_39[0],stage3_38[1],stage3_37[2]}
   );
   gpc7_3 gpc792 (
      {stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11], stage2_37[12], stage2_37[13]},
      {stage3_39[1],stage3_38[2],stage3_37[3]}
   );
   gpc615_5 gpc793 (
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4]},
      {stage2_39[0]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[0],stage3_39[2],stage3_38[3]}
   );
   gpc606_5 gpc794 (
      {stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5], stage2_39[6]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[1],stage3_41[1],stage3_40[1],stage3_39[3]}
   );
   gpc615_5 gpc795 (
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[0],stage3_43[1],stage3_42[2]}
   );
   gpc615_5 gpc796 (
      {stage2_42[5], stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[1],stage3_43[2],stage3_42[3]}
   );
   gpc1325_5 gpc797 (
      {stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5], stage2_43[6]},
      {stage2_44[12], stage2_44[13]},
      {stage2_45[0], stage2_45[1], stage2_45[2]},
      {stage2_46[0]},
      {stage3_47[0],stage3_46[2],stage3_45[2],stage3_44[2],stage3_43[3]}
   );
   gpc135_4 gpc798 (
      {stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17], 1'b0},
      {stage2_45[3], stage2_45[4], 1'b0},
      {stage2_46[1]},
      {stage3_47[1],stage3_46[3],stage3_45[3],stage3_44[3]}
   );
   gpc615_5 gpc799 (
      {stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5], stage2_46[6]},
      {stage2_47[0]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[0],stage3_48[0],stage3_47[2],stage3_46[4]}
   );
   gpc615_5 gpc800 (
      {stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage2_48[6]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[1],stage3_49[1],stage3_48[1],stage3_47[3]}
   );
   gpc615_5 gpc801 (
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], 1'b0},
      {1'b0},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[1],stage3_50[2],stage3_49[2],stage3_48[2],stage3_47[4]}
   );
   gpc15_3 gpc802 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[2],stage3_50[3]}
   );
   gpc615_5 gpc803 (
      {stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[0],stage3_52[1],stage3_51[3]}
   );
   gpc1406_5 gpc804 (
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5], 1'b0},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3]},
      {stage2_55[0]},
      {stage3_56[0],stage3_55[1],stage3_54[1],stage3_53[1],stage3_52[2]}
   );
   gpc606_5 gpc805 (
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], 1'b0},
      {stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5], stage2_55[6]},
      {stage3_57[0],stage3_56[1],stage3_55[2],stage3_54[2],stage3_53[2]}
   );
   gpc135_4 gpc806 (
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4]},
      {stage2_57[0], stage2_57[1], stage2_57[2]},
      {stage2_58[0]},
      {stage3_59[0],stage3_58[0],stage3_57[1],stage3_56[2]}
   );
   gpc1163_5 gpc807 (
      {stage2_56[5], stage2_56[6], stage2_56[7]},
      {stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8]},
      {stage2_58[1]},
      {stage2_59[0]},
      {stage3_60[0],stage3_59[1],stage3_58[1],stage3_57[2],stage3_56[3]}
   );
   gpc1343_5 gpc808 (
      {stage2_58[2], stage2_58[3], stage2_58[4]},
      {stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4]},
      {stage2_60[0], stage2_60[1], stage2_60[2]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[0],stage3_60[1],stage3_59[2],stage3_58[2]}
   );
   gpc2135_5 gpc809 (
      {stage2_59[5], stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9]},
      {stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_61[1]},
      {stage2_62[0], stage2_62[1]},
      {stage3_63[0],stage3_62[1],stage3_61[1],stage3_60[2],stage3_59[3]}
   );
   gpc615_5 gpc810 (
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6]},
      {stage2_62[2]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[0],stage3_63[1],stage3_62[2],stage3_61[2]}
   );
   gpc615_5 gpc811 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], 1'b0},
      {stage2_64[0]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[0],stage3_65[1],stage3_64[1],stage3_63[2]}
   );
   gpc1_1 gpc812 (
      {stage2_2[7]},
      {stage3_2[2]}
   );
   gpc1_1 gpc813 (
      {stage2_2[8]},
      {stage3_2[3]}
   );
   gpc1_1 gpc814 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc815 (
      {stage2_4[5]},
      {stage3_4[3]}
   );
   gpc1_1 gpc816 (
      {stage2_4[6]},
      {stage3_4[4]}
   );
   gpc1_1 gpc817 (
      {stage2_5[9]},
      {stage3_5[2]}
   );
   gpc1_1 gpc818 (
      {stage2_6[17]},
      {stage3_6[5]}
   );
   gpc1_1 gpc819 (
      {stage2_10[7]},
      {stage3_10[5]}
   );
   gpc1_1 gpc820 (
      {stage2_13[7]},
      {stage3_13[3]}
   );
   gpc1_1 gpc821 (
      {stage2_13[8]},
      {stage3_13[4]}
   );
   gpc1_1 gpc822 (
      {stage2_18[7]},
      {stage3_18[5]}
   );
   gpc1_1 gpc823 (
      {stage2_20[6]},
      {stage3_20[3]}
   );
   gpc1_1 gpc824 (
      {stage2_20[7]},
      {stage3_20[4]}
   );
   gpc1_1 gpc825 (
      {stage2_22[7]},
      {stage3_22[2]}
   );
   gpc1_1 gpc826 (
      {stage2_22[8]},
      {stage3_22[3]}
   );
   gpc1_1 gpc827 (
      {stage2_22[9]},
      {stage3_22[4]}
   );
   gpc1_1 gpc828 (
      {stage2_24[7]},
      {stage3_24[4]}
   );
   gpc1_1 gpc829 (
      {stage2_27[5]},
      {stage3_27[3]}
   );
   gpc1_1 gpc830 (
      {stage2_27[6]},
      {stage3_27[4]}
   );
   gpc1_1 gpc831 (
      {stage2_28[7]},
      {stage3_28[3]}
   );
   gpc1_1 gpc832 (
      {stage2_28[8]},
      {stage3_28[4]}
   );
   gpc1_1 gpc833 (
      {stage2_36[7]},
      {stage3_36[3]}
   );
   gpc1_1 gpc834 (
      {stage2_41[6]},
      {stage3_41[2]}
   );
   gpc1_1 gpc835 (
      {stage2_42[10]},
      {stage3_42[4]}
   );
   gpc1_1 gpc836 (
      {stage2_46[7]},
      {stage3_46[5]}
   );
   gpc1_1 gpc837 (
      {stage2_50[5]},
      {stage3_50[4]}
   );
   gpc1_1 gpc838 (
      {stage2_50[6]},
      {stage3_50[5]}
   );
   gpc1_1 gpc839 (
      {stage2_54[4]},
      {stage3_54[3]}
   );
   gpc1_1 gpc840 (
      {stage2_54[5]},
      {stage3_54[4]}
   );
   gpc1_1 gpc841 (
      {stage2_54[6]},
      {stage3_54[5]}
   );
   gpc1_1 gpc842 (
      {stage2_56[8]},
      {stage3_56[4]}
   );
   gpc1_1 gpc843 (
      {stage2_56[9]},
      {stage3_56[5]}
   );
   gpc1_1 gpc844 (
      {stage2_58[5]},
      {stage3_58[3]}
   );
   gpc1_1 gpc845 (
      {stage2_59[10]},
      {stage3_59[4]}
   );
   gpc1_1 gpc846 (
      {stage2_59[11]},
      {stage3_59[5]}
   );
   gpc1_1 gpc847 (
      {stage2_60[6]},
      {stage3_60[3]}
   );
   gpc1_1 gpc848 (
      {stage2_62[3]},
      {stage3_62[3]}
   );
   gpc1_1 gpc849 (
      {stage2_62[4]},
      {stage3_62[4]}
   );
   gpc1_1 gpc850 (
      {stage2_62[5]},
      {stage3_62[5]}
   );
   gpc1_1 gpc851 (
      {stage2_64[1]},
      {stage3_64[2]}
   );
   gpc1_1 gpc852 (
      {stage2_64[2]},
      {stage3_64[3]}
   );
   gpc1_1 gpc853 (
      {stage2_64[3]},
      {stage3_64[4]}
   );
   gpc1_1 gpc854 (
      {stage2_64[4]},
      {stage3_64[5]}
   );
   gpc1_1 gpc855 (
      {stage2_65[6]},
      {stage3_65[2]}
   );
   gpc1_1 gpc856 (
      {stage2_65[7]},
      {stage3_65[3]}
   );
   gpc1_1 gpc857 (
      {stage2_66[0]},
      {stage3_66[1]}
   );
   gpc1343_5 gpc858 (
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc623_5 gpc859 (
      {stage3_4[3], stage3_4[4], 1'b0},
      {stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[1]}
   );
   gpc135_4 gpc860 (
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4]},
      {stage3_8[0], stage3_8[1], stage3_8[2]},
      {stage3_9[0]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc861 (
      {stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_11[0]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc1163_5 gpc862 (
      {stage3_12[1], 1'b0, 1'b0},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], 1'b0},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc1343_5 gpc863 (
      {stage3_14[1], stage3_14[2], stage3_14[3]},
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1]}
   );
   gpc1163_5 gpc864 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1]}
   );
   gpc1343_5 gpc865 (
      {stage3_19[1], stage3_19[2], 1'b0},
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[0], stage3_21[1], stage3_21[2]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[1],stage4_20[1],stage4_19[1]}
   );
   gpc2135_5 gpc866 (
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], 1'b0},
      {stage3_23[0], stage3_23[1], stage3_23[2]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1]},
      {stage4_26[0],stage4_25[0],stage4_24[0],stage4_23[1],stage4_22[1]}
   );
   gpc207_4 gpc867 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], 1'b0, 1'b0, 1'b0},
      {stage3_26[0], stage3_26[1]},
      {stage4_27[0],stage4_26[1],stage4_25[1],stage4_24[1]}
   );
   gpc207_4 gpc868 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], 1'b0, 1'b0},
      {stage3_29[0], stage3_29[1]},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc1415_5 gpc869 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4]},
      {1'b0},
      {stage3_30[0], stage3_30[1], 1'b0, 1'b0},
      {stage3_31[0]},
      {stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[1],stage4_28[1]}
   );
   gpc1343_5 gpc870 (
      {stage3_31[1], stage3_31[2], stage3_31[3]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3]},
      {stage3_33[0], stage3_33[1], stage3_33[2]},
      {stage3_34[0]},
      {stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[1],stage4_31[1]}
   );
   gpc1343_5 gpc871 (
      {stage3_34[1], stage3_34[2], stage3_34[3]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3]},
      {stage3_36[0], stage3_36[1], stage3_36[2]},
      {stage3_37[0]},
      {stage4_38[0],stage4_37[0],stage4_36[0],stage4_35[1],stage4_34[1]}
   );
   gpc1343_5 gpc872 (
      {stage3_37[1], stage3_37[2], stage3_37[3]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3]},
      {stage3_39[0], stage3_39[1], stage3_39[2]},
      {stage3_40[0]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[1],stage4_37[1]}
   );
   gpc1343_5 gpc873 (
      {stage3_41[0], stage3_41[1], stage3_41[2]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3]},
      {stage3_43[0], stage3_43[1], stage3_43[2]},
      {stage3_44[0]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1]}
   );
   gpc1343_5 gpc874 (
      {stage3_44[1], stage3_44[2], stage3_44[3]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[0],stage4_46[0],stage4_45[1],stage4_44[1]}
   );
   gpc1343_5 gpc875 (
      {stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4]},
      {stage3_48[0], stage3_48[1], stage3_48[2]},
      {stage3_49[0]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[1]}
   );
   gpc1163_5 gpc876 (
      {stage3_49[1], stage3_49[2], 1'b0},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage3_51[0]},
      {stage3_52[0]},
      {stage4_53[0],stage4_52[0],stage4_51[0],stage4_50[1],stage4_49[1]}
   );
   gpc1343_5 gpc877 (
      {stage3_51[1], stage3_51[2], stage3_51[3]},
      {stage3_52[1], stage3_52[2], 1'b0, 1'b0},
      {stage3_53[0], stage3_53[1], stage3_53[2]},
      {stage3_54[0]},
      {stage4_55[0],stage4_54[0],stage4_53[1],stage4_52[1],stage4_51[1]}
   );
   gpc135_4 gpc878 (
      {stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[0],stage4_55[1],stage4_54[1]}
   );
   gpc135_4 gpc879 (
      {stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[1],stage4_56[1]}
   );
   gpc1163_5 gpc880 (
      {stage3_58[1], stage3_58[2], stage3_58[3]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage3_60[0]},
      {stage3_61[0]},
      {stage4_62[0],stage4_61[0],stage4_60[0],stage4_59[1],stage4_58[1]}
   );
   gpc623_5 gpc881 (
      {stage3_60[1], stage3_60[2], stage3_60[3]},
      {stage3_61[1], stage3_61[2]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[0],stage4_62[1],stage4_61[1],stage4_60[1]}
   );
   gpc1163_5 gpc882 (
      {stage3_63[0], stage3_63[1], stage3_63[2]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage3_65[0]},
      {stage3_66[0]},
      {stage4_67[0],stage4_66[0],stage4_65[0],stage4_64[1],stage4_63[1]}
   );
   gpc1415_5 gpc883 (
      {stage3_65[1], stage3_65[2], stage3_65[3], 1'b0, 1'b0},
      {stage3_66[1]},
      {stage3_67[0], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage4_68[0],stage4_67[1],stage4_66[1],stage4_65[1]}
   );
   gpc1_1 gpc884 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc885 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc886 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc887 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc888 (
      {stage3_2[3]},
      {stage4_2[1]}
   );
   gpc1_1 gpc889 (
      {stage3_3[4]},
      {stage4_3[1]}
   );
   gpc1_1 gpc890 (
      {stage3_11[1]},
      {stage4_11[1]}
   );
   gpc1_1 gpc891 (
      {stage3_33[3]},
      {stage4_33[1]}
   );
   gpc1_1 gpc892 (
      {stage3_36[3]},
      {stage4_36[1]}
   );
   gpc1_1 gpc893 (
      {stage3_39[3]},
      {stage4_39[1]}
   );
   gpc1_1 gpc894 (
      {stage3_40[1]},
      {stage4_40[1]}
   );
   gpc1_1 gpc895 (
      {stage3_42[4]},
      {stage4_42[1]}
   );
   gpc1_1 gpc896 (
      {stage3_43[3]},
      {stage4_43[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    reg [31:0] src32;
    reg [31:0] src33;
    reg [31:0] src34;
    reg [31:0] src35;
    reg [31:0] src36;
    reg [31:0] src37;
    reg [31:0] src38;
    reg [31:0] src39;
    reg [31:0] src40;
    reg [31:0] src41;
    reg [31:0] src42;
    reg [31:0] src43;
    reg [31:0] src44;
    reg [31:0] src45;
    reg [31:0] src46;
    reg [31:0] src47;
    reg [31:0] src48;
    reg [31:0] src49;
    reg [31:0] src50;
    reg [31:0] src51;
    reg [31:0] src52;
    reg [31:0] src53;
    reg [31:0] src54;
    reg [31:0] src55;
    reg [31:0] src56;
    reg [31:0] src57;
    reg [31:0] src58;
    reg [31:0] src59;
    reg [31:0] src60;
    reg [31:0] src61;
    reg [31:0] src62;
    reg [31:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [68:0] srcsum;
    wire [68:0] dstsum;
    wire test;
    compressor_CLA32_64 compressor_CLA32_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he04ccfd8e90a643a819766c428ad380b0cfbb196da3c2fee0f2d083cab825335702891abd0c9da8c632f1d3932fcbe25d5a97cf83752ac3bf35ac78e616d2fe886de19885988a3cdd08b631d905f9d9635ec6bee1c2e6328f6d3671498b4d5df2b20334e1c4a724433828843ce07e7ccbbf677a596b3aec703b8a1833ef80d2e493b65b2b7cf9cc7588ddfaf1197e5bbe511d02715822439d6497fd09289142b2dbdfc6b1710b057e806a77fe510c00002512d57e63b01893bdb85370b3b9a5eaaec4d0ef9dd0f07adaa06d8d615eac7911a794ab946818fe3a399e320ec9df4fc33e379f79e47970ea2c27c9d476a03ccad5d26b5e7a5328d818e6be62c05a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd5f3f1a60d8a3af0948d0194151e523a0d76f7983cdb3e61d1550b86dca7ce8272778df87613c5934f560458dd54dc034bce41b77ee4c312b30d7204ea72edce9e3084826d4d30ddd13e3f4a446437d09c3be5edcd54f1d2631c74b92972797fc3a602f8081211ad42388299a03b192b63df3c5562b5a4c443b4537b2d1ebf0a21feded2ca4afa6659cf83dcdb5655755649e7bdc0d8f3513ae9e97d851717497166a89de86e45927953cbc5b77ee61159b8f02c82ea8747f9775f8941ab5e1a71bde9e94235bfe89ba84022476631771ba84e568e54e2d9731a62b4fca92dab5c6279a5dcda783e289fb2cad9ab24dec8be504a475193097bdaf9fc9b9150b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1a581e02b2b68ba52228c9e354b3864f5d9caa7e45012d80241ddfc99fdf71568005aa6bb2dcaafb8d39af8ac961c0a11ae0749c224628a6a68ef047148abce28bc496f679c4cef5ab4454cd7592ca1c38a2f406c2d29b7d7267c263e3b7197512c949cc2e180dd3ca179fc63f653b4c165addbfa83baa326dd135eff2d8a495e31785dc46dfc9c53ce8465084b68180fe40c7b5f3a9f837512bf30d27bb85180a1a209f812084ec21b0e38b6e2fe6a4d615ea5b7b5fd1683a7270535658a3c52d8bef6810cd1ca1df23861ca6e414860307052c21b81703387046e17cb5077464063ca9e5c12d57a453a2ba6389982194956f9810a5bea2f4c37c0d4183865f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6b658c1ec1a1112212cf2227ed82cedc5f8cb744685a1649cf91538821998a985ddaeeea16661894113c366c1cb2dabd5a383c60d2a9486900e05dfa04ea763d789ce7324935d2418b565ed335046893f161b2738f17f82067ad9743d887122cbf79571d3deda4d042b8ca644749c62a8c00a00e43a555683d577416f8057300cf835209bbddb9547256869346804f8c1e2259a75f5552e3062cd1d9b9a7fbd1f9b9640fd510ebb27f95cc4bd436e5de8571ed758bace149e8eb4a1b48d1709cabc5b933f50ac0e64d2ea582e388c4001cd108a738e003159be49cc6deaf8a732aa0b4ed04701c8f54a52dda10e5586e09cbc438f8f9e76ed6e873c77b8c2c26;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hccccbcb0a17e04ba2971ab4e2c991f53e48349b7446c916cc4fd7d6bc16ca41e972cab745473c4a43d87e87c60de655fd9eec1f546fb67812ed00e1c4e642d558c515e683ffbf1fa256e3cc2ae820a087f3f11e3e44ca67b17e7132a46605bce2460c623068667425d3383c64244dc33ac8f654580f4d88cb1a946c20c4277555af7a0b624fcd73baefeac851cd56724aed61aa8ec0dd04e6f82a30a34a16ea5a222f94c2a714805b1e1bca9aa9fa34af8c038d350223d46269c2e071e83f696add36ec670f3ce83066ab9d0679b38f38b02be2a8021e207b139420f7305e22c56e292fe7f868bc3ce724d3f33cfc10b35c8b80401fef658ac0676e4dbd4a52;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he8580875e8a88e46dda0e7090801e9548a50cbff47e6b7e8eb5f78ddccf692a213bf3980b5d313a94be5935ea4c0955ee1ac839df6f811abcb728cbf57c09741a76342ea9c94dd0d9ef035d9eb464f6a16ace83d7f3f3511000dc027efb3921698aeaefb7fd56862168b91d6a51879044975148dfed2fe93c534a0bba8202dc192cee3e3181eb20a8976525ca50a60e324755bd04b5be8d45fee390992047f266482475de14c7bb667489164d06a51155b1bdee4f5312f81abc1784bd1fabebec4f96a871b414c76b35111c1a95d46d62552a82f74f6be6e1a8a83d93ff08354ea77dae2f4ea304a07d5c2615a89d0ce16703a206d382062161257004c14a23b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb22dbcf154145af33f789fda0514e6ff2d61a0ef07af6cbed9ab82f7987cd7a72b407a0a981c0a0b6a7560ae24ed11b47e88af23a78b9d3990ebad37af35d7fb04f663ba2c0df9c9457583d58be4edabab37f2a89f72542e2b60f2f4927fa0fbf19b11c7e94104b62459b0bd2bb41a6cef437c253c1babb11a87d79267a116bd0366fd0d800023d177099e50261d8a640c2f6387c5d595b3f893ca08beae6685d23eb75e8610ba85661ddefc61a1661ea14fde8bb7929a5e0cea7634d020c9e38d8ae544448bec033f86c150748e3e7b9b414d5e5a0d7fe3fa5fdffa0d69e4e69006eed05e6eb26a5cc1c3711922805f2419d1ff0e79ad260e0401daef574da8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h771c7a6433b4ede5f13f1d1eb8ec8cc50a0d3670ccea67fd947670531defd02a65570112a9dd6b7027ef9c281f88e4876cde91d8e35d75143ae304e5ea638b24e80c96427a5ab78b6d8193f881b183de956f844fe5298ae2835fea5d693efe7d3cb70023a02abd626760484894058387b4fbed014dfafbe79472838e7ed6669badf7a92c0c803eed8e60e1ad2c57d38871d1704fd7df2bfecadda4d314a1a27904009d44ee7b13034e0c01bed176ce390b23f7e439198fbeb3853748754f02ee1623829dbb0943442964d1f479c3f72acec0a528935d6f2017376550f71d6cfef8035ae4242812572b54ccdacebe1d17ca81925b3f5b7533e608a1b309a81387;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h25d681def7ada8018585e555b1fc7b1c1bea4fc1146c01415fd07d6989567bd3bcbaf20273cd83c614302bd08d725d61a8080f508ac1b17a193c88e45d06d83430fba3d4bbcc0ff8ff3f73c49b53238a57015cd5c44bbb0b29ebc059bbd75d9f649224bbcce3f5a178451771ce91b22b1ebe002e8e2373028060e53f4f144d30b2c82110ae472c6bb4085d17c0c38a512f38037aef9ec23460db676df6fded04e3d40d650487f4e663f653e14cfb21c821980105ce0dd0a3620a9d6c34754dd9fe0e9816f39a9eaf2c3cecbc23de2d04c658c201e4b1d7fe13a3278e800be64efebc897713f0c509443e17a1f79e8c4bc007bf56e38df62a45ac22f10a2db887;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8923764d8a07d149f2e92833683ae1152eb34ec62fef228b538c3111f0c8ae9084e71193049ae5895b4e2d2fcc97138ef6f7125572c1e2e2bd4ebda8b8bcb6053317cbcee8db30ad7f216b51460eae66baa8d944b998b89ee865401d1009750f02ceff8f523cdf4f31643f2dfb0029f1412a9c33f526c748da48fbe602c45d85463f5179eb482b645fc2546476a34b0d095de35db9c167ffd48eacf8dc998fe3280fdfeb19b6727b4054866f7c623aa20d90b5f2d0524fe07b9529b9b5f60a81b82c0e79f94c2d5c15acdf61f6a4a57671475ee43a8ea6d689f70009bd3f571c7126879bcfda12d9a6f23c6a9e57f285af3da971ca1ea8ad0ad2aacd157a1c0e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h169b76c862819070082a9111f007a89e0aace26ec4e8e3b0fe26c6109f84976355056c8e5059a1665275e3a1c8e7ce7d467514ec4a59179ee3d67f96ea97dfc8572aced06ec431cd7f909785186e58dd6bebeda26102d759414617d758c10e9fe44c550ecad3d4afd1da80feedd4e8c57e4badbb3919909c63c880c33451145e792bba00f5d818e2d82d3f3e2eb7f91d299b7251b6bbe13c1b68382d822a1c908fd5dc6fcabe1c7840a99c8adfafde7c23930f3d0ce4296a3747759909b4b58e1ace44eb7ad0c9858de60339c9089400ce8e0085487bf2ea59e7d9309900a7e7783c219a1a092de9f51f3217e1df63cb4b5aa7b5e4dd09f3f66c04388345ba49;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha4cd4cd6236c1c3d8b09de10919ff11b6124773b608d2a3f88c9859777c3ff011e96c38840279087b95112ec2d3316a6943a1eaf53050aa9b5b41ead68f448e9181c5de011fc3b08120cf20a02ed88208146ebfad172af21ff783ad32c61bf2c04b1e09bc42131234013fa6628f22c9e6d0d45dbaf88f89970b225b99c5b577a298a1847cc450c25d80254edce7fa30d538d4689ad71d5224cc11f217de22c8dece3b36c59e7428aef45d0870393e3c875478de4270ab045dac1110413f026886e4209d8bb96708eeee633f6de4bb565cf7a9f343a834094f82133db3cd0b5bde8d545056f6f61d7c9230230fe98cf8914f25fe0b9201145df7105dcd88f906f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h51a1aa2e78aebec7f70c6c2905a3fa3687317c547a3d04471266a49a39282ea9140ca03f0046d42e12167363d8364a2d57b88dfb1acecb47dcc02c1178791c8ba40ae2441a39ae9ce47a2eebf357feb245a0d717cef361ff966fa0789b3fdf434619575f07bd35dfed67fe5979a0464d9468b20a2856f83ef65ae5c548dba3ebd56da5746af7a47d181fb04f9a735754121e74e0c39fa7ed22b847d699a379491699f55117179b0d211fd7846da034d6dc882ba62c12eaf303f382bb020d5ed9fb69eed43d582203235c36ceb767b222433439244cff47c7c6a6741c9d537dcd8cbd680922509b97ec8abb19d89f05be443e02708c2dfa73e1cde9b90a121a6b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h87ebebb6d1fad6f0593404fa6601c507eed9d9290b4834a33ce262fd403089499ba71ff818911f0291ecb3f96dc582ee67741ea020fe99f89888ae5044ca6f2e08a61d42d382d8bee93830a97a6be59d27823dbf1d5962594aa8c0e209a47b80932b616bb96b8e65ffdd6e448440b7592c10e0801741ed67dd9525f1f4a9b04a1e81cf729b72efdd9329172672c37c55cf77da2d1bf16beef9de218f68ce053b06c80bd7e99cbfcd9ee4687e07ce604896ce7429c300f0d15656d215366b2beb0b5dcc3ecb73ba2341e0d161e0135c8204882653118e1bb752fad6e0879f228d5a77aa598b75846d19e90c10d7a7cc6400f45aca6f0b5bbb97beb73e5771645b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h70957f1c7ee419270c8ca0c33a49529aa1e3122b1e8fe75b649b9932c3218dfd03aa5e5325ca64c6b72398987447a47fbd428d85f2d198efc8afb162218e6fc022ef514300e9b3b11f5e9daf814b6458a37cdb567804f97b622378486eee6f37fb74955f537601a0e2bb4ece434c7a8637e015bde86685e084c6af79261874487f0b3d6946aa6598daab816b87d89edfdab452fdf275c6e5fd582d7cbb4793dcc3b3a97c58e2f287481c8c7779901200ebe30c8e6d87dfc457d32416637228cd1ec29b3d015ff0d6cac53cc2c9c0b7e573fdbc5c99a8ca105dfe1f9b7757a580da1c61433e24609008a8bb3cfa0feb1c08ebe9afe23971688ccc811f118155b1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb6bdfb598acfda66cff77ed99751ee125d1b9e383d79c6b784404299b6f88b26f48bd9792a871e69986e7f568724f45f2b846462cf9c6886f1b012ae877dc447a4452fcb14cf7fea92355fb16f6197ad48f9cad12e47f0da9c06573403dc21f0f8422ad079dfb188c7a5de5b8559a3caa51e43340c9772fd4d95ed4b471be6f89e0088de673a554a50710ecdc0e4306d2a30e19633785019595b70e40a6705b516d9069491690f4d298f7c3b14e26b9acb43e278ed7c93378452db4a642562f0d1078c736f29a6ad817c5673e1998a996fb5313e26a93d10cc5f8d2267a33e634a55ede55eb716246459cb5252f381954957f2f73b32b4c32f065732f1fd3fab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h91e9fc2581f1fd0b79afd5900d7460f93fed44cac900d6119ee251595ab6d9cb938cd91b7603efe4fbb984dbd0e34d6fdb7406dbb20b8d18ddaa7688d2643033acee94693b4beeb11b0883761bbd08168ca88dc5bc139f20241e7a1551284d07057ab267b451eebb7fb2b1caea6f4f85a709390862445a9a83c8b38ef3ba5e18ad465b3d2df51ba03c3df0eff8fcbfb401e8317b5260f76d1c5795354fe23051e6b9425f64682617e8462422652eea72f5ab20f27423c51811c2706d49a35ac72ba970ad56a8fa223b36b4d66a5d204dbd66848b8eb88f8a04471f4163d58b45492780fa61feb568fe01ad1da2c3468bec8b49c0494518cedd5b3f35a1dd3060;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb361a25dcb6f0f49123c9bb0db5c29db9785e49dbc5195ba029ede83be76294a7708cd01582bdb234cef2c29c6f06aa17a54194a7b540c50842a2b56fad4e1710e282609b93980b118bce7573a59a376fa374e5bb74918b1bb0d6bfd73e0e8c5fb6482d9960fab8f9e6ba0eca494fd75a55873915444fc7fec7f542fa765ac67a16cc4552047913c1b25c66d6c82c81b5904e909311ae22d17123a588f60c0886cefffde27f6510f87d82954808cd814051263e06a9a0f210ba4990502c903652fe40bd62ce06e24a245501b7c30d92bb0beddc64595f17270cedca929a6f11053e3f5cb072399cbcefce83f2b661070dd74675bcaae70ee287c970efa03711b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4e98af838f12394999f67322e5faefc211dd755e4fe1642e5ecd122523fcd91b9377480b25e17bedeb20cb8299d1f664907b740e48a5c5811500317332b87db38ace510093807eac4173d3be5a15252da969fbcba5d56685a9633be5b4a70480e4a79040517df0aa7bcbb50f25fa2c4680cc930285ddf8c45b3f764273313d046aaf3f0604de9e390b8e660b3a90e1469010e3790c10729a6fae7c9731b9dc8c9721c3c5fb91d943a022f30ac42742aacb8a53016edf16fe474f81630570c25bd13bf4c4e943b0d6691affe824b0891a592e7c91a1e5807860738af5e425d2ba73ee65a7bb004991326063cee9b3f65b6258bbb5bb5569588b5f4ccf1b23232f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36173557bcc0dc924b6a7ab667b160010bb37bd5fc461b018ab94ec03a3a06cc27f60d690ed3670ece327428e72cecb5c2b13cb896e0e2fc0185965522fcb49cf737d5d97d6b466598fdd11e182c93e0e51a04ed1a474989492c625b35d92b7c333360a023df6c5cb5d1623ea628c705ae402b5175595b8826b8ae756aa574f4466423607a2ba1770ed2e3211ce2340b5ee06446d64b55e25ea57af715450d4ed99735692e397b86daf1fed6d238f9ce154acae38c1cdafbdc4adf827121a70cf781ea0d508ad254e03c6991b22543ad18f5f51bbcadb0942503c200df15501547d7b123001aca3cd9b8be38fbb4402278e3baaf67333cb9770323b02e6ac557;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hedd5f1f6c7a1f2279dfa70787d7583efab9f8dacb63c9c07297cfc65c42b78493f1b83e5c29051a3560a413fe55e5495ee35e453d90ae9546acf07ad4fdc340cac7976758497f8ab5d3c442a788c45b18b5b1fe112ede9ab6a091aa489027e7b7227c191019abc19d81ea8875362d07a9b57a339369cb6939669e58620935163b65e7362c5817aef41c89e3a29c863188c89b2bd28b045f8b399137fe42d764cd462d5220370b4b2611cae7fdea90d0d155312056c554df682be45e6931bc25776a2ed51810650ebd2ef810233cb0d82297fd04159fac5986c7ffb5f0171ad49205dff96a0a5c30d2160c933b80e30e01f15e50c3c8dde44d7053e3292396d96;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h92477f1229ed94e0e065ed56c957d0102c8f7c88e6f5078ef595064d2a785ff5862f926180b8d6f2bc3d1e7c800e14d909458b82c7450ac1df7582e1f0fa225b14d507f931315cb8aea0aebe474f01f6b787554cfff812b85ce9e4342dcf5ca86ce36fc568c290dfe230f08a09c06ffd06bd3443a6691dc3ffb25cce260e9ac9f713e75d68b3c363e28327943c96d41fb8d922bbd20bc1d6cd358d8c3710df3e5ef68b1e906d0897c85c02d885f12ceec8a2162b8eb970b777cb411e4520cdd1b560966684a28d0569480220d041aa09a20f6af09301a2d294adb37f94571b11c9a77a1dcf23524ab3416a1023834b92d1df621048fd8ebc0c5c78b472bc2bfe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf65989b184b0fddb8ead3b90af074ae8e1a5ccac59e8123fc800e4f04172e10b78c566ca36bc2160dd9612264a1c2e9fef71d1c1588408a39ab27badb37fd14ff64e82d06479d963b3205d1405520dec5c683742323f414659f9b97bc75b381d019efb1ff05396a505f3c115ff38babee0014167e49487f990f11119054b8bbdbc39c9bca915df9d808c30ca6002982466bd71a7e3a5b1b923913b0598119d18bd42839168985ddd90625767bcfb6150ac07a68e6b52480194316d59474ec089b248cd598e51bc2b93e00d348cd007d89fde952cd714aa7e302b9008931ffff7c0e22adc943bb387cc953a27f0727bcd083f0fed5b1f476119691ca9da50b323;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdad1c29a84c0f61774ac74da06db819a4fc3e3ad88b36f3df66d16fab0baa5113ff75dce159a4fbdc489ef8e94df46b2918926d27702856a722f3d202ac7957baf9853ae46b7a997a0089fd3d057a129d4bd64b0f7ec6b3dd3c58a1728529d35057d77d28a43f4acf80e099d26320c9d20a559801e4c9f77ede9f78378930daaae3857195c54abdd431a9faf41ae9386fd0db445ee6f641514be025dc5a3730150b517dbbc647f631c7e79447e398ead6d4ac6e7d73c256dace834b7434adc2fa4a939fed956244e6a5f43be3b492730867b0bc868e5ea2a2c1ead9425bbcfb85f7fe01d8bc5e70a1afdb9fdebce2963be444c1b3d4de582dc6b0c327408b597;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h214ce024e1401bebd9d68f480a44144bda1f09936d0dd3c951acd8628ddcfe93b40a166ee9898a91ecaf2c688e07a873d76bfb80b2a4778dc77191065572d475fd50ebf60f49faee84416615d8267b3ee00e92ad6b66479afbb143ca8cafbc21e9912cf093a687a5184d9dd0bb87c1d96e1f0734ba31521cf01d160ba50f7c2807c80ffdef1c17bc34544e08734f2df764e4472b74bf6a967a08b7eb67db120d9a89b6efe43b2cbaf7bdc0c58c6328354fb3f3d7c20069761e5db6bb6e7b08df18a7de3ce2ac2a0706e15d3ab3908d3caf731291228a68b3d18d3f874135094b3d837bb6d3b40f611f6f5fb47b00663e73cb1acbaef16d41d11c3d3540c14f9e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he7fd1b23462f6cbdeeb3d21e9ce7b04991b016c635160df52ceefbeb3fd508cab7cdfe5bf41f219147d73582162e790866a8616e8063352e50c82568b384f1fa9afff73d52fb7bca36e8d2ff6c7df2d746035541a7e9dfe977b72654e353319fe72af6dd44ea29a3980bfee6c97ec44eb4c5fe9c69fe4fe49e182b3e3da8d1d32a6dfc5ad40423f21d670fcf50dae2dc4891f7078b1df11ca332bfa15255580a609716303a6dbd6fc9a984d1db7f10a06f9caab8c0795fb806a456625c576c06d63f7a97c30306107236de2dc11a3e5fc1605f1f64fd5627c94635493ecb1b414aa5deb1f508f67d9fd150264663e3cbc71485fb1ecf29f0942af7e361f8a054;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h664e8e1039c4cd05c00d0027b7ee3fa8e72035f267d7c2aab8f961f34d750afadf130140825943dddefc96b2ad5e6b33c70b0d8366c6e4e14a3c510fb7cb9e6613e35b537c2a6fbbe304d6b53afeecb40afc429849fe7deb595578e0cb1e193c235e54feed190ef8b89640779ba013c50a46b9a4094a501b5203fc359475d6ead8f95f6881bcaacdb3c47011686c8a0f38ab11f5fca19d6816113763f4853f2567011f09b0a5f79f4f86ef66ef4bc98a225e348625ed1c6029afad0af9eeb6299c5a07bc0c289dcd9c5e529db1a03b4e68c28233ef215d857bd3f2af0417789cc870247e89055a1ec49817bddc590f7b53d5f10c2463bf1a913a280aa5a879c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcc0d14abfeb5e77e64875d6fecabc9da969a4f97895616f5afe3efba42723540370e6aeb16bb44bfb7c5ddb8f0a01186c8760d65767c8cef1387d67fc9cb8da6b4ad9574592d898b435c21013619cf60088127026685d810b6b79b4d7c0bdd8afef016e3417a694347f5bbaa25803946c58fb8c3dc2c108f424227e46396c33b27ff02107414f1fef678b7493664a46fc36eb899e8155fba8300d04a2687e6afde1eee60731338b4777aaff8c333636c7d85457c448f8dfaff9a42c5d8089fddfd4eb72499b60a2c1078860ffac9666043b8927217b507c43684120f7f112bb97afddd2264f589b4747aafb0431eb2b56878df3cb2bbaa8ea5f6e2522ce259e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4120594c846d0792c75867eb7b13d094493bc98ff9dcb5b8e85fa16168df5da22aae29bd06f55fac1687a680b491c3c9c4d8ee7d864f29913850b7f8dd69bf6794bdca23bd658befe50123a5e2c38c964f70574a0db818e1883aade349f8d1a65bf6c46b6b6f2cba833b5b60cdb721ea935e2aa1c48736b6bad989a248b984810cc7f98777dfcc36393e6b27403752d603da1937ae3dcd1aad347b330be8c6171b843faeac06e87c0c0bff1aa4ae2e56b8f7c7ef9e7897f2527d259dd8801b171de39aa2761803c6175b8d0d5e281a22eba4f39e7cca60368b85579981f7ba02b3136e402edf24495ffe81aae97d92786e15bffad993762318caaba0d7527615;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbec108ab6d172e834892b4dc4a5389f1395de549262055a803aaf9f428e0b44d158698597cbec2bf6b8e618f5ac3b00fd708345754c4784da42f6c876f56730b69bb6eeba1f01c7730c3d483e8281e1e7d5bdd742c5a08c0d8f586cf4bcb4df8c6aa7f478e61a00fded84cc440eb70dc0fda9648d75b885a9cba06938f3dc2aefbd7965c5381a7c50c655d6c8fe78d58187302e0d06f2949932ae38573157030bfd66ec5bf7fd3e5c5dc645e7dbe09551e50ac57088a53c15b3106d922a1c5d92103b1b8a2af23e9907641a0b618ade69e791c427b9205a126f61a5c17bdaa428106ce6d2aa94324a9a6dbe594e49caec2a73b109e6e02abb4b8fb0fe5250d4d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hee52da5e7090c1a37cf0e1d88d223ff05e75721f4d2a61f101573dfc8d672c9ba06691bc7f1a14e859af2d36d8a765e39943b79c4687a73c76d3a17bccee446c11555a5dd921120f3b053224737dd96885d90b6047fbeaff7c8e9fd94ca0bfe43d9dc2b1f20a148363e1d57ef328a5e1b1e5b00376876056673549cbacbda694b7b047137f96c123cc71559e296ed14882b1443378a49fbb68ba07b0ca034c7d1a4a06ed3e2b73d9ba26f2d5925a4d19f33bbfcee5fc62deaa0e0833e5ba1dfa82d1ef78ab9b8ab8407e48d99366c989b6be49a28edb2387c67b07dabc9cbc2283d52cff36254c897a25bc92cdd52ee15501f8f7da0d206a09d0b78b06630e4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h22acea046d2e43f12d11be90337c9e4df2e686de9602a34a5beb16d7fe7f5aa0c9821fa40791a91e7be40a926f5d9c2599457ca404322c9e65f20bdc5e763f4417989c16b616690e1a3806c072b669e3b32605ad1d6a980d166bcd7fdfb92e1ab6b37b84a2abd9a7297a97399aae21ef1619037d3b01b760c8a4b04cf24e7d5342969803c65f2954e10acfb373aeac6489dceb968354316d9976f706a9af071ca6eee056f089b9d6bf0db66af368cfa0695fbf15c9de35706e85814d35e5ec2762daa3af8fad1e9bc051bb4f35739b69a2c4b49bd448f5ee43487123fd047f4b5b27fc6af87c8390f2203a6e975a674ccfef7fd4afa3410a7a86febf0ee69029;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h81919ac4c58fa072bdb6884236c2e961faa11704894ebc59fe4005c609ef6bbf6f8bbf5df467e49a0f0a96e4bcc1f010ddc9529f1ffdb419413200f54fb0a75ad3b87f6c05faeb82d701ad7c5abf4375bdc468feb6199ba596fe17b2bed04f157956f41f4c4a9c1938ffa2519c2050a23e5bcd1af4df039966ccf6e125053703003e66bc033ac5892ba235bc8e06edc1f23abf9d2f2479cad421cc954c565084c2fa9470fa1b0ac47a74c9c4e2cdc537bfd117e6df9e0079ede81b52cffafb4f8c28a74b63c4b738b10c7cc5ad809f08821bd94f3c3413cb83e3ae3c843645387401a37f5b80d33b7eaff6c9d36e758b9f659f6964624f48bafb6b2cb3f1fa38;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haa18c6ef2cc7682c5c8a5099cd0c2cae29c9e2e663fb1e193de936f2712b044436a3f1ff64fcc9e210c3d47a4a6a613bb76570447bd36d8f042773426134878287c3f30585a111c2352082988d723c8c08fcc42a17fa25f7e41b326005ec378e068ddbfde7a7585875ce77f43479de1a75c172f53f1bdf513419fb23d5d0eb6f9835f913cb85844a49c5ed51a9986384d94f46b46701e6118e16a03ad333f49bd786d292218a01b91a6c2e33f5684a5244099f825421e181624bd8db7218e97d3b4fb337330d61dd10d9a6a7d546aa5ee617d4f893e3b422d180f403a9683f8eddcc936d684bd415a77dfcdec3075a9818bb67e674bfacc8322b9cfa889a84c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1962270e740b9a72be96ae7bf5e936d1ecc718c9a135724ba681c76c7c281b8f27c0e8eb891b2429c0c0955ea6a2386ee7cc576e6725cb34147a015f7969ff6300b80add268bcfbaad30e7aa9ba7a2895048fa8b5564f133812db7227a0290cb3e8d80fac81ce4e2f05353d7b35a9acba480afbaab20c6ad9cf603144620774312ac492d777cf4b3eba0f65649bbd230927210e3eadcc773e6c137472d1217db618451cd68c89301cc8eb617d9a6b8703489e2fdbae80e29a95a77fba0193f353860e730e3c501460c98a364e2dc2954607cc225191a8b82c2bf34194fabaa1c9950c7c1e55057777f80e2ba5f6b0be081dfd13fd0a9b13e0a8f77a742d6c88e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h94c48a7d296b73502b4a6a83fc1f95eb764398b894323ed158a3f12218ebd13359309f6acc83889aec02c37508691364f4a2c8ba87dd7b483556e69947002b23546629d7ca8bda7ad3f92c82ac56607595a0857fb01d60981f602dd8c924f8327df7f9991de0eb1fb46262f34264743476a6ec3c4ca3ec9f90653cd455c17cf1c6cdca6cdbe201efbff25ec02c0465801c08a78ea4a6bbbd9bfe4bfdbf0aff353652a54bca061926c1b65f192038e8da54e2a40523237198da97a669fddeed781ed426cce858bd0c6e9c32422d6a7b5c4fdff546d74e27a83c1f8879c7891029c4bd47a0c904f77f8cd244f69489fc03b0a1d0b56306afa199374fe4a94784f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h18f14fbe77a10bf5d61a8ff793fe5f8551c4600087b7dbca02770da6c0109e7ce9a335aea1894405a706a75bf8710564f53299d8c9f8fe06d395b93ef1ee484ee6a1c88d8174e407f3624fc49049264ce176dba56fd940427461657f3f476bd9e9af76602d341c3e302e01288da18e192bbf741763d1ef896a3278f4bcc1b26b4d0b06f82c85b741edf7644aae9323c141f8d2ecc0556436cc7e7c1e5062db9f88d8dbe3e72109b726f21d39abc20ec015e0570e047c0b3d396e49edbae4a69bf49a1c0ffcda1b1fab433c1e419d5d04f771614a4ef0a93a9fda8e72fcb1fb2b7a407a8468dd5ba42868d6e99857f6bdfecdac9c492ae8495543a36de1444fac;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfe5da88ff4e2baeedd56258e91c1c0504916ad25d35cecc81d58f2dd50a76fd8a7314c4eba6d6d24b70de59e74d8fa46379a6051f4c306540597e844fdbfd283ec293958c9597f5f52e3dfa22ff64dd6beedb07269faa9e4072ca3a447b3da466924aa8f0ef51ce1f11a44620032c671c7aeb1f091d18d587d1e313c378a299ed179ed1008824c4b45e19d2784e43575e8554bdc8d0a852530657628b1393ff4df0f7ca5d7c6dedd43725996c093ea7edc9a77289e99661d93a8ec0f8bc35f28b9fdc4f4ffd8a5d4c07e7bce1bc58af1932cec0271abdd2855e04484bee7d0c8eb1aaf79f57486d78fa9b315724931ad3e9bf5df3c8ce651f3a93ba331b13998;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8d876d9c2caec50e959d1080c5c3f870affda9eacea1715945c2a4e55f36b966937f38762ed817c1149a900f6a4fbbf96b23238251a40e6596174d89350bb190ba7f573e07776a6ce726d61eec245a349f64b3335eb89e36ed797881b009dcafe2a108c6066d34774567922d854fae6f38317fa11c7cd76e5cb51e642a2ac0b6113babcfbea3884fa1a041c9074abe1c74fe1bd2172783f26b68a697fde9e68f704c6b69ee0db6b9cf992ace62b4a599e28cb4ea89353681bef17e27a15a74d4e8eb26418388246af54c38d26aa06771021eb9eb583c79afedf2f1ff97c4cfb78227896c2eefce7637b7bb62ff894f9083878266f867506f6d8546bf7313f409;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6b76592874738db1d200f5093d69e6066dbf653ce667fcb2f4e9306ddebee5d5391922b6d901ef7c717869809f1e2c869cb62782be00eb43e6e090c038d5440f31c09c6969da212fc85c990518b040b422053f2c8ed0606b0f282fdbb696555ed7c45bcc6d6e3545272e4b4ded3069134ae98732227648d7ecec240aae94a3683c5b6dc84c87fb85103cdad9c2d2127e49665fc6259fc949cfb4b95f023b240e7357c2d1903366f97563a2d2f3ef8775193a21b0f4173498f6de7c197bed8e094387fb3a3c363c931711c038ce8a80b510b4002b3c39df46f2e18f5bcfe162baa816df9ad959425cbbc702a3d9b887abfe31f80f28d7b7f2b6d35d9074fcb335;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbf530d7bc7db85b45baf73b6cfae0aad4fe6130c47608225ebc1fdf55428bdba605bea60166bef99eb2cb67923a8d1f578289f231d3d97836779656c56e3e3a6b65323f70971f3276c36bb4baabf34dae2fa172c44286f7225a709c43626755a4eff6e883ef1ff0e642efdae7f62ffc8972618f6a766a78933139c0fe5c43c405bd2ca37691e4b3998d7a2e161d21ee2a60aa21ce480583e8063542db781ea6569289585b3947b07adfdf41c16a00105f6293df62a4938d672b8fdfaf5ada746abea78eafc185be97caa25c6609b60d000e13421b33654256fe2d62c3ca71fc2c100b4983dcf85e16c9d27de5e2728ee5abffd647231d748a8f176bf67f21078;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcc2572ee89a70a2f5e90fc019eeb12a1e55514e7d9ed374927d871cd78072d08c5da103eead6cdfe3974789f5a1fec6e80e8cf13244121f05a8a278aec8004f44552870fe809f02f4432270c0338fc836f91f9647562332578f01f47f959ef40be0e381affb48ee37974fe2997d38f4bb4f71309ee21fb7d300e6e3e12b53e9b3304d426f592bf76820572bf93c86cf94e71eee7c6413f101fb5532925d6e79c474b11e1973bf62c4088b511cac69f1a60360adf00f0258e9bb9f547196765a6f6ca1eede81f0aac7a6863ea87bb62a450fc1438021d2fe14c7d06258330776510ff345ab636d26d5548b2b53d068ecfa2ead6c486757a8e7acfbc97f915e241;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f763302dfd7aaea89dabd0fe3a5937963b5ea814f1143c99e7098f098ab3f4b3e12fdafaa3520bfce15e0f3cc385ac4a4c8963710e4e16ef03a57f14c9eb628f765483de892c99f393e71349e7dbb97223d4fe8055755cd1c399aaa5fc24502f1a8e02887788ac4e0c5fd65230567dd22cbacbe082ddae1834cee37e88ea5f5d6c49899266cbadcea455259843d4ccafbc217260345b5413dc159a2489c337dc61899ac88e9fde5197d10561c60466c8e9dc3dc602ebf58e60e08abd2c0bd12c67abf539e248e6f55d27eac906549d029cf74bdb852ed87cbc7a4b4680c3d4f0d07d07ce7a554a68edb23f445b22db49740252ff43fc52b5060481a929c4929;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h461e242774fc6fd672b1ef5e0243deeade45fe0fbdadc4e34f40cee93adbac7b1f22d03765599622bff1aed3328f36e31c3655b91d1554d37287fa603fc42ca6ad3fcee616a96943d15369138de851e2627ff2c6f2fc35285b0f560139072d94ef4d6a1fe81b53e1ff80a752256e309aa2d83f782310c768c76d812e55e44320c45942267edfef471dae1c02a76c3008a1fe707e48192d2fe181fd3d5cebd16d8c2f51eeecaec674917c2d9b622f97fbfeddf49aad45bac046b9a8ddd8da3fcc9b331a30e372bdc5102e66af25266829abb4f6cf46c65929cb449f519de636e2c5872ec810ddf72c3eb4d533331fe66efc1413114012255b02d9a2b5836e9be5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f41eecff9347f077b4bb7cf4d9355e3dea77e7569fbe384dffd84c6fcd7974dd8bc7d8e5376320a03406ea08e4c5bee99cc7a9746bc3fdb5a827f2c5ce641133c18567be8ebdb805d292d15f6573a1aaaa62c0ca956c674574668d2250ab2629e2ae34c5350d7a099d91b65848a914e6cb001535cc2ea8b7a9693ff3dd866b183938dac9615de16afad820508b59a5c76718f5a651c3a456dd6b18914d5140b9741f80382734e673161899cf0457aceb4015747af4f35dbc1dfdef5c64ec5c893bfbcad0a15cadfad89558c246acacb64085fa4bfb488d1267cd630c5851d41ed09f42688f9d5819f3883ea200a70717d8e6f8aa0d3aa9eeec92d377fc1ecf9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h34184a0de35a8e3e8c77dde8453da60d98fe234e4acffe3f45c98008f5254ef11b712435d7b1a17657cba39ae5c66dfe526ad8fc598cf83917139a0d8a1344b78ecf6ec14f76c67ff98bf91c4c2c014991a4d45ec6d470047a7c4c6dabd31591527b7e35f977c5971554879ef6852f82fd6377990cdb8a58631d8d2594f52438fb49288c72e5e3da3e32f7b9f8a44bcf36ef357309273c4a46fda74ba68cedf66b956167772daa7b6c027e9dd87c43a00982c1b8f7e5982f699dc1667165886de4863abadc61f3d781b4bd92a142f4a02cef9a55c7f6925707fc82f6aa2e9bdf7e156828e8059f299126f0f93608d7f948fea1cd63a5a6febaf11a3e8b2c5d41;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h712f2baa7653023e80e6232d31695397598cd820fb3249dd2244f318a78ec611d4307329d6bb58fe326acbc14e39e67765c0e2ddd7c98b342ac7a2ed991f294337372e37381f769397b9c313c4cd01a8b4cfe07cf81b6938dcc04f75a291bae42f3230f7f9f72c7ef20983040acba5119045ada8d95320e368d98ecab3d6621309a957781dc1f20236ce9bfd106cb9ca4ccf654388564dd21b62a125510723cd38a84106da75145f8b21921d064bd1739bc31d51acda23183cf8dfcb9c04d323809434ddffba4b4e67cdb50fa89d4b60db1457eb72382ce608ad837eacb746fb9efab1cfea713f3dcd8ea17fa6f4201930170c82172be8c1467b676fb592448;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8125783c37949db20b43563c676628074640c248838e00f511855a350a88b8aec551eb42f5fcb3b9a2b2295e3693e88e55a0b408cfe8670992b2de6e2ab785e3886b32d5b8c989699e521b195ed3ccb49c956931133b536a567ef429b3cd81a7604c62e53c23906b0460e9b218df9192456cbd41c0689caa87728d349fed9002d63698b74e88587fcc3e0a1db504b5aef7d37bfbfd671c5c4a48e2277c4651b5d0c7b06648f91e0fcf6d3eca392c0a83ed98c766ea3627ca5f748bd37c96d0a91073a4433c62df734d910f3ea80e164e336bdf8c152878fd62cc55d3730a129ee817d20dd86b2a79d4a698856bea594888d8e765ab4ec7c6eedee0c7d9449b44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6ec1cbb4d81359862e366b794d77e299d48d16a56afec8b964edcd469a910319785a176896d4042d2d003b73db01457f55f7a982dc311f3871556ed9fd17b5e99392f7e1ef0a6fdea7c263db213ddd6a67c711ed34001b1dcaeff852382cc570d56348285d0add0fa64cdd4549caf6595e0126aecec58e946109308f7fbee6fc8511a848f23ed1080db74f133fa953558b0ba63118f37f955e3767f0aae6cc68ba1f7bd066fb02e75329fa0ce698feb77ec109a5a1127c5fc735b372d2bd7044c76e80ffbda63420a380b4a5a70d2deeefa5f4c2d561445246611c772e73de382215be91f6274c1f06d259ec1ef4e9e33c701ae419ec1739951bdf417ea87188;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h677a76a8c2c25f149217b5ba83bc1ec116b7f6d0b22ff7740bedb22336414c2abef3f72bb7fb24f4938e8f282f6eea24ffcbef9110a2d702553cd38edf9e4a5932a89c4a4b1c042474bb73fd392f90f25e254bb3560b3575c7c21966d7de1a98311d00929adb0865cf7c99e88da4993138ba6bf366696c5f772b454efe548059af62f1d827065483ce8ee26f75e5f37c5945251638e9a02d64e0916228f87d0ece18cbf6f43c7756132e57ce672882ad5eb922ffdfe0ea4c4e0aeca6f1c836ee59fa0ab11ab6f6c94a15a2636df185a890e0f356835ad053b6d93a26e661eb07afb45e2baef922cbc8640424f36259c1da707d222cf128cf5deb20a400b8f1bc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hacbeceb0113b96b488d1bd170c1e97a8a02fa93e599b4563544a800f573f46c0e630649664c2e0d4b8ae942c93cd5cfc042e77c52c2177150b8f9d0bfc6443fd2a5f418f7eed19bd4a4fc889a5a590705c8e43a7dcb1ba285e5aa8d5638aa5b4b6998a923162f7f909d19d2b4f60946f82862385d5e793538e1dfb58fcab460ec80b27c2e91c00fe725d05ab3452c61ad8403b343e6e908ee677a20e6fac3ac8cafe0810c8c5f9b1fe8eed853d8d472f4c10c17c3ace3d64fd7afb975fa17fc0a4c38be86f36b309d7cd2bad59433d5d439bf2969dffe653b9e2cb785f585c5f1be0be3fbff07c8e7de298806e2e58c8d1ef40966cb8c63705349f7757894a6d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7611a5455f77bf9f68a14ee276cdd9f3fc9230ac8258a195b67485f642e84810c74b6db3908378b3b53bf566d4f78abe5b051ae29e5fba8ca8edab563d889243a754ed6342b1de0ba6b046adc6efd1137639ab8ff1d6cd0e97c60ed5a9673e611c170b26d97375d9da0985e36e48e2df6075820158d4b50cb28f1217788eb2c440aa217d8168eb2bb0b2455e1b2febfabc0c5a3b9b235718eeaa4f4d55e95052822f699824deed9c6e5eaf91d1e95097c3b37c05cc6d5d17aec47c4dd261cc116c733a4119e6ecf29f6afbfd237d9cad40abd38c8e8cd22c34dc7ad82c98037f89bbb42699601da2ebaaa6207a6be876907bb8a8c63263594baecdc6165de8b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h157784b44059195cbd809e02cd7afc06e28c7db6da80e33a1579f90cfe6a6e56643955cd8c9e25505896d2128ff816e1cb74f91bbcccce0c5718c20255fe784f1a41e15b9ba39687cc97277d3490b65a8bf45ff0c96353da81103884e25e4543164456103254c87424d16962abf54d198ca6632122f9c061528cc251e891bd90bfd01a7b9372e68aa19ede6369ed5a6f5129ebb5fd29c78a56195b74e64efbec1493465332a03f19dffc59a7c07973d2f55e1901c5a6aa76e75792460c16444a608d0fc6cc3a22fd25155a23e0235e34c0fac7ac2a56ab6036bb80f530f1fe297ded64ea9261b0d9d34d906b1f13902b76be40297e23506b2f7cb6748e532326;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3e5fefc2ef6a2a6edd67e205fdc2804bba59ffb9c3205ffba11c9918d0e9702c11fdf184a06b490c75f19a9744e02b1a6124e7e09df56c4b5fca2c671c32e62841ebf175556d789a5b14829ad57dedc96b9643be4c57342de6de9f0e75e75e14d39f8fb24f93a90d05dc966bc9d8256da24e5c0784a1de089208cba65dda16482786a6ae82bbea508fb74ad84cae454796739e1c77481225d3cc84c1d8337491193fdc46631ca90962d9a9ac6d13b9e1915246af70037beb0b7a4a000e1e05e8d7e517f0b0c9c75ca7c19eb66f41e362ec330a671ca54fb03c1fc5ee497989c828340d8b2fb973091961e7851c5edbf69a00be5959758ce8ab70513f208501d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h88267c3c13d03fbf92ad8a5e278acb8a5e54fa3a998e073b380063a0c88e17eebadd1c8adb37cd6f14e5b59ced0c0aebd3013243266775c92d63f641b424fd411f8773961ab78caf506d8f95289e403b592290941fe80208a8bbc6b60e26f0d3b5d9f6567380dc860f60befbc0e1f1dbffad83e9cdb713a0db60aa62db60a36f6533a2ab116b3210e641eb9142c84019070ee3f6d19541280ad30eb7636c4e25c6607b1ebe9c2ccd8c27a340e8fefa3d4281dff2270b0319803f997a1faab080476e9e1f95efbb7027e02e30227268a2b2e55bf7f5c574fafaf08798cadd6ae32d6f1ad684206608d1a041cfe0c658247963067d67a7a40adc2615e62bedaa14;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6aecb208ab41f9fb564e777bf723bfae85d0e2b9e0625a0ac0ce7908e8deb3f35e5e167c42871b51a2e1dab2759254b59e04b933f83dd5a99f983dd824334d10b23e9cb548f91a00255652c508f412bc656d0c137e8e216e6af4d5f96c94983e740525840b0a4b620c25c1b6b7ac66a43b917147f2659ce0d15584741a9335f55432fdef981ebec68fbdbb446d171cfdf040dbdfbb3742b033f9d9fd04804c18d0922167855f72dcd5820e143f260e570a2d9300e25cb4a144b3fec8807ff92e45adf2edf98bf3215c5803f6284c0fe46ecaa4284ae99b7a3fbf6b7153bd2c5d33c580fd7435b9f3cde81b892bca27d58fa847f2a57bafdc60b8c578c6c19caa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6add660e519645022b53cb85da723416fc95bc08b1661d96c158f0a025783773715d08a904de74c7ef50282477b522c923c2ec17de4d76f365e14449a0ddabb3689d5ff3a1386ab19dac198e48b1d1e43e9a8ec0f8ec69c6b754b748d3a132e212be110361fd82ade413756e223e25c56a9eff66221ce7401e4247915b13baae2243f9d9aa1712dd1cc1cce529ecc164336bfd46e96bbb6c3941dabad670842f6c87bce9c4edce024dcacd1d5a472ee2dc3482b33c11da244ee5b0dd0d2ec8f6544bfb8a0f55814960a2caa6dd7d08d8454df253d351563cca8c870430bc893b7803d6feac8deabc678f858c04e0bd07be0d315608c34ec5e3637100e09100c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h312e415615e2a110c30cfe183fbc49823955689320ce6eeee8dd21010348af93d36e165d536b801674311de2b4dc5fd74204948998002191262fef973968131d38c7459b11ada4757c93b41cdd92499cc8ecef96bcd0acfd2606803c7f6dbc08a8f89a6e91814221abb4f19442bf491a7733dc7d8472c5ffa2bd869f561b21a97ff650994081dfa7908164e3b2bd59124898514aeb1d8b362d29a92d39a955c76b2429cf7054e7ddb607ccbc44ee03e95e1d12dd7fbc4dfe86379213a4233f07d0a472f046aa5007c4ee533920a2e703c6476b860b10c8a446f04be53ae21803558f27afacae6ccbcef9f5fa82172a58915cd0cec15832d60502dab5c9768490;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc4adaf1f7fbd614b014a32c7e446eb99a38400270d50082f83e08bffeb7643c30789cf9e96c3332bc9993a1d8747122754e5791008ef8522cce7d679e1cf3f7cedcd34c876e2b98e7216a58b821f3d482e858d1a8459d2891b58616b1a86d3b9a938cdc03891aab9ec61334061e5510c80743c14b309d1b1ea36a7fb9312f30238e55183d4aba69875cf77dc1398de1fdcb595d527a3c241bfc75b3cfcaca19eded7c2157246fc563cbb5ac3f2d9e626c508f54196c28f59e6e3c886e2aa5fbdd5820c43bb3cf1341d7689db7e32e2a144e6b9646b017c66b68f65e6c8c8dd43e90ceaea250731f7236e29add84ca7fcd25b203cc672b7238bcd8fa7881d899;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f5b9ed938b3df8e149e268538c545515d56c94e4e80d2c93af95aa6e4844864c1c342648154117d5eb3b729ff3dfb4abffb65a63dbad8922137f60bcb1c64b4edaf81a8364139864a7a0ee2c1d363fd678e00ade4e35f8dfcd614e9da054ce72cd8e8e87dddd67a024983b3f4c2878e720bb2cb247751429f6d12cb7787706a6a50795f20a2725f7d3c34b1e56665f3e3efdac7aa8b0f2a1be57d08ab88ef5013e73bcc9b0f79c42f467402c3e92240b7ab0f20acf083f37ecbf857f37688d69e4db856ef1ff81ccd485e3ae6a94e369a3720f2ed0e588eb33699ed36fecbbf9add43ea348dacee38bf87f633fb0b3d98f17b9879471cbb6f4fb9becc432259;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1d98c8f39125643f8dba1eb33bc09266cef47ee159d95ccfe6d99f9794f1d5b7cd455c90e99b20f729f6395e635f192abd4022cd2c96693e127a6c954b64fd7673edf70d019019f3097673328fa37676b6ae8304c2757bd6ac83f812b53e6956cf2ee7cf6ab27c29a542651ced98270202fb5317869ea6a55a88bf7bca07816d1e8790fb8ff96ac867905609ba0773b42c6c4734a5ea12877ab7cfd3389c7fc7a359e3e4bed3af0107188dd9748e727bc43cc2956d550b5608ec55f43a71ba859974013bd34e271c3d1e66bcf859c79eeeb84f10278a20565cf44466f34d3ec1c45a4b7aa0ad386c4ba4a6b38652d49cb02301084bdec20a952abebf08002572;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfdd078d25ea08d63fa4fabfb3c7ff4044103460004b1948d4be9672077b370bc4ff3b1475a37312e746d7e458fd040f384beefb3d424bce3812d121f1ba7c6a1f61c5929f3b6ecd8f06d88ff6c2ad07e8ffa0fdfec9e4294fa42b6f8458864e87222a4b53aa86fd5e765b249fd7056c0da04a8b8ddc796d5013bad77404e5f6802c4d67b76e0ddf462b177144d1e53123f84180527c7b1e074dbce0ea1c8b6f379d81a65faa546b7ec78bc51e9ee911a791a5b90c8d502e7b5f20181b2c544d90009c2c88b928abfdfb835cdc3987ee5b83f969433098571967cbf70a1f1a3526d7bed9687bfad460dc2db983b10fa341ba30146aded5f4366377a88aeb2ebe5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfd000832ffff24a3ef4273fb745293029cd15bf9874f3c1fc669960e37fbd6d888bb59c65dee15a04f550a38b2bd32e3fba4158baa3311d94aab55e1e6fb3170b032fc56a9c2346236d3c8792bd7c550a371d5a27a8b917915b88d1a17aa3731ce652d275e0663cc3dfb6f6cc2e7f078ae0b741012d55f594f92d53cd21833c0e10474009acf1ad98e2a71cebe0f995af39758431869f320a9942dde13f29d7064fd7c7d5c574f59fda139d647c173a6f954c5186080a15402ee9431ae63745725dd3202d4715bfe77117bb7428870c233bec69895eed73db73f3e4eec83fb5f96ed5e53472f1dadc4fe941374d225cb4c1b939d0603f0287dd92b315b4ed8ce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4deba5827413d216c8a90edf8c976183ac55040498dece8afbb6fba92fd46d2209be1e220cc816b7e9cfa8f6174eec5e60cec7773a2360d5550c0a6e8475da78148a71cbcbc93f9001f314ab264bca57b6e449550eb7f642c32e2d1515adfabd7b14f0499bfece1c009e3005dbc8f7455d922128aa83839b6df07cb3c22343812e626fcb59272aaa217c0e3f6ca4e702ba425056b2dbabf4bc3659ae188ac2d47e74b17a33049590dc6ad20968ef618db22a054ff90ce3e1b9ea9b5da5be93550ff4a8e6155fd45e7478bcd11344b45a4b7889257aee9b4a62bfc48a41fd7f73a0e31114b80f9dff560657b2dda20894baee47dc13e5f2bf0009723a44ee9555;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h64343f40624f25f538b87ce7fe07a6a799599c3ba2826433e7ee6da61fd5fbdaaf06b037a7c972a36f4354700352ff1da1784e096cfda24c7bfae5a39c9e6a3c70fb0c62267427d9d1683030abc2c6a6f35db975e988b61b3f30e52fd9c4242605da178ac925b79cdf1adad0f52ea64f1fc43d08c9ee700886243873e9007f0ab8313c5a3f9915955087fcebeaa945e22c088ca97d32683babf3d39720daf68c5ced7f63a9d5b18bb853a76910e8490159a8bbb8c7b6f06e28fb17997641d04e83ee78fce7fc6baba488286c8c82cfa7d4299677e86b2ddc0c2eedee225823b9db85a5d9afccfb8aa4661725b1b23c2725823555304ddc88dfa7e2aaab4baa4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8bd7c913f5a53e024231dc0396929a668d569e3c98b51934e013735778416072f9c1afa6987588711df799d3f516ad5e937c366bdd6a49207c046e049910a8e7fd4edf2311bcca43fb6a2a2c9ff967d444a6df4ed0a2a86b31cf5f350fefc38021c313c8042c39ca7b4008239ec3af3e014e15de4a0ad4cf2db1225fbea78b730d2036f6400b3c3fb1a9e4c68c387898bb4385dba01eb9ad645d8678989490edce1e5f436a8fddbec420cb73d0dbf87cfa1488d086a3d13557e9abd1dea7644f51f1c4a7d4ce27d8c542ba2cfb433193f550d95ba0aa9affee3986efd990a32ae14873f43468e291c48e7562a63f37e96d86041f87f753e21c79101ccfefa309;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h91aac24734f2afd1b126fe97d64965d8278c8d8809d7d95721af0a08dabea67a8810b9fdbd6a9f6faac6325d9c15e0af8fce357675a1aa8c8083f241fb91371aecd94b286bb4b262cce63b04cdf3d05c5e77a53f8a0dce937c67ec9c06ca9f66d5c7bd6312a132bdc57edae6a467ec79e53433b6e4ece9b28a80a1e6129966f7f77f96edcfdf18904e71b8af8b988875d16dbc6fb89baa0d301aafe130fc38c6582643cb8b7e73a3258d21ce589a76caabaee924f219d287b5e48d2212e87779d17162e42c067f333b9786e164bb7df0c106c5142e8e57a0af8bc1aad26c10dc1112a1b73d458a6b5f84ca4db12c6627238eba0d129a457f3af2d9dbded05ba9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc30ba10e84288e626fe337be893db21233e3e76be28cda30953dc3c9486402f27dfdd4e672e3cabae7d85f222d819ef7880076ce55fffce48d2595aea67e6c42dfad07402c1af132863e08e509b3f7984479a3788fcde3b05130af2fd9a85b67b4f3e4bc7109b055b1e319f874ddad882e9d8d93c44432a08cce430bf3e12c0bdbc5e1626d288ddcd20157fb14439ac79fb4f24117ba6f9bebedf793d1beed88fda21df5c582042646ae84ee2aa1aeea603de0af4a10bad05b85f0db42b454b6bc32fc9294ebae0d2274d81c4ffbdedfd60a9454cf2db96cfcf4d9a762ff1622d2936cf66e0717981fdbc1e2f5b143986d9989102f9e5871f0b9a1e99ca4dff9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9ec4b6e59e51143d37f228239e7c8821af5ba066ebe137243e6a433aab4b4d3012921cf2aaf2e160592ae51098a9f27b6bc9855d416009d408d50ac62f3c4156f6e2cabfb8f0c5ab817a9ac9738809fc28b53675cd3bcc4ef6e2e473b40e875580fb1b67c38368ed379be4d0eabe6e9a66038e12fae70b5b13375fcbf1f617af497a4e0c918062627483edcdedccad27a4639137ec0df4dda21e32033a1d2606cca166821f08a4dde15112132f55881fd122b057008f74accc66c9e48f84269efa9b40fd976654b83c416470e0f317a23cec78fc74db045c22cbe6b4ad9874b8916e8950629d301989d4abea69dedc896948710180a2c6d4cd7b9c32039d2d99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf55c6c0946b67c74be956f93064f1cce562194188e2f173331bfaad94b9f63e1c2ee295c8abbacbbc47a06220fb9fd401b57157d99a5b516c0e5c16c3c11f5546a82a5448d3a866c59511617369760440e24885f146964607b8350209b5f8b479c563bfa399a80a3912ebb095e0bd010bf9cdea9028fc55c828f33f2c9eb2495f16541ff944442c8bdd4e49991b2565cfb611e931cc09efd0f2ff82ca84fbf2e0843ece16132b79a59005053c4824766b1e3366ec5535469a33f288a8e07b28d4c65ada3103d6754aee18eb315757c61455f85620022625523cd0df7e5049b8e15f678ca0ace43cb8db30343baba35cca24b20c8cc4a381e493dd91f5b489652;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h41a8c94968e783125d821b797269a6afe1cf29375ffddf7fcee621663ef68c4d37fbd76361dad0f9bec9b0fa7c25c18c32a88a0a2e8b1bab0546159f3c3256fe8d4c861ae3689f250f736d5f3c8a66db0dfeef8d8b8cb2bf6a2278d42aede65e139d761dcc0a8c5e2613a85156984bb1507b55db57a711f62fdabb74449639925a8d04eed2fe0896c252bfa21e66a950b20c5b837d54978cc76774012e2609f04cb10176cbc81419127442b9ec3ead5a76f35d391879ee27bee78465e13fe8bb04fe4dceada50fb6d1f6a9d0ad0cbaceb185e0af22d498b8ac485fddfdd14bf3cbceeaddfcd118a7b65cf1d9ba19f91c26295ed60ff1766cb241b19faeda7d58;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4dec58e534b5a3671bd47dbc93c11f9eb043d347398557c90700ce8cfdf60b4386b6da066ea20c6c74790840da0034c9b43d68ca2cfc8cf2eefc3b491159468822d5df5438078b13b28dd88a66948dd498cfef3bdb36d9230e6b6f90fdfae9808becd8f82e6e2f61041534d12a9086522bfee1ebf8d48238a1bdba91c0ea87c25f3137001979467c90aa984d5625babcd69057f8432fbc085eb04f692e7c0d5a5a1ad401dda31ab35b750652210dfe1c94f03ad7c19d8741c6809a8eb262a4bbb16c6075cb435ada31b0690ad90ad65cb5656b1a55c2aac7eea8dba26ff8e154c91814005273362047ae10f5fcc7d240b078e93a35fa1f7465bbc0d10c995cf6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f3919c1ef4546b1bbfdb6d586086e4ded683df086a61815d69cc2f9e290815a39157c219ac0aa6db9ffe3b6c60de7264bc1bfc53860c1276f7f0f6925900da55e60adead5064bf1182478a88735099f1220c94988feeccd4735f122869ace165dd041eca4c710d40378384998929d117e80920169cbe841827d95b7ccf5d4da3e309b74eec5d220c75e07089c80b04a1b81eb305d302eeed7d789c5484c8c77ea7ad58b386405b539db870739b972911b16d8ff35ab8e372a5feee9c5485f840dd153e77eb36edee719c4797784d06ee979a7536049f6ed44af0589f2d98ef1970346ab31b3bbc924655d7d5840579ae899880bbdd7a1f4fb964bb0865c4a21;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfc7ee6513f2b3471e3cdf96fa2be7714fcd2e11ce6ab61bd21048399d841b93ed6975c606e951903027521006925143f241f2a7752b928ad30b073743729950c64c4fd232caba2f0f8007091d715597167b5a25b51bfb6e0f45bf8b60998bb46f14cee9ce2661a7ffb1bbaaefdd59661b84d99ddb9b1c4305a4336fb31ae078dde51d92a2bd5c80dc4883a63ca9705b30bb70e07efb0bfeef6c8400967f0fada8110409219d571f1e5e4262af66d99df1285483796476a5f3e0612a3555223899fedfbf0dd1e6e6204d9429c905fa634f5575627f8dd2ac488b2fdfd82acc4fa31b3a46c934e0831491babc6186d938b1046ed27ef41cf0c2703e3aacb9d23d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h88e7457624ffd886d9b8b1751984ee113755f2b4cf3b025ef009fd5747725616c36bec8dac091e428772c30a434338dea8a69e22cf86fa3c35e9fc8d166b95b6241b6d2ebba26ffc6341b0ae301f66bceb4b9d056d04a3ad80e5e1330d4d4a8d009c2350210fbdb8910f3e2372654a699f452237724fbb3db2b23892d7a0176cfc0213d21c626d530054dbb6265db0967a71e2737a7ab2d1aace6e732db26c3e2af99027a101817fe5a643a3c1042c2ff7515be9654e8ecc7f6b9a27ed56b3450660ab7de2b710a61014a8cd2d4bea953862e8d1219dc18d39f5182d5ca3a25b15cbfa7841473d07060972cc7027f0e20e1a50a55c5ff9b6250231d88c820bae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6a2348dbd8b08e8e8f4657660be6091f61277ba30a9024f6ff7ffb45f3cb59d83e2a7d9a56a8813ed430cba802fad60b9688d570f91b5930b09777eed552fc9a79e8763535fcbce3e8753bb3504522dc1e138a4d73eb50f9e3cf2b67a3ad7b2fc47a9f02e4bc8bf83d4ddc710bd393352f5093fe871ef757fd9ff01e786403c6d62b207fb6168c2c06d4d7230578568626d250c389a3224a27a2ba7d2b2b972511a956537778dfa13d5a2a6fdac705f119329ee0b2d4fa82d809cf9d4ed3fc1eeb0d896856f5db15fa74c501bbe64c6285090af1bfe44544564718555a57e810cc34fc0e394af6f620d019db824b69ca33c396e9f5a4c35a436502fcbf467975;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf24e595cb380ee86e68192e48adec5912cb305e4b9485b19730f023efa85ccfbae450e8db6d0f1e59a59fdbd033cb25866f8237051408bde0c3620bad2a2978a7c8cfa0a4a4e077336827bc21ab5685f8b587154f06732f58579fd77c5f2df6f999b19ee1cdf82fd0d8e7c747f124f4a93dc45eeaa129fe7ad0f89dff3a270997f897f97b8492d2088fd43c642ce8f9bfc0cd4e6ee39c0081e5ce7add8ac2aed13dd57d7a848d360e00da8f08b7d5dc9ed39e6148cacca500c89ca5952d37bc8e4569441e12846cedaeab96e5527da196db5d6e2d4cddded62c09ce9f8daff9d1afdf488d6a481795836c3db330dfe0e129f1905baff61ddb24651203e1483f1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3e38b903b2cb1a3b00961cb92b5d004acd180e981709a98195717d0adfa6e103679b17b00444b04f5b1ffe9af72e61adb13d39750c6fd985b56230dcde21d09695ed2e17c051a27789a0e050ea7bcb6f86429b13518095b3006c6efd2d8a068cf5732ab94042224bd457fb6f34fd1dd417f4a0f63384de9a5a42fcc0bedd7978416cc9cc6c73799013c01a65668e6b11df5d39caeb21847928be0b0bde0a7782dec2cde425b3b35878723d60e87a23b77d2af0f026b7fcac0fd47cf50247163dfe69219e7bb3b942eaa46feb0db72d1cc1d28baadf129a83ee39f96d1102feab53bd767ebb3f4cc6ce680e52e3907126c9407212051c2e0db3c206e9cf453873;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd0d16a95963d3e167214070de8fef878ac019b9ba15eb6b1e1627f719307b2a953cb83cf68342987154e69e6ae5cd1747aa3e430bfbcd78bc4d2e837a61f71671b3946b63496e9ae281b206212323540c85a16e382c7bd28b1f6764ae1a557c33b3c604e85bc6d15435119da8d7ddeabafb2e3f1b61c24d731a9b59faed4cf623baaeee6aa34236dedcea17e864cea9d2d7052ce45118d4d35fed8d76b1d30ebb98b5c723d4b191f100004255d2fba019006ff2d120caee127d5b7d7aed6f917f4d2802601a01c943b33514107b1308930f4b571f8600ee7b6d2648653dd7c6d361c160813ff4cd6007c599fc205acc86a18f96d25120073bef8428aa42d17;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6cbb60f1e04a60e78c9c229457bafea895ba26ba0cc9f63338c71fcbd6b614105d2ef9bbd9e93976147b12a4c26139f272b69ce1ebb538bb8f5586a056769697305195547193610813ffc1fe5b204380eba4cbfa1f9198682364d5ea2b39acfdb118d8ca470c4704eb133ed1d3bf04454eeb7fcd89c09f16142dc5cbbb0bf00f24629c3c8de83bb5e8bce0a739ab4668a62f498bce048ea123296c9c3d2884d09124de0faa6a947ade6aeaf5d87c4f17153707a3cc8d876a166bd96cf8dae822d2ee53a1ac103ac7b89a33416c1d39b09843f2acb23c0b74b2d7d0bf8421b8c679cd489bbeb19ad650d8bf89a2c41aa45fd57245d4aa4a098034929f03a124f6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea30ff91bdba0f9cf08772a1565f3bdafe6c4f5a0f55a18d70b4785f000506daa60ebf91068ff18bb3bc9e862e9d0813838002dddf2f220e8ca9507a44823f9247662d760c035aac38d45c36b00e8269c24c0f33b2a971411df1f99ab1b6855f6316da06b5354d16c6f9d218136e4ae7ef88280907007ab551e86a0b859bd8cbce1286584fe1de5cd59e520ddf0502f455a30bbfbc95f9e25e256899d7798628669ace12e10f0a555d1a13c96979284f9d7ea495e2dfe1bb489a3010da3eaa70fec8c6c3607c5093138f5c63dd2f1c278d6117156f44aa46762ab858e3d4ddee23bca19f5f7a96803b4f9804f25f617e116965c34580ae8e73199afd5e8b98d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb423b05ab8107842359fe50aa0fb511ec73d02b078bba933a55681b2826b2e42598036ca07138d6cb6599a9ff5675f6903789eecc21d5cef5c6086cf6bbdf55d87adae24baf8723bd9569d191d77879184a6f9afa037121cbacd581b2c4b96010ce05cb88268666695a6aecb898f6531714ceb44838ee2fb2f8572c47dd7c771f942a193af6125c75fdc389fe6b32de79320b8b10dab246fac48db81b3343f15b8565a74dc318de201a60184362617ff63365e23ddd9e932fadcba0572800f6f907a5a007976c44616b70de046c45bf4c226fdd0920cc49803abe3379235c5ebb16e28e66852f2b1b6567e541acf840ff7c2e70ae9192646e049125e2433eba8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h91f5d59843297f84194a75794a600e5013f2791d46e52bec7a29c505d87a3763be1ed924b1eca91cb5319199db2de75ce2483e892d45e9f6aef40387d39bf03a43e98be356583ccff24f7f7a4ffd88dad99bd5633ffd35d41221ce24d9e1e7afe11ac4909122bee7f6103a9efde181b8a2da8dc8a8cd4126f68a850d672521d639687d01b6c16f04d563862ab23a5bfd11143385a3bdea1edbcb48cb6912d19ae1910c92f18b54a226acbeb4637338f133e01723fd40bcd4a3bd66134cef69ffcdcb5190a8d6b3e5c97b37183a2e9932689418bcb34d39438a00bcd702a02f7c9353ae5b8f73afd01b12160e671231469d047bcde024daf939d252c1556531ed;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he957ce36bffb7e48def315f638a5f6f66eafc6d9f6607c924419ff566c445dac2e192ecba91253d003cbf182bbf617ed65f62b9a3c8864b7fec8869fe0ff8320aa45f7200f9a30aebdb228574eff94d201378a5d875c31572107541610b002402fd8cbde0c849d8ec0e208216d90417164d1b91e04f90ff266ab50aea293f955f18733e5276a0c4294df17e7715324075497cf6b783384b09997c0058fdba95fa2edbd6d4c894a7b10a85501d23314f9ade0c810481796de3fcd97f0dcddd60d6a487088caaa7ea3b32f2f025d5ddab1a50a88c454188400f2456326cc0ca71da86afcfe5a93ef5b3aa3bf68ea1feb46777ebeb8d38edcd9d95d2c8afe05372e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h15a951f3fd7206de2bc9d22088141217ec637ee69af7815c5ca29a1bf703c105f7626577913b7c52dcf8271b952101edd439192bade49dcc0ef9140a804bcaa07af88fb82c667695218839a7cb62fc230c0d92d176ad1739e341ab8b86bf35eb5aacdd4e6f908afd8ef170013be57ed7d0a91a8e85625b05c59140c33b3afd85c6c7ff81659ae18e0c9aba9421e100b31ca5e625417aa1ed41d84a740e59014fb366ab2ae5e6df30e2141be4c5c1a908e8138aba3616388b3ce6e0f9f1fee772b14b3b82ca1aa6934118b7f1ce0eff670d0d5caf6082f687408e8e471968515afde10c885be32071c1dc801552c79d7ac1e25e31ee64f2e53fe560817be9940e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4ddbcbf791b357532e3fc5035d76d59f7ca43cc60792294918c3ef0b606e2bd33cbe891f6125631a3eb9d11430887e298e6bbca116eecbd39e017aa2a3b5edc0b88f1b8a5ed1c3dd08738895a3d005749cfb8166c86dd106b0c2ec959f7828e536756bb661969274ac31784282da1ab85d5cb899ee1c7d0a53276410d3a7a2610bca2d5216c9576368279e3b31d1449b0a4dba582c94a20c6600d851be5bed169fa94606665b4906941f1b9c4fe633d1b6d91f7f794497056c6ed7b96e3ba0a885de6691e5ac09fa09fc760b98d4b0c262e39aeab5bc13bbdb3fb613c20b7d4eb456a00ea8e3fa8db0c690c095544c6294c072f8ee935b56a0d45b8c0eb758f6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h705ce65237faf3ac8aab8bf86d318651eddbe890aec5a7ec34c98e0be0e306b85ef76027fe5847024068d9afa8cf315f2a1d3fcd0f4926ffe4dc0fcceb0bc924e468b37165dc40d280ba11298887bdbb2d0b987667dd938abdc0afde1ca82459ed29a5932023c0e25738701d9fa7e142c3b36406e5083d488002bbe8c6b58a6f12bcc04bfd37869dcce704aa53dcdb21adbe3de44cbb7598fbd017af50c3b9f9a2cf157316fbe891b282ce6d01c1b26e73b10afe7cfe297e3eaa9559fa50ca7a7c721d4bed0375a5d0d6787db677b02fd4e6ac2af93e990eba4fc93a36c44fad45cb7212401905fc70dc6f9a938903da52e839293a3de11106ef60db25053239;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h103e6dba0887409ff005ca81cabefe204df140b1c2b420d2d796ad1964e2fb7a4558eac4aa18233d621aafec4984dfe8923a102d94dfabff0a00cb2e54a940c40da13e6557c3478b849e91d4cbc663008a0d4d7ddbc73ce4d296bb3f4d8ac69f7f08b1c38f6c4c344031f1f0fb1c9de392edbc3e3bcb082b6ed8c0b64eb6243af1da7f114eae363074d4dfa1ffdab33cabfb3d0e22f9a6295165d9f05b14bb0dfc13a735d9f3422fbbc0ca74c3efd04c896798f9a78f2dfe157751d16b183797940cb86e739e1622cd5c81ce3dbcb27f99dca2616157205a5635798f2e00f95a9030ad4013d15c7e1e497d01c215712e633c1bd637b15b0482e5aa7540dce3ba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9d201df87a8e3c60df4d7b8bc0b1d7d8a75091cdc0adf25874f08ee05e560d68c1359ee09f13ede206e0b01a549be3f192ab76306e41359e629144e21dd911b94db3fd684b892b4b872d4f9127e25c0378a9ec1886ef1cf19883e15d0da3e6458281aebbb71abf68ca9e2794570465dd11b5f0d4d0beee03e7520e88fd8e95d0157da46b193c8af975cabf8467d04d701fff20b9c2bb675d9fb7ea703c0b5c1a642cbe032abdfbc2dc00191c5e758093e9d913997bc5231409ac869a953f413d0a6a48e4c706ec89bf402dfe5364cb652553455f032147918b44b5bca7bf74a4a2dd3b9034c0ff47c9c21dc70eac0db058f20be265a6cc379fdde0b392f63e76;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1554ab26093960085382bc8cf5c1c64d7dfadf3f413b08f4d27ba9f2b2da8481abbdfb533d962166ef7df61f6c37c0bd95817e70132a771df6ecb999069c73a120ecad43a7c077d7def99b30df3c2909f66dfd8998430aa51da253bdda7135452471d3c2a7fba44de354ece90786bbebaf0e346bf6c320e483a9e495f5aa3a5e8d9ce6c344a87208caae085b27c060a1ce91bf72e10a6431e54f36ab93681f64c5325a90493ccad65698cb4dcbb49ba9fb5f5baf2bca7ee3ad93a691a7f0179998cd9a3465f6ade1d353a9e34f4e68eceba71b0fe9cf57cedc8ef07ffe5483bb8e5bc18ce13d96cb275f6a1482d8f65fed8c000d89a05d9c5c7655b97c74711b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h50a8f69616aea8f49addb35051ef84647a0f51a4abc52deacf76623c43c85d59cc90809d3a2f976a9138ae6fc005a741acc7241ed1f41bd2337a9fbf08be1caf5dee61a981dceb817785b300296b44a67bcbc62e35c175fd9e27c86e1be520f58d3756318786ada750cdb4014069036382fa615569d72e5c8a36f7d80468d70c156673883835eaef188fff3d42dd62fe5fac52736264722e3e1066e72899894705e461e69b0d1704b77e9bd60fc5885813aa1a11812ebf6e26b5164b7acf50dd9c3d1c14df627ecc03f83dee5cb495475dda96ae443447890bf4d12433710d57405b5688e04aa66054eb602b9c8e391018f7f027da49c60e1a337dde2fda27c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hce91af62d595db46545b0edd59f535e3f1c5cc088d1d95d2fe503eaf7ef48f46d3b53934fa639369dbaf756d5d0299d11e9c645b67b83963ce4bb88400cf022e694977951340161a1368029e14f9e32e8ce9bb12bf85aa176b5973d0c52a1d0c75f57bcade73c5139bf30f0f358843aaf3e40b040a3f4fb9c3670b251afa1901a745f887558574151c750cbde74888c978bd09c69fae0c1fe27773d3050ec44736f84a44c4e024c505be875191fbabe329b129d7b83c0c3edad583a314d355cc133509c69348ef10758d40d1ad83ed11302e6e5801a95b9403905540b8852e77c77e5c210f962914fedadefcd031d842e646948b6a32ae32a55d0e9f39735c9f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4475029d1b4793833f88d3ba2b2203a0c423a79a5cbd8370c499f5ccf3ab8a96cb427baed24d9bebfce406782bdc6036d89a39c5557688cfc37d4808b1a42db5f4daccba11b0ade98167acfe4ad3cefc89971d5173db023ab713bd098a2d1297bc4da3885ea45cdbe7bab56e89280d217250eb2fb8f16c8ca0f108dd1ed3868400b41fa2a22157c890595a0be8af596a93b6ddf516b8307c7aaefb98cba41a860366ebf02802f5217aa2f7713e62dc78d5d3a701b5967c2f243657713506fc7da5c242d8f9b9be6b27e1d3069cc2bfaaf58c33d1545819a54c6f3ecd486d9b40828220b30646bfac1dfe001ef544bb0ccb8dd7858208cebdba248ae796f49103;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h49e6c3099b252a31274c20582559c0ef73a550ed823e068a70dc8cae9238efa0311c0e1a795c471d01e6c9104eba6bca39943c6533967307e226bcbc69b365acc7cd366129e7c184254d2825e29e012acab60201d22131b0343c21f2cd9462cf14280011100dfe38fcce92663e72ffb5d452c19c8e5170ccdf1062808abae9cb19a974056065b2c8505154ef483aa5ed35783afd4de2b12a24bb358175bb470aa94be607e2957aa04c07bffc2fb14a98c6cdb48288d1332e5ec12795bb1dd5d43306b6b21cac789a4d1462f067c48e92fe5006bddf0e3d81621fff4a0090ba37bd161ab09ff9508767ec85b3729c88f005b86f4cc9b19aa0320ff59f201854f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h74240def954b0bb2e787e90ea100eef4b4d2f97a49ed556782c364cb025899ffbb8fcea3d2c2270c21cd93b999ba3ed19b94e1cbf59d46062112b6c7f292d4332b2810a08bb03b9fcf2df143ea1ed24941672f444bb327598622f9da3a5ae2e6b6c540c2c5cf57d386767a0db0727ee2748b109b7bcf32328b0d409cc92630ea435773780a680dc0b29fa55b532af6c94615442693b19bd6530a0c35b2ecd5b8b1c0d9dc51acd17ae922e00813a486fba38b302c31d2cda78073fc7622f4778ea7dd3b623cab347aa8a1c4d5b2f4c53140eec8b34425d6735cad6715fea47ddb2c77cbef5d612b1859036a9813648e309b00cf65c763745c902466356de789b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1dd922532aa37c97ce5118feb45b1b6a3f820b7d0b412913a5001bb84228340c14d4b3eabd620bd3eaaeea558f30d0a0b3854a54fa6c2504b568652810db62c2d21fce96e0bb80f06251a83880c4e6e29fbbf544b5a858af134a9c2806aa9b2c62d06313bc219e31d9368632ec25f9b81ad88f255958a2ac406bcfa1992db9bd5ac2e0132a9683537dd308118a6c487bede5eb58b8d72f06ee5fa70c7550fd15663a7dbb332febd095c0ae53eaf7bb3547fdfaa768ba9fbdd1daf69c55f60fcf990b6ef7efc86071dbd87cb2f1cdbf3bd4ba64d25693c208f13d9ccb69f80cac224a7bbadbc55596d79c224e90e5558ed80a9ef2741b26ee96263699e9ec8894;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h318388cbfb693f2dd58f9866cdb680caddaa665c7e72cf18189149422ed5cdbba555143415faec331e564b443e51621156c5dbb4ed7366736764086a0cd95691d7ded9bb2fa29405977a1e8db477fb841b6f7aba9ca4ec901a0b1204d384d12ee8f20a75726c3ba6aca6d822de8df04341e46a9fff850e89ba118cdfeb52b724c4402bfb9f370ac521006c1e3ef3cde88a907f2ac6a908ae8fc41c628116cc725ceb689d97e9829db8e0f75dda502210e5453718e58a7f4c5388e7c57b2974a3d9176d9c1e21eab92ef36f311915454b953f7dbad008d4bca5286c3374c0c7710f281cb2402dea6b27db33f9ff491ec643890079b300e6e7d547b35b5ebeef0c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5ca8f9e66e01150a01103b67cd3173ef0eaa10bb6adba13ce278da10288b0e04727329794224239294201a289229f0267fedd3eb5570594324c42ab6979a9ff0c661fcdacd2e4bd1803cdab4f0efa3443335a15452f4c6ed2de55c0da09350f3ffbec3733cfb99b6c375376a42b2918747014a6cf0a28a458a1d8d3cdbba618df65b39f6d7d057f9cc2f9d7e79665d5e0891d5f9614de9fd4cb25d0c539822f05777405ff02de4240e8ca22fb79ab6ec010c556aecf7271d2fa1683653605a354610b789fdb9eb65856a9561fb0b2895ee32a1b7c5f1d56fbcaceafdf53d7f820506e00099e3f083f49adbdb5b118819b2d9963932791db6d5de86f3b77bb919;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfcaeffb9d85b9d13a9c697d21a0b9604592569fdaff39fdb818cd3a44b3ac5b85bbcb5d8718e425ce0d0c0fbb0deabdcafd441ab7619c12964cbe3e18d06d291b41b3e945fbffe5d4e957b6742b988d9861531d20749b8f520a02525e62db8849d09ea1d9a07fc13ffbbcea26ac9659ea27d286c8ebd6682f56c2643a425cf8506dd3bbd04a06278192c1099e84d96cff83e41b2c652d470e23757998af4d4e62059ba156fb5380cd25f1e8a93409d24b13d96857a6bd4a04a8c7c91752508def23ec843076b5c5080d7e64bb040a3b47e06d201336bbb4228bb36b6c56d5c804633659998051b3c0c9eef025ba6130fff1f064f3969ec317e7e613ce26f401c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2d596a5598c41eba8caac3eb13c8025db7fa92f8694bd4f4b31821ff6de0c7b489635541c62b9f1fa9f52c85a17e0b730562ddddc2b81a93f63b37cf2cfb963fe5314635ccb6e68e55d255ff7cf3a0e14fafb7e58a5595ceda1b86938f8602e982e7426007179d20b8547f6b2d5bf5620f1c79d9a80b055c0f492e06ae0b540b0e682ae7257a446386e4d3c806d75a88b3fe371d7644b252da546c8430ed4e90fb75fe638a68260fc3952f45498d202be191f02a3d7589acb55bef1c8559e464cbdb5d7e3ed7b19e1b3317fb7644479b401d5532b7c53081b61633cc1d29f6c80b2f65cda57dc89a2c6f9726df01b183a97675157d0890fb9163015f67d25866;
        #1
        $finish();
    end
endmodule
