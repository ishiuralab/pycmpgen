module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [22:0] src24;
    reg [21:0] src25;
    reg [20:0] src26;
    reg [19:0] src27;
    reg [18:0] src28;
    reg [17:0] src29;
    reg [16:0] src30;
    reg [15:0] src31;
    reg [14:0] src32;
    reg [13:0] src33;
    reg [12:0] src34;
    reg [11:0] src35;
    reg [10:0] src36;
    reg [9:0] src37;
    reg [8:0] src38;
    reg [7:0] src39;
    reg [6:0] src40;
    reg [5:0] src41;
    reg [4:0] src42;
    reg [3:0] src43;
    reg [2:0] src44;
    reg [1:0] src45;
    reg [0:0] src46;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [47:0] srcsum;
    wire [47:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3])<<43) + ((src44[0] + src44[1] + src44[2])<<44) + ((src45[0] + src45[1])<<45) + ((src46[0])<<46);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fd8821a6a3a51f6d53e316a4c21f4cd4dce8678dccaac95c068fd71df20a73de4e4312e74e87685938d7a1ec7be5db507c2b329ed5c411187e16494668c87a35c1febe847b5279;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h852f381efa375d9479962da19adf3891f1ba1e5bf04c0461c4c86eea132f9719d53d0b90de762ba90590d244ce9171927ae48a73094652c1441d03a703aacc2adb93e705bb519cf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89b14300f74fe77d79e37af15fe5f92e6e425a282fa957baf887ecf37a4e725dbed24032981e3f58cde83c65b806fa3560675a45373af0ebb49efce882c76bdc0d341511afd69d9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h151d6657e867fb8c191de17106916f7da8c006a3ac99e70622d3d9c38d94c39abedabcdf6cf77e2274f2d03dad8b1c9bda97166c65ab825d7b3f598747895565f0a576a1e3f35ee0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h895dd6ba84b000679113eee73e0f9e76c2fe4ce5d077e61aebdd725831e0ed2554a269a0a577ad4aca8875ed79b7c45efcdd52f8083bd197ed2216ab6d70ebea4258e49ad2f22841;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1a9ec32378469f444f2892af76ffb4e57c80e9227137448fc03fb1a7049f32991e1b174168eb282551d5d2967605d33d1fc7f000271500775fd8dd23c832f5fa015da577362080f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89f01f9a47f361bcd0268927cd4ed0a8d8067870d75ffec270d6f7ced5ac7f051a32d0ac15f4426fc13e00d97d24d4e0b712a583109607753e25dd6f6f6f43be845273a8da9e36ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19783ad290628a29fbba002ee78cc7ae34ad3c61f5a2ab7cc01b8a987c9e40b5e38b076c2ea4e42e1d7babf0833364ebfa484ab441cb23f6cd30d86f2fcce66f34d3cab3480b6c0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe70776f0f8b443e7d3b9372cf89824714c179c10a6d5cf164cbd06fc62a1993c5ca62396010298d74bc71a45f2cfe8ec518fa8aba061696c6f6851705f9bb14634f5fa6f8446a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h870dc411275ae2e630260baa9e9a1a1b1a942c6f820f9ebf222655acb239e486e3bcffd79da886248978e0185fb8e4a4224ad8df5b1dc73d59fd1a89af4a654bc6d49996d32c422b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h493d18db6a39058ca741002a174ceb0660a9e45402a7991bd4c0097e2365b349160bc9ba566310435ca79dc9e8c64866a45392c3cc46b16707f87c62bf63c8cd522a2eaf02835678;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc5a907d1a8148469130d879ffe5a80a14749cdd9393e10474459a9f10cee1a417c8a11750d8b4df2186b55ace4d17eb64a87d0cbb633a2ec48409ae3eff8c064ec9a63d53c1d394;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h892caa166d262da718283a517dc68309fdc49147cba2b163172645081cb661c1d31e2b2048a55ee998d61221f6eecd801fe8f7b3ed343112a06f9b5be42372fea071c0f82fe9fed2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a43d41744c783ddbdbd10d63cd696b61ff5188abf9df656e6fa171c830a2d13bb0f1631c51b700ca735b943f851b6ae15b5932111f8476e984553fc2f79a4f83b1d28a8edbd9681;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eb72829e3bebe8d05a0390e4c833110244065a16ef70811bf44d69ebadc961e0324c9fcc98606cd6bc6709c838e9e9a527425e809ec0762f16ca7822a732258e20c9f1bb1950a5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75e430bf8d9ad89a5a8e6beef3cc621cf292f8f3a39402aa37e20e6f398ad5d43aee2fa0cbdcf576fb7d113441a4ba0f98de8a9b1ffed4a86de5eb132ae0aad59868126653d3b09f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4846a16282c2192fb083e470c29d50421442c9383e19cc4e93736597b46c919c21ffdec236d1dfdb1de5c8c5acf3e4de79a083de4597ea42ac776b9bb60e14a3c9fdd8bff16667f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab5593891e88a406e3db36d69c2db8b5b05e22b1c0a0d8c65611114f9afd8249a22386f9a5d20d50bd9ebeb734a13242b73f8255db278d0300659c2cb8512a5e9560920842063ecf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8c35a0dd909d305f5aa091d0e3158fe7d50effb33497496f7d413e828a2be630d735e672f54eea338448dc1980a9989f2e86b3db8ba44c239e4a53ffe3fa72eb20904a5fdc5b1b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccd933d3c650f5897abbc84a4ffbfc7a9d1c6c97f543e9a6133dad8f7b028bbab829a89097290b8522b66f861b80caf7a57f5c0d56b8c8d0a7dd86cc27581071f1888b48dcda82c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83c4e63ea648c46e73488d177c8f1fa4d33e536061adc51f8c03b33a724f017217ec5d9a8625c6bdace68cfe8fe8fd607d17c9300bd5722058b23dc24e1a8997125f268755c64ada;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20e9018f52cac015999a6bd25ac81cc89f2c1876742ca82679e19b3804036a54572efd63383ae81da2bd99f9a57321f935438a871a0ce7e3c21dc86996b96163676a8e02ab2401db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec449c83d563d56f6def7b5247aa094ff5581fa636211ec21ed6adee23fb7e50b8fc023a7b20fef388e3c9f64d4f97cfb7e58940b2a190c0d437192892d7620e4d204fe8fd844e81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e41e17c08a5b9537576b5d2e3a5631bbc579f3c358643b86f29ac42a69a4b3f05ded3197bd78f3816015df8dd5bf1fc1b1b16fdfd8fa76ac08e3d3d537e0817beb55825dabaec9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd41c5935c69d323c4c363e042b5c6d2fd4155ca579869e94f2c38e8eff24e30a6e0a71d22edc85c042ad82c6941ce6bfcd5d1cf2eb59e319dabc74a067324cc90a1f12e75681c2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7dc690fe7bd1a01298603afca9b354022357d3c5f4eb7646cc7dcbfb0f46690a0e344eb5857f66edb08ea29a137f2d47d9fde4af6a17178a3deb9a3ada2e9c7b1b3cefc9d3c68dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f75ccb04786cb268c0e97455a74bb23cd36b3ccb28c142b4ac196778b191ec47a6aa99a5a8829e6d1df8d599609cea7afe2fa0f4c2e2626a7da49b8c5b86cee3698f61e65f5537a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb65a2e3b90683defa227b181bdee3e7337daf7fc62b1bb5fedc3af8055bf2b78e43d2f30926058a346fa29a3d563b5caa6ec4908fbdd42c95adf5a79d4b02f1dc8da99fe9e892223;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56430aa248aa64071465154ffb61925880d1d4d354f7801c41324ba2af2f27db36b7d138a2d8590b43ecec8d1d5d7dce5124ca01ac67e44b210a5e93a4577a5d6eb9b167ddb82abb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddc4d33a80434f477269275f32840ddfe808956ce1beec1fd7d9eaa24a2e24608c4c86a34863d991e40ade538f27314349afaf3653853544fa217cf9e846b42b32b7043ee387cd04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae5e4aa57efba31c31e3d8f9a4347aeb170cfe7b5296bec47ccf6cdef098e9843c265b66725b6ea107f49f97153231b5fe7fc66061510b0b09466728b1282dbf24909dc77be4e083;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1353450fea707e5f61e65c4ad80b9ed8450968b6e23634c3cf730921fa77ae7b4e2167917bce6802896f8e98d000b6a08744759bbc3f9d88ad6256b339babe5279bc26dace8edf07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbd34469911a5855d3ed82790f62bbe5cb089c2175d82a6f90a3b2a3c8555693c0db0dbf07fc3931cd66bc1131ca1fcdf7f4063d9dfa0d9bb3ced42900e4b008655b47e909d5efa4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9662cdc4c4cfa82be68d608edc4ce36a17934de7ee233f190d989092f993698be41d122573f8b5baa2c8b39701507bc35424cf6988790c73133bf712a7e342bde4acb045fcce253b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68f074e6772a171d59196f1815681a1d04eb0b8a0df7193bbfb673dfd4af7d92da78a5cc8a2587ea69a571b60a0b9b2b6a7d9ff0ef8d24e802a69cf7278c1ee27d27220aa272b49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he37a4430af9e143d3aba1898c7fe9453047df037f9a8e024b3e4ce6a8a1d58d9e0e6de70ab73b13d93964a0629aa13c4068a79028cf8bd1b655f91be8d4d5fecbc5182341debd1ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e998b9728dcf693835b94337eab0099dfc97e060cc30ae831165c690c57aa5ff86a796ecb64cfe1ebe92b6ef451ee647e185e090322556ca6a294ec1e836ae609a17a8db18d2495;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6032e332d8884a27a0965920dab5e328b25655214d07a3d9c0f4cbf1b5433a006b81428c9684380a5587f789f1be51dbf9e1b0601488a9cf5f700736b61993b1f0b8ad7d85430949;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e324071c4ff63f19a0fb0b323fefd8629e73dfde5731682a2a9d656c9aa2ce7e3190cfe1296dd9e61a4899f20511b7b4ae0870c8f0c8dfbcb09b5ad273abe694a201dfe25423d93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2b17d854e43c420818c3d3b8203ebcebb685d4d4c2f85bf4519d93c203e1a78bcf502c5166b484bb615405c314541c47e3ba520aa0b4e78855cd850b81e435ff85a56600eecf2b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3120c5358fb85f0141666cca6f1971bfa799aaa2e965052d476552ffb644ccb410443acb5361ed5620bfee9fd3ce11f6b9d179c8b43a795447897f9dd2937a909cf64536a589fec5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f0e1e9442f1642011b03a4821f0b824a530a489cc46d30fcb2d70b00fe4bdc3fb4cd7997c1e64379cdadce45db04d308f5b3e6f48c8c856502ed4b8d08d15b549309f787fb8c194;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h243bcd643ffbe4ad37ecff1d5ecae0399aae6ef1534d3cdd8121c91dd0145204a25c4242ae95fef0aaf9c16db18f74403d6a11780400488c53fd5415f31dc8e4c08c67c4440133cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf89515f9688ff853aa6026c9ca111ce50d361ae0ff7302812c16d33ba356908f7bdde4cf1bda1996a3875b18a6670fe5aa24bd16687708afe68030dc9e16a18656742d73a9033b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7a90c08cead240901bd9901202a146ca359dd35dcbf84a7d055cf0f179312e23959888b6d48d726420ba9b730ed6cd16cab897859eb382f19957cec6d07c47eb528ae79ad71fda7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he71a6e666b6db75a95d64a5c9fc2896291ababe6e59fab511208d0b033a19b0c75ab3e9aa200918a5723f269d158b3bbd61b0b4d51f120bc0b2627254aff2db14583c7e53bd38e77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h423e16f045a05b8bb3faf867af6ac6908c14b9babd4f6d49fd1bd0d0d243bd8986cfa8d5502841a570044eae5c2ac4c9c426bc0667c9894dc5cade7e784cacaa71a73f46094352db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1df336ab2b4e07fda07c0ba24f91238476bfe2bdb35f15c00f8ef931b8d811121486da01aa5d5639d7e52e9d20772ec46fc41ccf36ff7f8dbf46b79238167181ff8311bd209c122f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1f187a4ba76d91d644ba6ab12b0ba7e9fe777e4a3df8bdfd599a45158edc080e7ae2eda5305eb1582a93639f900e46eda0bdcc4dc0d791fb1a232a1cd6b93894ffdfe0b0441286f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h379617a501910c709416c3524baf6851ff9470608de571ea77ebce35a6b864ec1a45fa6823ac1df2b10c329397ba5dfefd40b9f7c178d6d21b1158ecd462e4a4d44a79988bda7923;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51b57e536d3e239cb3cdec73a7c18488d1fc2b12ed8b55a6ce12e756e992ae6729f4593c2b19ed3fc94487e8bdc5d8ca8f1e4d3cfdd1b7900e6c4c1975a905e562e8b9180b546d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h355ec5add70c5888945765114c044c0bb9da70ec5ad6c0ade76ea142e90e37f1bcb025a48555fdfe0ffb0d32b500af2a25c737a278a365e85a91a0cf6c2cb3a52c9527e06e30ea98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habbdf9cb948984df8b8891db34f15d178a9b8765d7beb5ef851bc328338803278ce5f0efef21f8b72e80e19648be35f38c64b1dabfa47f47d346006751970c96898cd8680a42d45f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2623e7a76b33a4698198f2a0c73b32b9bbe8fbcc07f8e1ae260abc1e81c57121a1cb93c5540ee32687bb84ef0b571350f7337b6aab7bbebc242367072936c9d492c8983a5f5ba3f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27323aa7ca146bf535c7b6047a51975c3f4674d1f4bfd59cc05d39123eb9d196351d808821bb4473ea393c9946815edcfe3941e16b4da2fb6c72f611f3e340c2a674516c8b381ca2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94d16cf0c9b5a862ebb6e5e209412219dbc06dbbba61a5974aa6c3228d1a02eace76a3633feb22d1bac97145a55439cc06de27771779b5af9ba812a323a87a14cc00184c3d32a4f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a7a36b76be155c1a7153f666c3c9bd983a8ecb320fb0cf9d9644b5e675fd32f8efe70ea6a916efdb58c577a0a7cca76be25e8b931157fbb42c2cf65352d5ea273541abe6835baab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h265587f0b26caf08a125e4f0cc752200d44e7cc6f1a36b55abfb9077249962340a659dfeca5023f85555eb705e83e4447f75c6a56108c28f1ae85c05853066383e52d1b98845e6b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac8a8140c7ad043ed1c028c3c8b77e1f81d4a3ba2f9306b57a7ba89c89bcec57a0cf884eb4ac57e73802b9ffeaf0c85822721b3815bf0f2bf911fa2bdfd0b423e48c8de3b141e012;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e39ee3e6e5f0bdd7fad9fe8f0c733c288d6dbf77f649ecf0f4fa3704e2048582fdbbf42d72e1bfba7b15e238c2640014a46233ea7cb25f74b51279fae2ec1556041dc1834e3f476;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1e88239a3d41ea44242277acc6a964459aee9f0cd0474f976233bd7e8bf7f3a7d460baadba9661e70afc2a22294d3fcfb9ddac096791ad814fbf8836ddddbc24c4677709d5a1767;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd15d1018e14df328fd6f44df721022487ca832fc276936090fd8292e64e367872b340ab86ddc8f5bd5a98d761612e1119007d26cbab0e3b8e01eda70a088d5dc643c37c9eafd9e1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82300b500b340299c1728543b00086e68289b9f8781f0137cbd9e816c71651ec931929b94cfa34263a5299714bfd7fdfc39777810e621eb6b8d5c046ef140a9826c5e625df0de4c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h200882e389f9962c62d0e6b10d0e4d421bfab3d5d17625893409b546028e97d6657ab40440a66fed5a440573ab870ed36e796e4664e9a70103179129862eb4d13096d9d4350750aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96900a8778ab61c5050fe37da4296701938b8711dd6d1145f56b74384928af1e04e3e0715895c2f56a7a73c81f9c84156e1f034c9b25bf03c73e2141cff639adefb2af6b39e63eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1238d0bc0d3bd398ba849104eb21056f18fe0f40b42a2bc8b52ff3a10c3339b55baf13b95782a6858f597b53723ab439daed37860ba7990f76f913c1f6e83560b800f222d6668b64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef543c812da37d4cea60cc69797c3521d44d5de805363b85245636cd76a3f3bd4be5ee6ef73a565e94bc239190d014cd61f556bd92ce383bbab50ecc559a27dbe53f27279d4321ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ee7fae6dcc9c7fd34445c95031ec1b7042008f02b034a7c522495d170a2d4b864694ebdc580b81f9c15de6faf2b23e0c4bb9ea92a8457112fd7bdef4c9887f697ce54ddc0314313;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc17b09c0050f28066305d1504c8251b1de54d890fa225187f035028e2361f733e5e65fadfd8388bb0b07d483528a03fe3bc586d1d14664b4a7d257f9037a427d1820cd056f30e7ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b9233175c524907055c3fbac36e732a2fe1e56ba6b31139c719c0872b31325db50b3816490dff1953da8385023c908610b8bc77de130b6ad44926fb6d6a391131c315c2d1ba3501;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc58c79e1b680845f3858a2301451e70996fb7679b81b1256f92d865976f5cb4d862380f90619f789b8f76500219b781d73bd8bcc90ffd25bec1b648629d92cbbe678386afcf7ec35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35d2b56aa04bfcdeb12c63ce681b0675a2720e6f5b3b148dbe52d2bf47a7b5c8acd75fa1d4a37beaf72a3a3b43b4d45facf6046afb4ecb6dddb10d3e80336366e674b3fc3208ef72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbecb5b8f29e4a072823654ae848055ef47ab935be1d06f9aa91dfbafd4adffcbca51d7e6259150ae4dbd7bfe1698f4598a4cc0010771659e6cdf017d3db074a0fc3411c0dc42718b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he71a8ffa93c0b24b4bad5c11ff57a47f242038518062974ba6ff70960f0c5ab127c26c720f6c9e2b19984f110dc208ef41bc6a5cab1b679f551e2e85aba7665875f2564b19b6b271;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc6f5f438280f36f273e8f1d61f72fcc09b55a5b4a30d3535919b21ce7c019c5cfbf28207408f9309e85b8aaa70ec9d5149d4c3dd43a860650b5a59f80a4d35cbcd62d794c2753e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb2f1f1a265b8b4ccd809bd2dbf71e79f4e855f02d0c3590cda034a8513608c23da94651c0c036f310723442825793a601e2f34bf606012746052e74e1167e17f9eeac8c73cbac2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48428726a5bf8e57f48812915bb0b9d79ab504d951a04cd4184c80a1023fe672a3f559f831d4b6c66145d0ceebaa39448e3c97d8932d22e4c9ed61ecb6078c7bea9cc1877a3e1e6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9e32445933bdc00f9c7c4295bd2b832e29c600d0bc83277e9a84293b804194cf96593905713c35c04e1873aa57bba509457e5f923addc420ebac2877aed471fda46a7996477a024;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b99b4f990c5a4b51e2eb24c0b16eb882331dc6f04543eb3031f5a45d103326186075155f2f26ca0a59995ff2ae9c723a8464e4c2a915cd04eeebf3e9d0e919fcf6003a1985ba10d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36cef0613be406775f932ce540dbb62174a8827162cdc288a35546e1393e47f4f1912f0d0c913e72d2050a43106646d05be54121843d12385951e3be569024b683d68146dcd2a610;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc52cf51f5e39b0dc48dafa89cde9f3a27333cabcfc5fe078fb85d9cb509bce0898475580aff11c6b35bd92105eb51a24763ff4a6d5dd2b496f98ea23edf3101b9e627bcc6f818d08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb35e349a43551813360faf5a5394c3c9c69f7fba022f60e332d2f1bcffc43b6bd80186b983db8f65d595e4537652699f424c7589700d1a8ba099b9825a48a5b5fa75951140ee36bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2419017528c6cc2fe70bc9e32d94fbbdb66c239b2074e2c62da79932388ed30406df25dac7118ac68f4a752eb2f8239fc7bdaf6b2a81d8c43baf28f2e58bf1f86102e70bdd53d3d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfff094fee3ea8c622824df830889fe00f85ec350d3a7370033ef98c66c6564a90bf7bf17388fd0c153e015c34214967f7e92b8cc4f31e321a59a5f0bdc715bbbfd615eea4de06de4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3ec00400c71c105283bff2c146554513f08458b42146710efdccf679bae3e1d48ea3d4191c2f4e29e1c9d5983ddb51b35f02baff49c75f39cd0b5e93ad43ed287f0ad5d14ceddbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h177f5ea7c8a5df64248117ac78005dcf0d34002e12742bca2d98a77ebbaa7e7046aeb446363e161f36c3fe967bcbd56a3ff4788c60e3650dce3635316f69d9803a23229317b760f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeaefba79e11808b2f56276fb89822f9bbcbebb9432d218a29574032e3e24772ac9dee8dc7d51766ae15315180733bb0cbb7f91ee343d3a0b0ea81ef4826e02256ce6f7f40edc439;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b31da6c53d2b4b52dc4c1409470fee7a9364c40785491e6fbac13549e539e370696c5da1e7553fd1f927c329340ae60f33da62c61b8f381c10c157eb5289f73409efe3623a3c281;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb639a6d5b5bff673ef8c0f39ed2015b607a41049f1421878179e0dbbffaef41f5fe8ad8c9892e670cb5c6d80fa30f2e88036edb49eb97cb0dfc8e4578367876f021c54e6c69af1da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f50a0855a512084279ce2711d831f98b53eab171e15958ecba7c733bd9e18aad6ef3951a184a2949345b8a701db50488af4e9795657cd2543a9402ac30f05222719f57c60aff475;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h562e74372a3a9a57871755c45a2eaddaf78217aaddd18885066c70de329dfe4fefc2b293f1998cffa626b8b9db5efb9acf1635cc8de1ac4c71e7d426a517467583f9217bc1a9f90b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cddee3fb756deae046f24bc0c3bf4163efa0c8e4a9ad62c9e4e1e913897b223d548223b4fef7729a18fd1e0644da322ccbe88f1b2f97735d3e1cca22ff3baebc8f56f833b0a606f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85196b2e704bbf1f09de6779738f70d3bc2b26a3d14dcdc203e90159fa0a2860d6040018ec69fe3b910f1ffa581083ece9b3691ea191e31ec24d3af3bbb7b6ce8bd42a6e33ce9d7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd992969552fc8c6151858d78cfd1d56c45c3556722ce3fcc28dd980329f5add98494a418371bba0cf9dab475fcf669b74b69fa073988ea74a8a54b0824f42417b04132066b5353c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h471ad77e7a9aae2896142750b5f119f57178432752508fc9ea83fa91fd765582e934f28475cc935658be891b9ab708e2faab1e415b91cf072a99c8195ab044d016c26e70cb25d286;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3cd9f7381e395030527c13f7cc52acacf56c3113a51fa5e4057d17daadee983caaeed06047d5a1ed13a9a261ceb6b4bbf3fad781ea5644045496bdd3d643996d0f61e07a4a2097a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8bf37f49f80dd4018a63c392de68640ebf4e42af6a0d13a0fa565796a7066186a2699f17c6f29a7de8ccffa4893feca02a59c2c5c2fd6db3dca387efd0eb3545fdc68700d9e3fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5dcebbdc49e99cb8e65679b69f91b82aa00a8573af9c5b6a7079d13b6445932675509ac3f0425b8f4fc006732a8e383a36fbdb5c96dcc15fbb4be9c54857ff273b974b04caca494;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h252f52175a588b0f84c169d1bc1ff1c5a119244400cec62df30a9fd7a021723c7a221264331be1c08169ff2d72c41f833894cdd8e0b8ebb7497a0078da69161e6a6c2010f85dc4c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80c301d4a6a8ea558ecd400f5da0ea3cf8025c21677ab8ed7fc8f6262aaebb4d2a3d425487bc779a39fafed1db846d03210e6b7133d537a851ef60e4062c8d83be8bce5ff3158cd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25b56cc349b7da88f3ca08038ce13ffe36981291e9b459f7411111e243b50b794e572dddc4cf8e6ef834645b9c19f84853497aff209520f22b4ef4436708fb5dd81e2454985c0da4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce8a014fc77274d138ec8b7ddfe57dc8ff2249375088253e980b4fea6bdc978446cb03303f574701bcbd7bd61cee3b98ef5f3bf6c943d06ec4429784afbbb65b56ee6df6b80db25b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31e0186e37925b93c426261fb97f881991a7a2f9a8559d92a59ed3092ed47bb37fa34e929f252a37a3c19b28213197bf0c31d91206cbcb776d909f5bdc7bcb95318280f0367df04c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0d669b3b9ac28244feab2c375c6bf07ba570e6f713792c5369c266125feebcf888d3b3d99d5206c493fae10a3b98017425d0fdaadba7e28c2013f348288f099e18d0518f277f791;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82555babc7bcd35971a7825e7444f26f0cc65f724199f937e5866dc227c63a96b6ce3cdefa7d7dab6f12918327be952d5bfb10b72f30dd53c1a37e8af8a5c9db76d7a65c7b45b4ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34f56a80ab80f47c82ccb9ae7d156a64c02109cd4ea2937321f4943c413c13ee9c2c50a16638009ffcbac16c64bba933a77d589fa28634a2a2c13b06e65e1d829d7f1d4b902bea2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadd813318f4e43e9a3b5af8a76fc78b4ec3b5a3a0a4e0dd74434276c93799ecf6cfdb997810817cbc7362263e9a1f490a798b0dd766d306ac1e0a7d1af6ddbef56ead15708499c29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfe3f9a1b054f4a74386f91a4a6d9dcd4e1d04ac0658fac1737850fdc379e04f26a1cc37e61da7a0a3fae1677291b7865baac9a21ec5a88577b5580a312c220f07610286b21e9d51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96c7c7708a8dd5d28315d6d5ee32b5995fdd374e2142b33b836998b1768d33042de486443bb640f46574a88e09bd7fab24e3d45c55ab926646c8852daa07797ecdb7302771d6d45a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h178e51d082dcc34b1ed35b1e69abe5bfeff979210dec6bb7483bf063e6202218407275a5db08a8e1490f6dd692a29513afd766c44de83f5bb92094b16136f219e41335254bb04f3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c255b6524402f918dc615cfb3e5f5c95bb6cd527ce8abea03088ec42a7ea90bdc4d41fe8ca747b24d9be58acebb9453efd61a18c37b9a12982099c26cbf4c46b154bcbe6872752e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d5bede7f0a9cb3e20ecc2093ea6d8dbb182ed86b1ba6f64598f29794e07fdfdfc0a0ec311557184ff1cba873d2946b5134ee36e98e2c7c6135afc8555293301c88c5630d214a2b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he19caf13711619bcc6d71cb27ba6892035e9e116fe427e5aa0a6aed95b8cc4b42a9d5091ec8fe6194c9f8fca2f6ef073a03aa6aa6f2b2507aed7b9830e38a3554dab659c4c37a60d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h606dc2467e9b09bb77874ab394999d2114db105c6b9db7af938ea6ff56e5283d25a8030aa831f0a06d336942aa7e2f8e5417523416ddd16064efec2ee953b244d6c92f303feda602;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6142a4ff4990216867855b03e7e27341d4b3f3e9a093b059ffd75461e627205aa2394e8f7b1ac1ccbc1542009181797853a2d93d62ad80d6d192905aa85f1cbc3806e0a40732ffb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5ebf5732a1745fac4acef5b0fa84f9eaa628f292259efd488d2e8d9edfc26fea3eb2a49bab03efbd338f4918f2d0fdf8a45f31a0b6189bc9787de1c0ba63eea1ef276b96e7cbc03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h575502fed37a2afa49289ee204c2608d0309d9c41d869f18a1605ae25263c68f521291af1f042ca22408a16df89427f9a9262475d44d50dd551909b69cb58e760e80fc99269fb09a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he28e1e233cb2f9f884eda467f14ada37d2da28d8c62bdba471ebae449f60d7b66611e832e919f538a0f8f456965379b0ffd00c28e171222dd58939260d6c81bc3fcb4fa787763c8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12e3d299a1c7f1a8271d6edacc5c56f45967932c88442e1cc59a8232118beef669e127c1a2516bfb4a4fe48ca21d7ca841588ce1395d16ed9cc325aca15903965b305eea19368e7b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69971a3af5d36977b7e1ac54fe4cdc6176bddb67850161ce790ab0593e4ab957bf90e0a796a27676b0e49e057910258376c8fb6fae02e2d1488c48a5f062555cc1074c05b8ce6779;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h149785cecc2bd3cb640f93044a5313bf80a057cedebc6bc61b3684aa0dbab0e580e7245cc2a3b38c3d64fd903eca0ca20ff70e4e6057a4821aa33242372cad3370b9ce4f59f4aff1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae3913d02d9266d614e53349eaffeec351335183ce0a92eda78cd250774b3378e39f1acbf9f2ac23863ed7ff95e74606d2bc4c5c61cab712838cb7b3825f5e0cbb5763ca3a931c10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcac331329cf8203a6450585379a137e95faca401d3ced250c0319227a4e17234da530938273d63ed664be02db04045e24339c3877b52e5a02907b61ee89b492b0c83ad724c75bef4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h132a1dc8ab819d7b65d2dba82fb7ef308b0d860992896f1db38fc0c8051cbe34a8f5eba2601dfe2a56d3e0187bdd7f3bfd200a65f6869f3692cdb26f8b4c0f4ba2f21d310adeef28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b2f4fd2e84986f9c94e9051550a8f179b60deeb86c1e8dcccb406ddbb919bbac52d4efa2bea6f9a7b3d93afb14fe1edb06767a908f6346f30f1a20b10df1cabba89658d4d0dcc5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3b01740b03d57faea40a786bbb6839956f834306b40cc1ecc41b3eb3a9ee17a43cf446f69511e6b8fbc077519e374760aa2dc63ef21c8d146295eec3ea037390a9d92f15e105d4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h734c5fd775be1d9e1ef2fa039c59ed6fab4ad377aaf25a8e1fc4a977738fdc6d4dd63af089712ea41dfe217c6171ac2c431cc332d1ecb02438c71a56eef04b83758877d19f5f1dbf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h199cfc6f27bc2d218cde6d29ac37c1dceb71e387d37c0a1748154c4360b31e5cfc7116ca0fe472387498cb77b9e0f28374a6b62f46afad0e088215c7632fe953274f6dd9d1f35381;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c3b1aa1a3c935195e0281fa5b4e70a97dcbc1a8d533bbdeffa33ed4753dda429a971dede13da204d4d4e8c837f0b048ee865de51d81652a011f9872660a72b8eee298a44c075552;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ba0dcaa6a44104f5179121b9c3fb56fabeff2ed1bff868e6193dbca9f3a8ea1db71c051d4293c15e3f3753a5683b0b9b095bf2e1327943dfef201034b01787d9851eb3fefe34592;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77bfee81165d3b6e4b295b8dc7bf6153e1ef7b65f3df4ec894081e5a8f83bde2139af927b57bf676196374b053eebb0713390b3f20e613628604b71a9d881977fa98f795cd2c47fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf82d60d2f3188718c355acf64ab0044bf8ded9b4845abf3607577f35e01e2ec5cfc4111e546daa782ec570f0bf694313a10a808524a48c33ec8c60ae13138665a5d250419a04bfab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebe593c5966840709c8e0946b3815f35a89e3014b74d0b2eb587a2f6abe5d1559c18679fe402f7402939f1b0d893eb107a3d1e86364fcf0ec8f066670daaafee5c010a035ddbdb50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91c54222f82771e5a180df69948574a9e0ae8da24e402ed920dc67ef25150d0d3b3ae7441acf4a95a806c7ab2b31c7f91d214edc6e04f29237992ec5a392b545ef5a2733971ff626;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1902db61f39d9388f0f4e81ea2432391cbcd8c3c9d4e19a9a5c74320e952d33def936bd3aec3068cd9c801836fc9df0aac1a2dc02d7ee589efbce5c894612decc5179066120e7c14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd46c378e031548fc722829e0d9400b768741ebc9fa31020946758a4378014f8d1856dd52af2f38987227879f442975f304c170444a43a7db6f78e2bd253e862b59d0b47c83f3231f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc35c1d12567cafb8a6fd58447686bd99cc6ba63107ac398d6136dd7f278129906f72f828b266aebb01e553d3ba46e2dd4ed51c57717cf8715dbd2ad09a3fbe6b1332697d88809d2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e13a90e1321044214f7bfb76267611e705adddb39a37612dc968d1784f53306d11358bdc2c0dd31c53aafc3256db1855ff6f5d4e3e081c7c65d94b8fa43bea1866335fd6a3f614c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64a230a3a2ce862caa8b9462b4c0c866bfbddec446d66d58f2ed4a12633078be4850ad5b3f5642ab36745363a3b4257f342832254871437c438af038c86becd57db0bfbc79db739;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h438b815c847e252dbb3f4407578a9d5c674f6f8428f38810d1e86cbd53b5c151ffe52d24d458aba312d44f05f4ad40232689fd92017cf117dcf4773e03d6395ebc958afe36ea79a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe43a80c83a5a1baf7b2f2ca74939d363e2679e4e5f00589212bf1316ecaa4500c46e112184d40e8a4d97c324eb5948da7140015f3c423d1907cebdc0506d1ea3cfbc9c634ff73d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f8836ecf03b7ab4c1284818cb6a865bca1bbdb0a4eaecc1a8c74b2cfe9159f5905339b4e1a8e9ccffe192b30f3a557a89c9624078a5bd2638adbf9082fa5ef45c1083aa525afc93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1ec38aafc76106d0f69fa6589b3fe6170f3070943903467f7034c2eb559b0315293d9bcad922895247887db4c91c139b027bb64f7400c5a32d71a9e2ca50985a2647b8b6b5f1c28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc143d0124143e099f7287532429fe9681c5ff9f4a3070d0cd42be63a3e4033396b05534ac9aff3e794ec3d3b2a98ed9f130a8e769e8e01d8701e407302d4edd892e583a4ad1d49d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cdc3672706fe0bdf911d6b4d94e9dacd82c395cf4ff959e798452c0471d548d5b6ad9e25040bd608f872bf1c85eeb8387f248b16b35416e7ebdf0b27c4bd4cbea69c2fb75f1a8ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45bd5cfc08bdcff59938df2a682c53b5fa916140d0d049ac285b1b444d6d0f0c7e6b6b5c3c51f7f046b308b7d3cf9793032b099ec2ff53d6e192c6350f148fb316b398d234d03f66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h249419f4ad6b153a29131ce56ba1abb67782ed58684937774495409d6dd855590aa923d069e6794b399c7a28d0e6e5476d0163ecac3ce1edf2e5abe4a5eadfb6cc8268638682fbb9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h149e75188abed7f55342f805d925f3cfd3ed60e46ce108d8dd84e944ef5903669435112b777f0042c033bc3949a923ad87682160141d5bd16fed09b7c4dde16fc09506f88dfcef94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h742ca652ab58d4b1f3098b5997416f71cd449a91956faffb43c86f7b9e06febd67f897c0431df605bd6898d0b2c29afc446e36fbdc655bd21a4d80f2f742f104eda7b098c4f3e4af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3dffc153042d8c28fc344ad57f7d2fb160da64d0cdb55948ee80ab56a63aab1ec45f317efed412ad5e75920d897a14cdffd348eeb8ea1132767838a1e5fe578113439fc43f64e88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha202f5c3250882ea1ad78bbb9d8b3476bdb3d1d50a0b15203376e4b5b3049cf24755b3167419dd6d43fdf37afaf473871dd699846f753468ca9deb522fe60865c1d77a779c1eefce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf53133934da7b9c63feb7d9ccc67f99a7bb07d5bdd46a05083c00f3c9e29485a4760d9acd367fed0fb261469c431da4cfccf8afe989ea21ab5b84ce025687b0a9e2da5976e595fd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5e97ed8ceef100eab5b81dd25a306bb2d517ae7162349f28890dfe6db74c9d092f7e81aace96dae0acb7eb7d8b69631c76f65ab8e301356d9349d3c42a5a15e9fb095f11873b643;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h731df18822883fc3ccb51c791e4fcf2acf1d531e6e842a705e989d046ac9d14bce72d2e1ca25a6401498df0952da06572cbd9c0aa53844876d34906e098e0c611ffb0144e69b25ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52672a5fba221b33c898a62f75afc764119e1c95f239473d870c9778c61cc7a95a3e7e71a929cfd07aa7af97ccc4f0f08df71f86c14eb9027a2ac5f1a40912453b4e15c84f70a33d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6e1a5ce24941eebea3a46e64a2a19014a74881d181dc636ac73d1f4b1c55ed99e8fe0eecaf4ef881df8c502b237b64a8e4e6b769c32fab0049e0a9d411f5a3432256dcd89a72f50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7863d79e4e0448ef71b888092df05b7f8dea4a1a7d099816f1417eb332297f55399cb0c1aad026565830cbef30fa1a5b6ff85230d63f5c5fded762d3f81a9caf8ad367a1fe446e1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9602e2d524343095ae8ce4ecdd83e7b82451940eb35a3139ab776013b28cfeaf1a6bd5ae1bea2b4c57f23361827bf227b360ed2c44ff3643727eba2c006f11a85a125d115c2f5773;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c474870b85b696b458d62977e4e6fbe1c4969a7db9cc37e5b766689f276b1fdaacb8812a4e00ec2953bad743cc06a24c9a1cb24a30b2dc70e89b75025799117f1d60666a214448f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2226608b535fe7ac9b10e10c30ada7776b1b6e0745af68b9048c81ca3ba97cd873113dd52fe9603e495a77b1148f4625430f82c3e53a6f4149aca5f13a505e7f41b54bc232a65022;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha833780d9e01593d919b2d9509f5b452125eb64c3dcfa095a7681a0c6d94c7ee0bd852a1a6f069b2ff22f6225b8b8ee64993fd7576f6cbf29bb4f6429d30f387ad242a7a26bbb9a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf13c8b8526becb006ac55539ec921d023377bc838258673ab8453b1fec1b1ab8c2c68bd205a0ae465ae57ac11d43100b88fb362ccecb70a2707bf8b4aa0fa91c547a5eabe1fb133;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac930220c1f86b3981e020f0b55ee4baeb67f83300c1d10823f679d37e012a2e44b45616e72fec07ee03f28b86b081ea975fc8d524231c55c105bbdf4d6401e44f223e04e6f520bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ee8f1e39dfcc5f5a89a87a8f0012106fe695725be8b97aded524b4b881b385c3a933adc5cbe2a04fe4811e03f360a42056552f2107fae806c3eb999337ac8f1d586ef8d456fa54b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2a5ff7741c42271ebbc34de63117535067946f3b151d08cdeac32c9cc0f0a0866154217c0121d21f09612bf574df34b5714fb32fc15d672a48cc46ba859c21d33fc9055b421deef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67a5180ab60baddc9ede6ec486fa8a20718a21bbe9370679be0443886266b85af1c7c6d1919ae62479b8e23f2b030b3e8792ab44b2e42c875c12241231f6897d643f0f6033471cd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b4af1d56e0df45082b414e55b73e6bb2d8d89d3074be6a90767e706d81e1bfe878ea27847ab08e2723f08cf4f7982eef11435dc9f5ea37f56de78fdbdf307893ddf346cbefdd2b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h963c19664c02e480a103f790482d0f90d308c407978bcb96ae6b700b4684d6cc9507bbabee5bb0f45de9b05aebf9e993cb5286faef8ff28eed5e46110c7e35df8d4a889f8e67476a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54988a64d9f0139580cd55ced388080c6b3694c62ce8c00e2372ac1e911fb0e86bac535e59a77a92fc6b597984312befec3fe27305d1fc7b430238cd68b8e159291546177b4f8908;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h312a1d58c3e009001a8a463d429e9f9d550c1aff017b6c66118430601b139f8c19011d9d4784ea7bffb44c8c0c7761e8149221405cccb65065404e1aaeb51b735a94ea270af331eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ca6c8199bcf0362087d19bcabb76b348a5e20b2edb7cf2c5ff8a8fd1b0073c3ce42356aca31f7fe3dfa4114c27d2a0ce40e31c0f173b1ee8d7cba7a94d7d8670599b00ccf2fb4a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha42770f720fc14636ef51b2012e73bb390a8b1a9a2acf9e93807738ae4221c5f4e0030d25adb33e7113d07b6782d73da558a8ec7a39e63fe2a28b63daba2df61c2c178819717efcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb1d35a14b12e89b8845c5a36b05e832d388b5d9a1f589fb188848b275aabf668df5015636bfca3fd41b57e81538a04be0e6abdeaaffcf1d17ff6e4275d74ab0a38ed4a0b75b61f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76477095d164f2b0e13f1983ad6f7c5166b83bf1ff05ace77a93c979ed542d6704a562acd80ff79856ae325d5a58d9b764ea64b667f5e7317e900c2d523588e66146d8f0f4878819;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda1bfb67f25eec739057e3de4498da1f93b9393eb5f6480fe40bc033077b4c0aaa7cc778cee14e78bff086e572fde919cdd4340d4cb8ef23e428a8cd9f8da68d8fb84d747403f68d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h263aa7a58a952d06e1b154df287ae72e9eb398e3555fe22b1253b512b9b19960ee4adfdddd1f90565979a841907bc8e0b635275c1c43d2d9c0ac38555d89fe2b2de92727891f4bc8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6396cf1aa47d7c5e6081d730e88b462bed0c0d0c822fbb86fdd161d17e703a83ba29433978d62f57144ee1d394d3b5599b03c1569b75c636d539b0970693acf9bc38f7cdb581fe4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83f5a92e42d24e76003263a6f80b3444376771f511dd5dbd956cdf41d62e77f14a1fed263831327b18cd7953dae8c906ef499f4a9a18c2f1c02b48de19826d9bbae064c348a4d363;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e3101b9d0bb1f4c791e5a1d8859ca99a7b7032f016854ce7ecb33044dbdb8f9c55e0cbec976562570b7cdf95a77e19b0bcea7ef36d3eff20105af8b011c43cc618c22f61426219c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70c3cc80f9d49b1da42623f4ed4fe532a23330c825afda328cf1dda68decc50e2aee2e4d0891d0b0aa62bed0980c40a521a40a3ac313aa8d20f3bae8bafd2f8e1d5200e441d4e319;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h704024397619378522419c1c78eb085b7a4f2472b40ea5f08de05f1ed03ca46dc796a56281b2253f8f5b67fec323fc962851fa1f37b89be5d4a6f487c9c4232561178022ae560784;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89aa0ad083d12815ef2b982f3f3beddb0218971a08cb4d591c2c4de04678b8ad5e6e2f51875df6421bc13bd50360250c9e33273bff2e2291d34592254a6b29f1e6b4ac684ea3c6cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb46f5ea27b3fde1d55ea498203489df220291df26fc43535c6a572cea89b657b341e3e8b2b6aac12b2bdcaddaca45991670182f4367de2249da1fa66e83d87fd8847fbca382e00ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b62d7ac33f7c004d9b5b389d39a1f5eeb2ed991524fe9bede6874b9ab676b3be3a1d560c6d97210f1baad73c007af2af9283e852325814841798638a0ce02263726276abea3333e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69e16fa85df00e287752e54831fff0ffd23ce8679ade9f4e4cc7136010d90f6e37dd70605355bfccc1d178a9198181db2a018d45e4c40781b74d0db11a4b2449773bf846930be480;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb0a8cc65b7e30489f18492d627f0a5254bafdd41edbf82161680062351fe229a7a51e13271b31c8b8977e73456606c0277e04e1ee5c772627d687610da568a024ee8048f5870066;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce6f993544037599a99b5cfb543603802bbecff8bd6b06596334894801a4d873dd03b4845eba356e656f972bf9e860a6f4aaf5d116aa1e8f64fcc4cce6551fd6576e97b8867c641a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf930d00cce4f69c7a46ee5393bb709ea321dbdf78b3538df1f8e309b296f7068e0e7abb70cd7068da28c1b7efa21be0a862a98a710cd2ce6a2a0fab13de1f6a590fb048c0a56d62c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc84bff24bccf6e75c18afb01ea01bcf6e62612f1a05c637c30c17146853743a64eeee1f5afffa23b92df1d56a4cfaee1f9ef136a70c44b8a0f1bfcd9d8104da46d5d1da842968059;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h738b2a93d4b4ad9b1b13336adf7d18ed57a6848ceea580d9155d3afe0739e6f457120d538f0c99a90f9280113cfe10b5057e0e4fea1190217fbfdc69142f6541cadfd6e0053aeec7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5531aaff75422008654176112f36c20921bf047e53035e3a67156082026caf3517b118d39a0c238c3ab4b3296f052dd76d4ecab32cd46dadb8b0dd5cd66e59acaf09710f13a189f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1310400696ce6d9e271853a3f1f311df1f5df65c1a40ad25eb2158bc28beacb5db408e265e0a4b494fb35302c0c6f12adcad11d5bd647d17b65ef9a89f4b573f07e3ee979f919716;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d93425dd0b09de5f7737a84b8522fc36c595853350f4671653ffabd050a361ad9d3dcd6ae0a0eb22077d0bb0143a112e83da8edca1d40015598f627eb25ec5667e655fd463989f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h616a7dd21cc5e615740a241b8d9da4972a3e77fb8918b623770f52ac375e958e334e2e215cb32f989519975ee1e2b0ab588d67cc5e67c4cb4dfbeddee6c37710c22c9c3d6d11c661;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb68db8a4ad4ea3a1ea5d08b06d140a1ca431993300173419deb65feaa3d0142501af7db052e3d26ebca980b9e9b50221649e4a3774d8b6387786d42d4443e5b33872da97cd59fd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84d104fe97ec6a802fffa886de59dc075212d4f342dbe974180706af4a524c52f8bd1cd7757fb741b38855843ff8ce9a0490ecfad963f55ea9be2b80e6783eef8f424489cc4c4311;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c159e08054773a1a0f4026fc1842b3ff88b8c37d905753e0096d1fd3c882671cef154e5a24c46df4a39067b463b8ad47e73789007ade5bfa19bb22af32165fe1d2634fe6a0b7a47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e38376495600ccd80f5a02ab633ae6e85f4ac842c5de2e47a13839c75568aa66f97189e8dd994cad40f075ad53ac5eb85c3a6df421dcd0c16251f644a03a9f5589ea40d66ecc33e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha24b98ec578e3702aefc778980998ca924c27f227f06f3968d235f03f8715e0ae9b55d5c95390442e6d2d0278fec4b3c131a598f8b5f2e458cf8fab1040feeb34c7f712a4d64650e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4c1069861b6ba32cf9b31fa6fe30bb263785b765e6bb5133c33561ef59570331353d4e661a2723f781a283694c2d952b7608af0665f717b6a6946a5b60b1cb847dabff6ad1f7a95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27585953f09273cfd459950c08448eeb1fe7d2f6e82d8f3b03adb516d5069ee20d81922bbf185af7dbe05921f4a64f8e34705397ff619ddc39aa894f8b2c860911d411c9225717e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h136b44b5f4d17ced3908ceecfe591dbe7530ef900762b2004413e517c0c13ac9d2449839ca99c35d375ae92cc551c8173033b9750318be857c9ac6ab3e6160a1631a112597124420;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec92578b0e009bf6e1a7e3b62c7bacec3718504a995796e2cf1731b0c42eab8740d3b24d604de72197d6471f5579b5bf1f5c78f630fb4505d3489820f3e1e538ff4290b2317fa74c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96d9c1ca819e1f5271ce8ff25d0cd75ab9dd941b589d97db8a1df301759d4e9ee9b6d54410dd3ab921eb0ee7d6a5678f74e930f04836c75b87c33ffbf2e7274bbf750effc52a60f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60e981164ca233dc2ceaf2012f50273cb47332bc4925ff34533deb5d56c4be30f54174df3ddc57131e7ddc60c8aa3bf0b1490ec7e4a6251dbb52184158f91e0b118145490e3ccd44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4050740dc8e62968d7da459f4f5ef434d110503c3b17b6b56a5fbbe6bb0bcf3394808d91f32b099f8f501f4c21a8078e2cd6112925fb0a09a051a99582556793f34e431aeb54247a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6989f03b372e37119f97d500aa8414257d49efc39f04d8408fc510da03711ec9bb26ab986d57c4b9187a103a7f70801566e72882083ffd6a1cd172b48e51eae8cca070305a95ec9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee7c21b07fe4c3ed14401e635845e49c4e719bb43b2f5d996fd4d26eab18495990b3ca91107048c903f233a556acb9d3c2f18c0e97bfd6d31257117eb6a42ac706008ee6c0dc6704;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc75c619c5814eec69eafe6f77369b5ac4b10745fe9b7806a7f018e8e61d0d63e9b98144bf035cbd859038dbb06d3968c27f46e22d89faeffe0f14e5d89e9f3718c346402300883c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h492e62450ab5a81d2154b39a2c6f97fecf14672402f55f81d00d4f519d836867ac3ead70bd8ad7aa0c646e6c50cdec7ef0a6836bea5904eee6b7fd2541a849612fc54141d8429120;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99612245e2f70d31af8b5cb1f800552be7f2a890041fe0073923b79159453a467364d42bfad09f33a17bd4aef44261e125dcc17fbae3128298cab27f1335c9286e6a7b5325ad9188;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5df36d5d9758aeeebb65f5c3df9b12db32c4400ab5bb670419224c7af9d8be0e60184848c91bb7e5c5f1ee23736144fe150c9172d380d64d7d3dfc0d585fa3c8ea8be4dbae4faca3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51f6159dc22e94b17ddd31dbe407c38baa81affe3f590d0fbfe72cd40d3d496d70823282414697ad3a429242b4a6cc58e604b0633eaa05420721f5994a91d58a6e65e247a0195234;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d6d04da3c23d48ea64920696940dc8b64d6e7c80456e113e0f30e6dd223dffb8b30af2dc75a20373a628968534d1f55b1e4c3ae472d9ebaa00c19fe73667b070ff2dd68cb1c915d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h360a1cc61916b821ac69c432c6863fc95546818caf772d1a21bbd3fc5aefd98ba8d75ca2bd50b1ae602b6c8f67ebc0e781bc791cbef45bf6a1740399ea1ff1c1e055fcc90b50ef14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9488b2e69592f43eddda0d987de9bed638b82ce62726509c65bcc70605411aa20e42772201c31fa1581950251d7da6395e8f127ef516576c5dcdeef91d077265e6501121d17ece82;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbaff204c971cbcec605e090c2b79ab314e8f25619e7b52b57e1efdc4408d6c78fadff6f1f71bad3238b47d3027c058a020b37bfbb8e717f1aaca9a806f372f4846e02f601d2dd438;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfe308f57a87474e4743d0c3bf79ae29d630e25e45c98797ef00760996cb332f2b5756a4404a9f4db65c503906796e234a9218de3d94e074449d6285e6a61a4c13902f47b6a024e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd24a5ff3444561b62a03ce26b175a43f777454a8607f66d8e28ccd59a38e99457c30bcab9ecfd88a65f4f1ae10a871f6ca013f44cee8b4faaf895defc1fe5816f7b83bcf9c67116;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd04dd2c0746b1160b696edb4d36b4ba8cc5f7ad2be43e84b9ddf8ece709d2d93cafb99440fa0ec21f40552a8ef1bd02b866d06af2b9c3721b7e8da703231cfbfeee67f745fb69f4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12c53bafc8799b82cea3d0aa3687904ce26c75d3d3002e6d09343392141406485332631a107b39410d6d39ac19cec7d1dcb0d899f5a8ceeb403e8e18476db64d34f72eee55d2331e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7601afc0e4e0e86c25718b832131c44d9389d1835de8f71c060c35491f3871c4f1caf3988a16ac09090e4e4d8829a5f7ab6e7e52daf5db29224cc99aa4cd87f892a964ba9db6cdf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bb02488ea083fcbb51e70ca4a24063b36d0957cb7bbc1818b8bce60fa2ef961ef123cddc34c92066cf2c6145483299b5db20f8a9c17d5b702d21337e470e463b4be04d12ed3670f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf91e292ef4fd2e6b2b6d080551f3a37a71640ab6ba2e21ee795f8c3b77a85ff14b329f743d9b5b729f655854c1d2cd9d634212a925964137c96e2b472203c3b8324235852b38905b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fd8e0e62f3aebca67b9a85e1461802cfed95a5b5a407a4005fee7602fe361d5eb1f31c999350617f1fad57f5a33bcaf3b12e700e15841b869a0aec4bad14eae887fd5da511f59f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf63feff0efdcf674f3f6325c27a019c90e7cd405d0f5a5671b08dfe1e8a47c3858479d7a7ec9f5d83621b3b9efaa1fb903fb9e579cf37ca5b3332f0c1024579f6974c053101e06e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2774f399752479619cd67ea7c487b7612d7416f71fc8bc62c319e0c274444a32fb3e54560130045c0016e88d5e7fa7bf6d11f439fd7908ad9150b32432e22b2149fd9fd625834a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66ffc5b7a5f73d03e1070bec2e9cf27ac0964957a1a69e9bc3050cd5a2fd2124af3a7d975bd6cd1416936651c5906b0601b0fb13e162113dcb47c89c3841d6ce29da45d7cb6c4899;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91844ddaa56cf96675ddb981f4d60fcd71fe74dfa2585294e701cb4163e643164633db8a2549160e10ff3bd008a39253edfbd6f9be5614cb856bb3e174f66586b9920b24efad40ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h692ffce94e2f2a507844b6a66ad807cd5a63e705a9a48580607ee445906b7046f1ed74ed9ecbf506e22f7e1fd0846a7e88fd737ab1f68ddcefbec660e6eb62c38f0313d1e372e6e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f5c97826db412658e43824d92c2ebbda3af277dffab9c96da089c832dc7fe7efc8d2e8fb9af07d155bf55e2ef67bbcc092589d7341ee421b98c028cb7470958b8482361445ecaa4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4cb0d8db9671a835ff80fd2b7718e28b090cd29a0e2e883694ddd7bc1f984f4c03d03ace6dbe42ff195bae1ba7c18c283a83649cc0a2b940bb423fc7aa5ba9acdf570d3bf5ce0f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea7bf4340baabf4edaaaf63c427c7714e2d6208216976926f1d1be8539c03cf8363300b8ec7964c6c279c903483e936de6ecbd3eb788278746de50c1a08c6c3e9597397512936a78;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf0bd3437a4fae19fbbf583b46933b16a2e7240d783591d91bfc0240e1f9bd427da92a4d02e847313801a4323532c986a1cb4af3365b4800260feb570416239784eeab6409a2ca00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc31ccebd89d007b3461424a36a5ffd53cdab7b0d08a028b759256a825798132a811cb5f6c8b9016a2b26b3b4cb9835a031eeb6c8b0a5db005522a887cfa1128762dc89f4ecc438ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48651116cd3b0c59935d013ef9e1a1c22d79c063a465cad613d623060b66ddf4fe61c3a1b558196bbab76dd02d77483b78a4387f9ce52eabcec53009e6c6ba033aedddb6c86712db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9da62f0f26972187258633cd1b0bb2868031c4d457e56d6d3c2e503c1de97c2d3bad2775d04c90ce4622ae27f4743be6e1377409f0f8e8ad4d00f233d128d8d89cbe35d78df01a3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb686095f0c21fc37640c8e1e94bf0162dd6cb581229d32376aa5a0e9afa74ec3cb4ab1691fbe259f277c35458b6c649cd09ad218b3dad533c82a5555a60a15a3f4ca158d5f3fe55;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h824297497c7c23086b63d4a014b18f82649cd727bee8798aec0f2e25ac8f24e9bb8ed392bad3a9d514cc01468967aaf1ba0ec25912c9c494a735aef8218eb238d1c95af8b0531c95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4caf973bff0262f1ba27be4bb20e24c0cc67b50d8f32e805269d408cea5e145cd3d656db856b56538149c5e40a908231a2e2ab827daa5b38dacc21d90e6ca007498955b26f6b3e86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h218f3066902a110e1ec8623158b43a8331628b46cf47abfbd939a35d9d5fcf690cbebd1ca64cf9225eec91bbcbeb67b80abe4bacb8485979395057d09fbf1d4bbdf3aaa0d56a9f21;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7df0e4576b4216fc5a5b338e9b24fac25c2b4f76917a1eb670ad6bde2cade0765f00ce679deb08de0eeb0e5b2f307580aeb38959059d51ddb0eb6358e93c1a7ba01ccbaea8dfe2c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98a7183d4aacdce8e913ca8c21ebf098be2cb405594a08387be1237a32cd18017294e3952c8554202a7c9e35dc5ca10f144332835c72db32b4c0320c0a06b682a7681bd442af16dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8722e523100ae22ed6c31d4d29bc645cab2b304bca109a0ab656d336239bd19d7c64695b3f384bcb5704702b44f4bfdb751d39e04fc1a52c0323ccf56856d295a63707c3bbdb408;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4965f1c9ea33698bce740aae476806e98d60a5d7ed60585f0b17651b0dbb72a42c8018ca7abce987ae1ecd048ffae9a9e7b1d624c475062a285e43ad6645e3046fbe476f553c6d0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54821e503e81251a0204f01815411058abc2d7d6ca09c80210f7a4842b9750baa08d10b9d8ac50d3e28c97d8f2a282db8a09670c2396d4d642d51ee2e5c4aaddcdc84bdc1280db95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0cba331b77d0c8adccaff30d54ca2616aff7f19ddcad6d8e825ffabd34993104f8d8b393328a9327b6320eeeb58f4e8df3cee801be23a700667ea9536a3022ddd58d4248287b087;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed3ea1e09005750527655f4035bfd3d99c3ddaae06b19d0dd04c867ff7bd27ce8808b229b6019de73867689c9808eceedbf8c643c79c253e927b10fb062c968875a4d63909da4504;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6815fddbaba778f8d90d8f71b20c6b7920b24421e02fbf1eed1f83cb18644a0026bf839fea3fcc678733fa36992dba2ffd756de2009979a047a8d5189f87fa58f7ce4611b3e0af30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2250d64c92a962020a4866bedfd9023930f30269ab791030440bc8de21b777d6b971532a77596f515ba7f46a2dffa4fe708410fafc15880d3af9c0f19725841f1c8ac82d1b23ccc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fb298c27db084de2e586ca809d624587a8bfcdcc4629d444a4d9c7bde30ac426feefbdb4fb28f14a6fe7ecf79acb3851c558fde66ce2085475164743937094044e63371b1bf2213;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc95b6267c464253657d83673505446c8bf862d02bf4d56be7a4c6b38d1daca458d62f8dc95c3e4fec6ff4329483622845a5556617fca57f4ab053d7c69f49112224f145235a3acc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82cc39063cf6e478b1bcbffd2b8c924b77782f3ddb61769a72c2f11037cd1c786b4b32bc048a457115df467a62a366fe7152abb6870afced585bd92c81a07b73ecca68375ffad24b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c550818e02fe08d81b959a6cbece00e2bcb553ac9e91e04d2b2e150a50927c2aac29e5782c7f4689df0c0df2c4728058bf91d8f4d88584afea7c07f0aa62351603c75e1c9e76acb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1dff76ea52ff168fc1323490990bc0d7342c281fa2f5b5a13b58eb4eb527c9ae3ff6b88a2041b3e17622a24c551bf31f4b95c5617e43f970d3db832a3916db3abd24a06c12d59d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1b904d550ab0768dd0e4a41fba25cef38c36248b0ef874bd06104752296e9f3e082c6c0064daf6d1f5378276b96ea7dd4269d51e9410b744e30ad4d0b380f5a077e3f28ff6e05b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63687a4c877aa22190e54bd15dda5283ce065ed55b0840ff26eb93bc539d9d9bed1267fcfe03d0ba01797323e37f4552bb7a11f8883d81069520c96384e2ccd6c778b797d7c993ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8611ad39b99ea4128d421319baf653998d242d4cfa125fa2c96c46550a8e91978cc559b21bffdb698a467034a4d76d9569fa729f98bc1658dda5f384c8de3d5c77051d6cedf0ddab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2155acef647e928fd8bf22edf7b95e7977e0103076ff83be01f1bd9a8d987282b123e31b885db90fd451612091abc5e69600a09993212ab33b9188e50ce5eb9b506c898cabee7dc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1793c3a147fa8807df8f61400fd0065a4cfca9fad104181198cf4221d2eaf1d6b3dea3e816358cee32aed9607f857e82c7a8c58b40560d5ec19e4dde06fd43730a44227af89d64ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he86f8e6f835cf7cb38095396b303f7e66086433eb44844425f4f5da5f06cd4dd28893bce4232e89e14087b90edf95420b1b3a7d34029d4a6c65844a6847165dac43204d9667e3b8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5e5dd81ddc9c1ffabdf0bee350fd13aed1dedcd25fff6b6553934aa66a3ae15cdaed4900b093210a13cf60f62440a8364bd17c50d6be3116c3bd3b3bb77ccc773810e0c53adb916;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c7dd454c624f09c4277713be3128bbe414ff760b1400674b91e10510f57e3ac8ab99f0dc7ed0dceea74235ae00357cda7a07e5bd67e5c12afc995e7a6ced354c68f0e82247f722f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25b3020c65f1d9ba35dae39427bde7fd325a86f08930ca55372295ea0b0112dfaf3fa1eca77b1ec54743e9d4dd4a2d394f84a1bfbb1b66aec794a8b67bafc518c43d5a470e13cdb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb217ec18d31a680ca0dc6234aa3093b98ee9ccdcb4de9922ffe1ddf506c6a39af18a5a955925045af635afc01c55cbceda936fe5c2ed6f97c1111542c53ed4b7101ffaab9349fb9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he92d76b2ade809ded354075cdb81323c9ad05112265f56b8389b46f7b99a9824da7c28a024fb9e743bf0d887795268fec71da84957b71a3926208658364d1ab514085aa97398d700;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7913410fd0111322abe3a49a6d0af9af662969462032a58a97e78d353ecfb10b1971751745accbd6e9ca1dc98f10147755b07dc38d38e369b8a6a7f9a62a42e36fee19738dec2cab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9dcc4b631236e18b26d67676cbafcdb3551b6801d3b4139dd71975e4bb2547cbfd7e7980cfa0f4a20bc379ef203cf9b19af37182453cd3024e7f98a8f152a4ab0f18570aedcec05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d4c0bb9086b1aa61c9fcde84e0f05b245bc5d419111bc622b82f3fa551fd2f1013fd68925a84308e4028df938e8fec5c2ffb3f04bb17859c7dd3e0029d34d4b96107cb51b22891b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d6d70b0a36aa7309b902fbeb3f907f6cb79ca710eae3d6621c34465793d9816018d76b0aafd29a02551d0def324b3c8b9336f207e858540ae8bb4481b005c24dd47f1d86171e1a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h545b957fec207b082019fbed6ddbaa3293b2caf6ae0c91e642a18363feefd619aa4a967deccfaeb3d8b863d3be4e5ea8d66dd5cba07d9af41d88e6eeb519a355b8380f99bc41c866;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb87e44c1860974e69ad10fe84be680091b69afcd86227a323e9e31504e60afe0c7eec8a34fe2973d8d3d9f282d52d2ddccf50ff05786a4f861575c2583e8f5f33d54fa02451138e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd71679b911a2e5efcfc54c1da23c003c7728427dd507b561aaa36c9175b8c025a04d42af64048a0bf9df177936e869a4f94fa061a8398c8ad10470f73ac999a828901c445114a72b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49a3844af28bdfd87dc85162d0b5b30804d3f71274c6a48b61fdaf44b9282c7595c42d2a5b6fb687c33226f211b46f21bb371b2268d81ccd2c810ff9b0a25a7ec45c0c6dfb5758d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8b8dd642c3ddf73ff0ddba3b9e674c7e7f828e40ecf5f217d2e24fc8b1bb08bf36ab74e112c05ecde841e035e514d92ae672c60679726dbfe3e6f1ff1c02ebfa6b0f9aa337efec2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65b3f2bec054708ca8d4e43e9f0a38e5f76d2e0207d862bd2468a81250822b2bc6f136c660cd74f30f7c03d22e14a36689a60c0595d1b10a40ff99914e82ba374e72a925ad818ec8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h765dcff94fd90bb7b74f637a8ab77dd649a9b5463216f81d38cbe26ddd076ac4c9c73b9b6647ff74ac5379937a2cf5671ceb88e3a2d2e6ad6583a115c176f886cb2c24f3bec851ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc312cd7f8a35c7dbc8662cee5132072772d6bf82cebe2672d12f45e4144ce782bf6b8e37d170e81b09b72f568c52e643e7ac7c6f501d59976117b1674f23106b2790daa167b22664;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1152f8dca2970d3541288c82a67baa8dbcefa7210072bd143771bf85987730dc44c509d62969efaf2b470bb474e661e03d95d969d36ed9229bd40783508a4bec9cfbb3b6e008c032;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba615e50da439a20277554d30d1d904d30d5ff24ecb1b66fbc017d7912bbe9187830999740f0b8246bc9568a9e2013683de275c35efe5cbbf20660009a872a6bdfb87a85e3b484b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h796a66c6e0c1c5e1d70ede834e12ca6216b3111afc00d22125e7857b26050b4cb66cd9adc4d4360a9ef8db4bf4f0fd97e77d1c0dd5fb3615d29ccde0d04887530ffe55f702cfc45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33fa153473a3fd5976725a71e585d5291fe5e9eeb4685a69049a0f1f95042eb05757c889e20a74d6eb097bd10543e623c6d88309c4bcb17cb7cda281a2dce796184b9a2fc47ef8ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa3401d1dd10d2173076ee847b465cf529782d7582eaeb18d1930c8b01a048d8d641cdafba2860e603ce96c054d9c41062b1235da83d8264c41321aa002b3b53d5f5838b922388c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha08a534cf0c9f9e173a2f32e6d92c33b8d91bfd393d270777d2cdab314455c13e12cf9a791186ce3a406a5686a943a958afbbbb3f65464c31036483db777598e715864db7dc0f1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14ca4e656415c4c9b2c0af8167555ebc6d28c9e8b67349c6632b08a56fa51c4145344b4cd84071469a438a0c2d019f2c2b6d0292e24cb6a39ec087931973ce426f03c417df0ce405;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30bbab401bc970ad19324d47ee624469ca741dfefad8688f303f8cfb28c976f1539384f116ffc99688b78ffd722382f1b4f711e2e01059850811cfd108741698cd1b0ebcf1bf4f5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d6269fab7560252714d5ddf90e8b877db12b2a5bac179c80403110be7c876e4540adfc0115ca021a13113164576fd8ca59acda383d626cf835f433ec295eb1957c8602984bf71fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e441b2ac10288a720ede32d664909b0cf4c39084d65d8e6806e16736c4de7f276149c5150a5ded0bcaa467c7ef46dc73e65bb57fad5a80ddb95e08b805b583245a0c79fe18a7ae3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc399ae7487a22882543f5a8157510a6eebd693eb0d20e0e9da2d416e52ccc90c0bd9b20ca817b814a20a35c11cf5b5c45897cf5e7b0f1f8fe568626db27e6e7a753a16c99b99de3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbe503ab624f4060982fc291b55d772fdb67280d6d4b45349c03c58ece26ea371bebcbff8f7ba12f246baa2515e4298ae478b1a8a247818892d10dad6b4b7bb718497e0614d95083;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18f36b48b70e4cb0b4d5904650cc810d09e275199ecd00850c0ffb31d62cdb3a186a6a1dd93ddd9f92c3bbccd781a69ceb3a8ba044fbd363bcfc9345642295fac3cd38634bbb1d18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0b3dbb71703e02763f58f2efeb65b4fb8e677adbcb8db1a1a3d46af0c150699bfddf6d4b75a1e4f97893d57db8d49d26c8b667725f87c2288660a585a4622175e95dba4d66242a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd062ebe17e6d0b8f38c0b15a4c17a0b6ebef2f780b812ffcb1c88b1ea148faf8747d8a8a506ccd6904f56bf63d4ebb4bb88f277d75717bef5e5e4d63d4a95ba32b9f6b7074192103;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9ff110d17fcea689726305a32476c6a2d8dad823176012ca0954a26216e95e03f907819115f3275583f23f9e57e1bfb7c7582374d4e52a7b9dd8c032e5df606bb408a120e7b5774;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62abc4d881fc24196b78e95d11263c03ad6b61ac09ba854be164c95748e3df74b4ae3295a23e684899b7d76b1ccc9d5af4bb7fae933831603d6450553bb3fe53cc90c72b73bc3c49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd9effb13afe55dc6fef42b16d4ffa5eef87bd5bc2c9117df7e597dcb90a233f88d4f5a84df65893ba271e7007e8a990ae4f62c7005037834c5286270704f877aa21a15dc0182244;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d5570d704088694c8c4439439c5f16ff8fc80e774d11c6ed8f73ac4959ebc799804de1f39ea2191ff0ad995a50b7a53e67c75609ec00e0a93468c317e4f79fffdcdd36c0e2e3563;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he491b4f4f823765708d4cfa4cac34d90983cdd0ada95bc11c08864535e98aadde1f946b735fd0c4475ef7e1cd27f247200557bb2531b82ecb5e33ffdbaec72a062a738de0ff12308;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb682f0fc5d6c558a0f3ed60b81e9ca9123e9315b2c5e0ea8abc2b9bdbfb1e2d9910bbaa6cd6cb0b47fa1e32ebe9a10db075271416f8bcc9ee9cba2ef435bf3176c8e5b1a294d82c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6733c412ceb66e61d8999570d6353ccbe6881e5ab4b5965cd7cb4cc5932b2e49ecb60a4b42dd8a5e5c91addfebdc0cc49783901df027f8c811d2544214088aabae964409ad8466ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92f1ae4462bec387daa093bad838e2aba840c8c957e00cc949a5d123394e614d553c51975fea50d169e634d19692592193739ac7e3e3961154043e9eb75a65dadf4b10736e49186a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb41dec90a719b6f3bbd0f3e5c883d750f19cdaa88bbcca34ba5eee0b722fba5d8830142b10efded006ac53cc6db99f3204cc07c30728d7c7108131fea363e210ee1b3ec8d27d0254;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6261bbf3d36e5c50abf26a19d3e067d1830743ff4bc6bc563b513679e5d3c94a768f06f461d265f6fb787c4fb5201513493c60b83fc831fdd837c099b760359feba2d87401a52241;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2b47bf0f19c4e3e90858052815a06633d7290bef311c2d629ab4dbaf59158aa053ec4829f9c7c55d8d9c31dd7c5fb7f039a8539ecf57252b1dac00f5f70ef9d2662ff1c96766fd5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d59e414a5566f2f6becfcb661ee01ca7fd3fd08305cb2dfe23ef4ce755fb636b75a64a5e20a02b666b3a695870e356992b5d0149f1b13d3c7e16787513fd0c7867caf0181469b93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h500dfe25e99176dcdccd4f4dfca4c48c66f5d1a77fa473d86835a6879d2692f9bdd26e0be4beb8bdb07f578413ee309ddeb55be11462e80f7a79a787c61c15f0482ee9abbe5dacc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9e3fabbc3147a8a4ea9513ed21cb9a541683679b08e31651b40d7eded8c5476aead83507c4f00428c2032693c7fef25da142327ff348647922a437e45612297404a022ab95021b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d8c846ca9e5890f7fc4123146d86f5455dc008dce858a31d5ba98bd6db1074684574051fd60faeda7c1ece16a0132824c34bd21b0c7f39ba220d7d18a0ac5da5203f11393ae8353;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca24c1e1b912fd65511a1dbb47c22903d9d1ae6470a64d1cf5b9ddc0cc11725d2215338be83d8ee9d24f0d998a01620c09dd5c92a4c41d1e58bd1a12a731e70a3c38915cb2a093ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8ad1a29503dcde17c5bcbbcc832dde3ec1230b2994de80038aba0211b668879b3d3fee1d8dc622c5c9e9bc8994b4eb25769c22d524faf979a1cc81ecebb9dddbf681661d089f5f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86577ce35948b9dc9d785fb701c3324928b52d93fbaf4d4d6e00b42bdd0f52c037ffc3f64aac1af4abb8236e87b3e339810a31af8723bcbedea01296a1685172e1ec7eb7e6d38c77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8c2437da447c0d5ca6e82dc9e485b82cfe679a3f6f15f786a715871fa38630928df9bc24bc04fed7d5c0c7890a9e0ed49eefd16313271cb94a4950054770fd7ae8f1e8114a600f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc005a131a149411ea54db5798e862dd2f6e233faa3311941868cef01da801ef98d92da342695081816b3bf467c0be2d3c0c97a3a6aa0ad3859d5fd260e7b9a12e5d145f55a743dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aced5f6751d0fc036bfd6dd7c9ba59289426398cbe86e54bd5c4104c0f42c3774cc16a416af50a4dce39d24292013b07ddb38f75ed988d12e33d31e933300b6762b3c2862f69124;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h423a0f015bce02f7dfa32f690d2674a84559700f7793d6a275fd2ead09f8474e894d990e8e861f0b35f32549fa548736bed2584fc7d4dfc617159245400e8c05708ee268bcac454b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92c16c2940c5f3955bd36970756534266015d8b13a36dac6810a622622ddfa6a0a5c29ce421829e9c301fe97707de69879341d22c9f746751f28726ae19c707402c9a7ba2e2d80be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11ece0f102e6f3e2201e7002c8dbd7684b6e48bec24556debc42537a5aa4b2e438a31d2901ab16c04b9f813718f3a131394a87a8b1e1de7d4a19166b1989c0bd9e86973d40b21cd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49bd4f5e935b3544d094e0154f17dfb3d31745c31497efe4a554cf7f2380ef067dc1a15d9c36330435a35b7067327e4e25908b40151cf2a6575b189e4510a9806029a544d2069d76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb687e711992dc6c9d3824d024e424f198464183ba09451abc90449d808a5b0f0eb31fbe5b21e79a47548d81cff0eabda6dc459e1763a079d589955ef44e382f670867e89752728db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcebb1770ca9dcd5e7b22c334111ac9a4b27f0fffd8c8e2890cba554b1c17bbbcc17d7108db602caedce2189190b45d6b36a5a191259dc3bff3fdc8f2dd4b5d14beb7120df8cf8595;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13f8b22d7aafa6b709b102e3cd1614ffff29283e9ff8a890837cbd06b341a51d7814bb7619fa938afb79137fc00029448002e842f0883885cef85f1138589bf4fa0f1353f97aeb30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91e450d52fb5a9de3b13c07adc21a987151eb7beacf7153eaee59d32a4c94747cda11966b2d8359cfd0ae44f8d80ff7e679c902aa0bd0086725b31d17b4d059fae789fd3bfc18171;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc205a9ee87fbf7d08155185c47bee3b7a8bd27139daa8d5f10aef14f96b04c4b9e7709fe5187b11f840bee6e1ee2723875a1137b6313da4e321e7af49998864fb51bf73563d87bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36de0236df79c684e0f47e8e50b03cf939054c3eef8e8b727192384d6c1b27f4f0c054035b08bfeeaa166a4f3f15e4acd6071fbc3f5f437e2c064ad825f1fa0d1ac736726501c3df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9190f9d8f37f8ce805b8ef4abfa2b45f7e825a597d969d27658db955a74b4d6c61a36357a0e749eddd635e8a29fe01f98d7c16f188b28cd866bf6423340b4847c33467d3477f21d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43db21c8bfdd29df0a4948dbadc872dcd5a1def6afd64e14cd71889e52a729dbdb64eaee37da39b1b6b33c7b3b6a0a081db57d1bdfb69b68c58363383d072bdda7f52621e4e9b831;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26b442933b8a82aee9da6e89e16c54ed0547cdb2132b622ecf71656dda554a2b25046a3b4d24532f44d83b50539be737dc8daee12cf708107898c374936af9bed59b2d27494b3cc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8ae46ec41558af8a3b3884ce754557c7589b0f0b032b340190697c4253332a2717c93110fa98737ab55ff3f7e28f9ef14fdbf6f4e5aecff915b744cbc17c31b90377cfb55bf05a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h613378fca0641ea1e1a398f9ad690e1e6e0446e27522ab5fb1253a2770efb1201fe9d318bf22683fcdcfdec0ad5cbee70df0b6709c8785d468865a07d465982df43d343b6f3bbaec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b5cf596589e083c00fd119ed4088fba2ee4c247d802cafafdfcbd5ccf177d09ced8af33e2a34f520a0eeaebc59e5ab780bdeb236904ab22546b8af00ccdad5878173f10496afdf1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h530801179b7fe08df5cd55a9f4e0e2b72e9ece4143e1715a7e6242143d2da2980763868642bd3337ecc7b458e2c3b371f5cfd58a7eee9894655316a86b8f1435d99325bec3eecb51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef143e53dbc650d72d7f879fceb7e22ff0511c91dbc81fa4f756c276fd2980b7c3dca8a42862cf99b0eea302e8c4ce12e0d57d8322b22c07a80aed46d3a184b871af996cacaba6d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36f28f23195a8edf89e2fc4ed8365254f849a3af20d150de7b15afc2d570d3c2e22a6f3f6345f59eb65a38048e6cf74d28fe0128f3a6cc0bda8639e58de513b4b1c5982653d1fd6b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14e9d9e96857e0a1adff018d8645517b114663a5e74f5efe4f8443707c05c2568d7a9e1b0c5081ed44fab1d54d4aa40c1cbfb3e262454c087b21cab241c8189de289ba5e528c5e4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h741f8d4cc8379fccfe0632c2eb487872f2115a902902f2ad9dab6131c25e6a29c1dc36488949707755cfd0bd341c1bd39e0e73bc70b9abb59011ca978c4277efcf868f3032e59d95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4165570e4163a03ae2381948cdf403fd07acbb47bdbb07e834590c5680774560098e285adc068efb61072e0648cc5f2a67b0033b4c977e489a2f6c8acb1f60b7186e67263bd003e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c219f35c4ab48ba674fd0287fad4a9d3b5f696fc93e08bbca487ee1c858ad5c83d83285775149ce1591d1dbb91461844bd9c3b7bbf753c074745b940ce05c9dc3105a05b4c8dfed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h549d172ce335d45d227d38523501df1925f32aa5ce16d75c3f40adea3afd6bdbaf2884e2ca693927aa8328f291a1930341dd0931d7c6f63954d2207a72269e392b79824d3bd814b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7724d772d34818f99bfaecbdda370096c9ff7089476829935cbbafee83bbf6ab42c1da419b109f02323c268220cdda8d215e881191325b9093054e710550d92eaa500b9942492e08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36ef289f9bc9c195aeac04c13d51916069df2d2e337b9c5ff3c2c03355caabd35675305de352d3688a64f2c1da705173e25d03c8f1b1ee914f4beb6e3bb0b628ee9526fa6d9509ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0b46eb427043834a94b6b3fa68d506bf77df9cdb35aa954dc9554d61b71e355f2d5c9aaf4e2fee797e1ac54a61a8602159eee0a24b09b2d23b9c3d8fb86705c3efb5565ce130a8f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he088a6c970cfe289f61106ece237882e26ecaa8b831b783f28c58dc7342db02189af6b9ec037d11b55d79040dfd3fef0eedd4b816b7e6fea9543ed0ac3ec30aabe403b2fc26abe1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dad05830ff1499bed710116319e4821c51dda9fcdcb517e08ef19d154308274ea81b13984a5fbce7d545d46a711b59868dac747f424eae44f25ce3802ba33a1d4711dee17b2f168;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc704638ea2924fe49212172585617f1c6de3e60eedff4552bc51e9893d0024a11721aa740b3981717712d318b99955ce48b45f91c585b8f98307b1645faa6450e17e6f786d684957;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h662674b83bdbff28f8e3bfc3386e3eee74dc5d0fb0c7adfe320999875f2b033e374eca6e63776822a2e04b5f14c7ecf7ca1f65bd3eaae18cdff6d1ed4c26770b5609d8673b76569e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had3ba423ba7ee361f37742e0cb2818bebe38a890418de5fff1ccca8fe29d473fc913ab00745a329bbe46052402f592448a5ab8dc2ee62ae2454e85a7ca3ad99ea19d8bd0981e050d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha864ae9df93d3b1fac471efabf9f15ab33bb79c4751cc1729800e9dc691f3325504be1eb74d4bb0eaef4bff8d70373ee7943845b6bc7440810d4c4efe1716381ecfd98609e70c260;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cabf5d4e93d26b2ebd58a27d6074f9ac4186afbaf17503d8f6ac31eee4e4b5e9326463ff98f57ec10ca2a948d91b9744663ed652ebe005d66e38b12db645c6a4a288a3b72a30e80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7761a8f19689403b89eb2c65cfff0e067e59b02661bdb873e8052d77f6f6d938c85f2be8b47481089351be30a43b2a0e4b83b075bb0cbf8e319b58ed8c0ccff4f3f52d4c34cd11b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h550ca5b4bafb0f9bac0c1a670032e829028a0ab0e41ebb0e42541c3a4c63d3d924a3b071c78bfc301f98831017fc887203c117dd96a93be67698a9a436327cd204566bdcbabcc7bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hace662e8a881b0a8afa56fc13f2144748622f6bb04ca6a926069546779e3185452f915c8d65dd6ecb0233f493ff686d07d6f3c538996ba126984f835e119d0c6a597ed9004d78ec8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fc7959479db444764f1cf777e4f6d0ce35f76c7cb826f7bf720bc4f859596d35e50504a91b74ec18cedec98336f8f60a027d11697953407814b1c20ce7ffd51f23998ba639c6b13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d20ef3f0be3a2efe4c2ef9335f14d392524cc429db334fd2e8e98093fc26118aeb774100cfebab7359cf1f24224332b08667919f9858ae07f21313bb91f617147b6869b5a32029d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h135c2791810adee92fb3a896a036957936dbe90dbe4ddd7ece9a7702616d8bcfea453193ed7f1785f32d3db46b84a2754c525d91dae6b6c819c9d01834071e26a6949175f66c4f7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd83423a260690f5d1b74d0a391402a46deb99980775e0fcf421815e99ff2b3f404c08fa65dd9edb8d0608973dbede670f999f6faba56c8ca97f3b9d96fbfc40a170dcb3cc1bb5d30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha442df5e3b65ae7137b8459bfb45f1f65121874f60a0938ec602e7597d687a0e584185a272996c55336b20c665750cf9e7bec7d1b6cfd89166a9a09ae3f8a0e8b99a5144163441dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5069666ae81f097cb6dc298c4dddcf710c5d66ce1ddc9664e03758847476297d71bfdf48d9110e4727e07e3cd99bb2b7110c3032726fcc446285bccb548a5916d7b2c072c25465b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b7d50d576eec98db0a04e6a7e0b17207b2e740ae535f4b0734c698593dbfdf48354c1951a284cfa15505187a6ddb02783d3c1b87d95b792b5bd8adce770fe11724daa179b3e1256;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h765aa638664db2cee33ab4a25dbbb32803e45ee964f8fadf4114f10617c92227c39ffed6ab5a392ed0600d0b6c3187b922b5857bb95ed95686ab50012a854baabeba7c77cf09d372;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha760c096daea4097ec2660f0e44c1a6e9bd1eb76c8e7210bedcecfef781fd52768dc4631a754e7f6e2731d8dcd5467b00d966fac29dcd70ed737a490fac47f28b97806fdaeed0d1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2206f37f8de9312ea33b262a956d3dd2d29d0502508eb4577ce7708261115a147a3ccd076607ca93420c2468b012f9734eff5dc666786c09c5ec521dec5047d35c5fb170e678f0e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6917288c30d9a264e2fbc0d0fcac15eb4af12a3ede5d956dfd8d5e6e249aca737a856af1de1690fd448a7b3b8c66c12fb7baab917b4fe6341b03fc79793560cf0a34fddbaaec1a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb26a2a377ee75980088d9e5ad8ccaab59874d9e161b844f3a3dd4565bf8825c91be2ce69149244067fafa9cfd122fbca011829527e117bead15a88092e35cb843f7fd5d05351edb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha561f1e49e1988a0d3954c79f2cdc7b010ae9f6f9d59c696b5fa14d513ad3868f6f5b7235489908808828db2c77d2c8aae16d4f03ed10ab85be30f21e963ba358703f8be6b47960;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde50e83d1ac31f2490be46133eb14e7e97db1826387ae5c92c752ba9eecfbc4bbfe43088fdcc6bf8150773141f0e64f5b9fe176fc0c911cfddc54d6799b975d97331b015f6897ec5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c8ce0e4d4fee72ed421b03bf9790781f59e6f1dd106d3efce1fb70e944180355136341a0d61a6761d8a339998e710d975787f19de0aa638e40b2c8f358afafb72a33c788a7c3fc1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd42f10b8f2d06a492387d88ec5df3e0e3ec5ceab6789601d1d5b0990e91d419ad2e5057b43858a58ccd51c20cd415d9e8a2fb91a12d0b09d68b50a39bcc11cdae635a95b9d022dcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f3842d1f3e9635c3d9da0b2da8e4b1aeb0469dd3bffa38c3caef964f86c267eb155d6666d45c6d68e06f5a8bf876ac8b4daecf11a8b0a3099c5190c198044252dafa761c8d7333a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha26c07351d9ea739cc7f665f256c224709b133f06a621f352ff551612b3fcce979a777837aaad85bcf2c1d7bd184d6b1ddce920cd7dc49c47b5731b23e0942c2ea6524eeba2c743b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22626277d100d6f1e20528cd4379f3db7de464a37ecae2b5e12a38c9caa45be73142a5474922e6389926eef7f2e079df537f868bbf03962f464deb846167956e824e7b8f4f264931;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea30b80bf3e3f0e0f161bfda28f03ab912e278cb4eaf7ae09d479edc40166bd7fcca9e13eb487b470c03a0cd5b219eef8ee3a2c7d009ac44507a0a6a632328ff2fb368e2c385a4bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2321d9c6a6b922b56da6bc30b12e4af3077b6de51355bcb9edbe2674a0705a19e3362f291a101221aab870035412ec480b682504145aa6ec1f6ff4bd4307869040d847ea03856037;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc11de3a67b76c1e86c74d90e3de2d72d62ec52f8d13a137af7e0e7ccebb449c3f827e5ddcf55af1a7d577c7e9d2b18e1b61cfc627893525fd4bc16cb800ef4ff8a68dbbd38b3148;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6090d04842b8d7e91d609bdfa4a908bb3b5eccc23a9c431572b851351dd632feaaf4ea4ff1d8b3c0036f1929aee7a19020e402bb13b4b5757c28af47664fe5732a6937381b83d7d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3478ed945eeff21398b5c5a59e808cebda5b59959ec6f15d80d5f7c31326b1e7ae424fd321f81a2f9bf85e862fd3126e3477c7af3775acc87e751aa47851dd8592f545ed38587e53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8744b075cef0789d7a76173fc1aae84efa1f84bf166986329981d755534ff9c1d6782d9d00bf3b309ad00b3e517fa2e21ee5db5ade3db0ba18f759b0c3304019d1d5c213b30b674a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48d4098611e66c0d54271527d69326d11f33126e74167320699dd7d9597cc32cc6231952d1ea850b032a1e117a29c59e2f1cac6325bc12885bac7865917edc50decdf4e928ecae80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32e8094ffb9a788c47e25c1b56dbe3f867474b9f32d169800a21fcffccb1752cb4d99abf0058767573a047d3424f530c20af33842270353d5de1364b528513fc4ee9f6c5d67b1d08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51dc0b7706cf9b24d454d4455d77d8ad297f86718869575a4e991d897fda4abb8795ac245badd9d80357b4310fa9be1d72cdb91dbe4057fc82e1171bc4cccb84604b7db06441528b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h779f60b9ac224e5b9beca89abdc65233f378134a36b1706bf7aac1a974d5e4a3e7471ecc6fc26c7263a6192e5c86adec2d2964383d8e61b5af8cb434397feaf5db5da11360bc24c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he82524ec7f4eafe65cdc53e2e09a9fdb387d9b7ae7a42379d7c7b401be8219d0dc9703e8c2340527d00b1c3dd27d29f16aa94067d486056c2ac419ea672af0b4f7111f262010f975;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88f8a0f9f591e26dbf22e5b55cd9dd2642607f0cec6fd5be9d30817a9120780b72dc30e6b6acec1e1536e6fffaede1e4b2e212851fb3868ab341503d168c0c4471ddcbe50e0c7740;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc7e8d950f8950c59b974978e35c06c5437a49d74e892e49fc293e1ba433eed285f83fc31697515cb13ce54ad21bf05dd866a25b1ec3787b8800499cc8f7911ab35a7779f459f9fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedc646c6b43a9c8d2c24c08b485c91c60fd35ff1e5d02685260aabc535d9f121bcf02e7c05117c4c81bea920a1c82b1901abfce3e470dec9ba1878d75f1942d679da0f25da92e830;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69393566f67e215352756f4deab730fd488c03ca75bd7236ffd44e0bad770bc73c5b2b1f6eb9a2192064a4802e79829d81ab75fc7e96ae5e58aa49c50eb567a04dcab504741b0af0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf3f8fb302ecabe31965e23a772466a26868aff83f6d79ca940e47c6df83e28689f03a2a4eca3abfb643e825ab16683c78e8996068536b7256e87082eba1183e754e9af51d4646bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3267ad6f627e561262279503376eae42e41411a406d0586bee74495e9dc3045e4c7be9fc17d4be938742a46884ae2350ac44c2ed6bb7d89ca5c7038288a5f6353a12994ae28aa098;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6799c984de9e6b33f1ed8e79136b5150690dd911f494832cf93880fe06cc6fbf41f93b99ac65ee3c6431f982015bc070671d227cfea573e3d7f0528fd4f38ebee195d00a262a1033;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h705507f9ade0274833cc412fd09ed96969c2ad3fdcabc0fa42cb34f25505fa74b77e895e48b11e952e713d73bfed747bde05cb1c24654e202b2a18a87a0aad592172cd5e75fae1e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h655ca3ddf47deb17fa402d1ee73d6b801ed22f69fbea81b69a15c6609da9b4565d49982f302849ff7de0e8589cbb39a1564f6a51bcdd37137fe353559e5108f3988e9f189aef9c0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb97ca70cb237add3990b967ca3e6dc3c05e8e1306aabe852b1e118a3b910c9b77f74e8da43948cf53a79f5a87527beb4c0551315c6bac895a012cf3b17924637025c433e86ef667c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41cd2fd1a78076fd86c319a6d6575362516700ca2561e330d846018f8273bf9f433249d8a5791cebbfec6181a5ebdf8d30b46ce6bb543196db41b47e27441361c0f36425f3bf55fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0eb6f79e60fd8959de2f1711a142088b601acb0e01ada03690e0a7b7a4f63c6c3298d4fbf952e2b2e96022ecd9a04aae192ea906c1d3a7bbb76fe8b95ca595d2043200df9d84138;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e8abc5fce0aed1fed96c2914158f3883ff80ebbb34558532a7100eaf7480bfeeac70e0ec9f366fda52ffefacff9c8366a53170df020bcecdf7d9468f3b63fdb34b38fb526433774;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f585674efba05195d0a8124ba98714bacad8cc10c954c4aa95c9ba7c77abe1002068910afbfebe54e856ea108f47d7219df7fd3c67b47efed19d2f7b45bde72e9ea838336647d56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf34aca3699ec57bd0106b257b02ae9bdaa34bfb368c87cddcd8d7b6c4eb15b7fa245ee2285fe70cd397897f39366337a6e4203f162a5b2b4758c1d788cd3ae0f25e978025775fb1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba3fac45df39aa40627eeae5f78096667dcf87ef9c8358dc3ce058baff39742f3f03b0fee7ce1d0de305a48663515fc65a0142dd926e02e9646adbdb018c80b3f1ff871e2ffc2987;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he18e847a7b9573f52c8246c904fe461c7c1533d57e12749bc799cf42e8446e48242124e948f96c57b21a6837f2d181f2882fa783551683e3b3295fbae1af9935c96d547669c43651;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h702d3cabe24a2c6b5902e5fa82ecc15ffcebb4e672c9d47e561deb93f2d565e226610b43b8bf19ba6f9f623c571347a722dd8a0ce50b742089922d07315034d45e408dd60ab5cbf0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dea47c7799654da0a211898546752a264f89cb1e52f4d9833f0e70dc9a99d181e9425ac89b13be46578d828f6dd4210e8c6b623943a5f3b4da158210e6e3a64e18a4bfcebbcd8d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha795a205f3e13c8d5f2a4c9cfe23cead6e059a89021a8c123834fa8ea4ae14d70fae42f8b29dee1b0730d62be482269c5cf23e9bdcdb9af0c3963ca6575de551f9d9a4683dd50407;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f28f2d728d8264e3db31bfca89fcdb02cdda12a7906d95551dc2155aebdeaf0e1f3cb30ae39c4b75d67ffb058713d0b66127887cdd447550d27c0edbe405e5c7e6ed68ea0c89032;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h467b2ff59d0688465b87f5db99b120f67f683937e6ffa29d338fa7695792d830889efbea92ee69a0b596cf3079c56f81f3a406922119e1846ed6eafed2a9dd5cc6296b6a0956a88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9adb39709885e27358e3223e34b164218e388115d30e2463a04f895f8b05775b76b20732d0da060aeeba79c29dacc924220e6d6777bd0ebca479e33043bfd718add31642fe395c4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc513c3661b973ccbda142f76189bc363caba9c23147fa8e26ec1ebb63b8e433f0d85c71580fce19a3cacb938861416db9c69b443851aac56f1850b9ee1570956c63541d7e61efb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d09d1e8f0f0bbff50fc07f26f2cb826ca20e1b5cdc2f8b69cbc3230f875b16c736e7ae75f2cbbec3643b1634f64be368e1380fb98fc0d4bc873a467fb29017b0b77d2fe60b6281b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0a239e937bee886f41614fa7ca7f9c3d5623bc322fdc129a2b6ac55a9ba372361a409df5c075a01b7c2781b1b00b10573729f4fb1753a57c73e015a793670998fce95cedc5632df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31b6482e585affd3afa615ca0e474a8987efdf3b2d56c2fe0835dae411de5bcf7c23da034520eb65a0df37b90cb2d983b7f493b1423d4560e5d67aca3da4a82140eafe06866690a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3979a9e38c54a3f9cdcfe99a046f570311a829ed8d102eac34a7f611c79af90d2c4660e6d56e1efa41115809421d29ebcfac31e40f031dd677500d8d67f348a0f9120582f710aca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16b277ab5f573a51f464a159d7b9c6e55e22d7958b9d5220538425218d8139392a957c352e9d31d301a3647831f98d8128d23eb5522ded69b2199e3b5167982adeb748ced0e3d6a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb46757de7ff01d3d916ca2429fa8e9b108c83371972ea5f0e97d7ba49c86e7a9033b68a3a0921446bef7821e35d5d5cb97483f86a8dd0972d13582254853004bc18e43df142841;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf81e591fd41c865dee0cb99d69fad9c6175b3d01bcf30a152a23eec046d1db63f49c44180a4375cde5596d3c5163bd2282853568d3ec0c15511a25426f8c3c5a3aa56abad0fc3daa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99584b5d57ac3bd819aad0116789e8dbabc68353a986bc7a0adc04e468a34ff8f3255f3cd442e36b59a446803d7beee663df810d2896305e50ab2a6df3c26114b3c5284586d809a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b27083f079d1819b7086f3814aa64881b526014821dd7fb309dce7612d7d75457c80952ec5cf19dab14d4b717b558d06968319e02d49c03443d2a430cd6632799886ff45fd0b0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdfbffa23fc99b7290680552fcd9ef3ad8d1b6cce3643176fa1378af24772a5ea457e9cf5836b4b4f017af5ecbfbf966039024c78cdcb9fd87a87ad8c67b48a1a08f2914080797f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e1bf8eb9a5e16460d22922affa575c62251e87ace6e0149838233c4d3327e23a5c0e1cf76b18eba90f30fa3dae3af71ef0cbd7f5a715d95076a5f1e968244eb5ac04dd860cfc7af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h132c17bc981da990dd56cc2c73d0d713a3893ad920024e105670127bb5f495e9439590fd1f9bce5ebf7b933cea2f95d843e82b37b9042831f30b3d18a6a684f2a61576a6f371b386;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b48169105f5199d262771a2a335cf8031363f197aa4c7a8ef3a59986b828958bdead2aab9e5bb3de9e716065cf916dc1317c593ab15c6b4998c5d946fd5d769b1bcfcaa012759ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfa0e7c49019b3ad9dfab8ca326cd7297f7030633f6167430ee00a2f5498d87f2db4017f9e78697fd06d03213c0167f688573413365db38d2e676af8cb2ad4f27ac94af59940a02f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h412e9d5866f4c603e2746d704c23eadcd4df02791a27df1369a9de6299eb1d71fed5a7042daa42236b91eb6e62e32bac2e74a0f048a2d843b945737969f7c6399987cf2e7ed8f4e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a0f0787cfc475bfeae2732222ad3eb125405b4976a3040f0f1e6d4610b97f3b4f3e6a41d868899b0f4690953f9bb7bb27f03fa9b975b843e4f62decb7c4f2d403cd1828185b8aff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf3133ab81ea4b362bafc10c9f947f9eace6ecad3d6f1d26264ef887d8b05544464f90c1aff684bc602603b3713f6ab0233fb2ab3f41e9f57b9e69d63a8cd8e08e7bf5d09c976b7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68a5850c7071e33419273a5bee19c758a516e5dce232750c3530bad73fb5e36bb89fbb6e3bf38500708ad38fa440d86f5ff4dc7860ba16f8357289dd45d698ef2503c63c4ec47a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h500496068f7519fa33ff87f45b0bfdcb2e6414b4a45e2dde12962be5e3f39e644c57e9796b1f6a85541cbb5391b79be5a2800b87886af03b353eebb9f5ea191b820a3807cbfe7292;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he651316eb706b360c31d1a0d6af82a56f0932c079f5f9855783688cded1c23fc5d832273f87b2b1be0d4cb176df5bd668436c9cff313a4e78c275ac52898ffde2dc79aee38b0afeb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h129b12031b14252bd31058157c3dc280035a6798d60b292c6c235e1af3d10dfc2a06f6a6cd56d305a7c526b73916db8185a54a68662e10f875029676e007c17e9989d298b87b2b2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf9b7199a6d22b5ba4375c1c84a998b86aa48e02c8f75ac1b0763a97624a4ffa713ac3247ab4f5eca5a68472644130be2000bfd4327ef769ac1cb08d631998e6521bc5a4f40bb3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e98b4d1e80e3ed699e86074201acc5a2bc95355918ec51c4820010233fe6e8337f362407a2618610638039ba90a4ae64aa0b272c8ea3e363a9a8fd6f251faba0693b7f3e70deb8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce66a05c19d829da85d47ce277db531809bab53fe4feb39ef4e3a40f80cc13fcdf59a4895e3403f3752ba7f33d9bcd2d33f9d4be56121aef5ae454ed47a61696883e07a04c295b47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h277032849b6a1963cbb1e2f1154593be9574d21def250e4804568946588b606ec4fe33adb8f2373a0fe4378127026c77989bd7317a8da237bc188c2b7432d51ea04993cca6a04b00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2561b9ed2f10b8ec07e03b3df5742ba14c8a6ca25f13a4cd0672a2ece2afe4b702a543cceda3ed9316ed3d7981ed3db96bde68c6c491526d5c56e21b1bb61e09be39e866679b76f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26b29e5ff7f0c7b5c1f6a0839785d5cf439e0da21f5a62782259c08f56e6eb11abf9e87ee92708351ef8ca3548527c7aab5f27c51402532827e116ab9ce7867f893c7887eb378f67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ea8f36f5f6d2907d46b190aeee004a3454ec27b2555088897028a372424ad34072470a7ac05be27ceeaee848cc29ec0bd60b40fd665fb596a5fedd3ef913576677ed2ae750afe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58756a28ec4467f5cddf029d98582cd3696afc03dd2c11a25dd031700ef315442ceb596564498d0e93a49f97e613d94bc89856dcf5f8fa118c65e42fb2881e565fed20f9aa604afb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87695ed0ad267fdd5a06aa00215f0aa1e1e8212bf9ae505b0a879831987a33fe82a5da91bb929052bb747a316cd64872fb2c951f28c45e7a7484c245191fd8b718a2ba40bb931bc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea3031e5d255942eceb772eb3309519b88b99c20252b9f33e5f498291f7ad822619d22810f860db35fb22a41b326e824f0e6862f45d7ae892536cb6ffa1c65dbc2444da8e5e548df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb60e52508f7e91b3f264d78b7d11c1de2db61d14ab840a0c300cc8a0c380fac759f581a3f1ecc4c0eec577d5a304e5a172153d99c0bbcc3d42ac1ccb4aa2c0039cce3577dba3551b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2b2c1c7a562d8c0c1c65850c46780c397e4f79e3934c41e28cec96225c7488276dffc71c72c7b064acbc2ca1048e195b13e82390708583434151621108a12b24271486577871adc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aef0042caae02fe2ff0a336898135bce8662c1706e1fa6b84b47c64b1e62d43583c5fb1dcdcc3a0ec1a767f5a4171a3f739cde3ebe010cd57b173a0d82cc6950dfe62f4bb8f790d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h642f978049a86c67606be9c32157105c8c6ed652f3174652372835b3b6bf9d890c1c9e4be45dc6cbc390aad8b54d9a77c8a54b2acda46da7a692ccc46128f56b02ba3f1ccd25049d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64c229d2324ca8ed453a54dc4aacf71ff6fb6702fe1732a55955511cdf3e4c2417e1a5246cd9224cc9e192d1f1f9166445ea4e1f6fa2f28da022859a8c12987954dbb39e8169ce6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed02998a2880425585463c506db2010c0e5ead114f7a8463f69b8fda1e5d46546ff06c144f3c99d6adf897f277ff99f509edf610957614a6b6aa5aeff5acf8e816a8bd8772d2d52c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab4c28ca0c2004f3fa36bcc32cfa05eeaef162ae7dc6ab336ff6c13286bf8ef3b49350c82e39abc4e62f87e0f9870f9d687ee1f62d3991bcdc00f958a0b730646331e77d12d7b437;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2863de0a02bf9830c4100771256f8db960103b2a7e823e28e47760e82cd41c0548763268612821a8a0cc05af7c571ff7bd718768edaa0c54573b8df89b0d1fbe57f08796e6b9ed14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h164169700b2d46ba20c0437870982b989834ea6f966fedd6c61e43f421d4b16dd36c64e26e0dc4148dfa2632fd8c11d5b1f5237ae4c3062b7a5bdf1e1d2a6a0e407dfb8e956273fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h793d31f0f78a96b9ff6fd3ac37c6d3d8325c9f363e4ecadec8060f9ce57e8d204358b436f26a056ac47432d56f3632c28d81c970ec0a7b49fa969650d2aee3941c19a032b48772de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3e52a59b470eeaa21b1e9cd3ca38a5d8c2f3a3a500e2eb8e6d3477713ea0bfd1edf9e23a47dcf17b261959bcc2a4ed1c820b35ecd343b2d10135e4f4fc25523f8dac55a445e79a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f50c20421ebe67663c0a1c7c71a25eff6b7a522cb21139223b8c6145776a13de22b20d7ce843fcc88dfe78fba5f29f8df7325dcaa5ebdaf5fe1bb07b027f0e19048d67eb57f1437;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47d04e8585b04e6f4704ae90607fb0e98230cfc6992916d977518a3ebb33647e11289c1bc3980ade67448ed08b033cf03de5cc8d5172a3cd1266feeff37fe5dfec84323d9b56da79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf00b7ae60e79b465e1ff0f652c08ccaa7c81377f68bbeb0d8c8a450980cc2cc447c890b8a514c4899bc06b98d7790819e520af3de0bd70f5772ef0fb9b988fd85cdc506ad100ed9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5eb126bfe1eee7974a6f96f34ce75379f2430ac8e4001a83a3dd2b7b6f96ea4a37b789f34da5f5802e7a95512c9b071d47877768f07206c00925768034477e0db2190a48558949f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he05c1720745adeb07812d2c778a0ce558f4c64af0fea1974f7ac91ae938af9d391aa75dfb82989664c7b16f45ffb03b31a0c12b607c4b71b82506913e774889e28805a6bc06034e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h283984168df4ff18b488c09451c8892a6e04702c688549dc6a0ace3b26ed539dc625fcab96fa87e1fb2814b7c94f89051656a066c0179eaff307fdfb93707c1379b853b942e49193;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6132851877900893a6d5595b328399efccfaa0e5235db3d450ac405cf7c49593658871b03a3275ae4abd3e48e8a295a9bbabef48cf6f1fd1948c3418f1c18af17e64e4ed0c69b264;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h111c856b414c3eadd8fb4df201a0289e6ee40e6b00ce3866010739ae8a26118773b13bfdff5d71ae5e1cdf38779361f946cd1094f52cb0fe29d626f7931f9e8d6bdf88dce73b34eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf08c07092426cb2c4951ed11ad1ad56bdead433ef9eef4687afec8837fecfec9da733d7852476f561d2ad281620255cc726cf127de6339e5c62f40e777a98a0946be0dcc1503af1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fb0aebc1c1e4fd8fa2c381b60448915d59244f98bd1505698e1c2a57d7fc83d10ae699d0cce2ff010c9206d1344cbcee66a4663bf0ae4a4b51c17f0df3b2490e70b067fd368fa0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d98cb49b5b4e16130b9b13cfb3999accba2f4b066d8a536e1807062422369f8224f75ec99ec1c76cd4386fce892e1569f10cc556cb4407854ad0de7989f792cfca912b2a5df6022;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7fbd904aa029c066a7d1420c67f7fd3bca218ea8b8bcc93b606956e9099e6bad84e4d3f0875edb676a00d5ac5b309ac8bc9d67d5ab54123ebe8d5ac402e82785b7fd7d53305ed65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6ee352097371be9283dedfd0f120a6d56a63691058dffb1bfc14d04d4c42a458035981ec1c6f4650bacca25cd8b55cc8de0264177f6c8933d6e1ec32220224b847fac5e0603969e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7519e6b423a230f0fa212cc1122141e09cad675827c786e633a37ef2964bdd88f157c4c4637421e6c3f95e341b3d0358240c27e16d993bab1d210a371866f168952e0c38148faf2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf675d679901145d8c0f0d0d263c435d37258f077e67a534d80d893c04358bfe75973fd8a91984240c9c569ca8d94273db7b0aa4fcdda816d43138bee593f20f829b141ce6b0f1847;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf55b7f950adfcab1ed6ea601e476d34796dd9442a046c37a3337ed6fac2d05052c32897977b06b83cc6ccc3ca233bcaf1ba92c9be44886d62e6dcda0d5ae9e51e8d2aad163792a91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc67d1d904515f5d5bf64165065631b9f0a292aef198186517446cd19efe6f1e7a883dccbdd1528ad2767de2af522fc23bac734a7b4d8c3936b665fe813299bb65335539dc8ff6eb8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6b6cd153b3ee36b29ba1f69b25ecce82fdcb78f7322d6837b6bd9984c2afab9deba36d2a68e3b34590b9cae755686b60cde076b0989d2488c06ef6e24521c0e6163e846113e35e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafd25847f6cfa3b2dc142e576aadb1dba98778f1b6ab45a339f7850b006fc1f9bc339b80fa3e86b3499206c02660d9da24316bfea22e52f0341d5e8659df3d34b01635cc3057af50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a705b7f6fcfc4b7a5bddd64a134d70baf4761efc39e51f9e008a9a71375e4dad2fa187d80d9cb410447b6ed21b301593a816147c610aad7239b59cf876959e2bb0ffdf38274cc42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91705a5b4d961fdba771271b87865c78e68943fd6915b7c4c71467d6588fa2860e4eaa9993d0e5b250428d886bc82381fd32a9cda7b259191b4e68007db69dbe6cfdf439b3a51e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79e37d7083f77e667d24ba21530e230ce83c5f54da9e05e3fea7d85c21ae14939ae080cc5fb4c64fda07b44e6ce8e16cac56b43f825213bd77502b3e0c9c794fc4ced21dc12f8900;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h219b38aff40cb4f29c5ffc1e71dc04ee68349c189213132b9ba705c41a2968e7afa733ebe31188fe6dc4bcd08b2c0ff273bc97b1df33797fea402b34eb7bdc31e0db203f2d1c3634;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f97f0dadf703b690cd3b7d20862625c0bc61673fa6f94c56882814ae28cf2074d40709132f40ee82d847295764a6ef25ed5ad86204776e88f53e50f7926d353475155d82ce4b3bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h765c52d3baa6415248cd11c1825dd306c73e1ae356aada214bb7214ff1d1e154e00c46ebbabd0ea37d631433678fe4171e75fe64ffe9b12b856b61048710d0aa6171fd88392f78b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb06d294da7588d817461ff44abbc679cb2b1ef448e8bb5957da1401449af27e018701265300c3657264dbb2495dd6ad6f322e6123bc145a1923cb4586644b344ac5c0459f49ebb45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5eb2fc5bb15b66984dbe008278263b80af67c3f7115385e94c23d24d873b1af022da69c00768367ff246cf7475dff9c08e58829bacd3b2bf9f63b31e6302f92ccb172b119c272d5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9a2475b20d11ec8b61bd8de19d7f549a97d0a94b6a85a5fca9bb362ed26fed19f3a59183e9bf05d78212b48bb243fa569517e8ec04b2a4e2530da7f6070220b147a17705519519b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f753e2487d6b2b3dac4cec3bfba9753dd6686d9b2417b49f7aacd84a73e2b78a15bbf6ecdc89b5a393980613de924343e2e8422031408b52ed220aa9ae8afff8eca8074aac488c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2031f70e738bbff24bd0db04ae6b6e460830b0f797441b114fb0a87fa5a6792e36a3377445ccec0b1896492bae77cf034d4cb9fb6e883c7ca740ce9e7f7e12d0ac4337213854858c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haba20fab94979cf3d386c79e37cedcf675f3b756d6840e2aa593af1840177db699ef956b82cf7ff21a8402d6d96ed3a1c266984f0ae0c1d2ac7d44d34dad4519ae80d1dfdc60af01;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0833affe53c3743d03597f6cb98eb6826ec48da28fb07935c028c90bde68f9157cf7e3e2b84b3ab8ba458541584b54ad1e479fd9e5e51241a195c17f41d9e59e9c872e622b7ead2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19e7dc6ac9683834ace71443f1d475927c85fe6ad85fd791f16c017f35de54b67f56bae5c083c38fe2cf63dc4a77b8fbf151583f6a4cc6b47ad634a327e967c0c5dd40c63a07b97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbf63dd4a4ecf82de50817e28d9511ea365b8685eff976e2b10c5972875d7b2d18f766b65e07ee7b1934ea955a9ffdcd77e43f5599f83cb3f0485596d66a5c53c9f03da3a8c37084;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h806cc0063a715f6957a75206a19a90751a674eddd4d8b07e8ceabcfeffddac496d8ad075a3f057e165c2ede3755f59d158864ac806c8d731abba4eb361e0229a729d15a4b22f1e53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18702e6380d2104e018fd1e5b6e4552ef82905e717640980a76d189793c6640877d2e52cafb1643f87c1dd1a5c4d89de04e0e30754d8e2ac8a36a3ad96062b157fda298362353dd5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a110554fa84ab6176cf2eddb6393f235838e3c6e5fe38d84a3623b2f8f5f2663edaf1215121effadc09c6f953ed22f0fea44120f66b4054fb2a2d075d7e10382e645afe9639ae25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he53169004e2387011130bba4bb78d80870c371bb9edd2e1c9eaf9c55120497ec7fdd7f1d5e29451dc0b2b65470b6df15b2b2f1ef2f0f422ee1677a67e35449816eaa8e61603dfbfd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3fa10ee443c3fb084d95d92a53aeadb065602129fbe5031e2d31f7afc828849fdf83566584e4c5e2e1cab9a1bad0e09fc8845f03c5e8d2c385eed54c72ebc14f7d312847a20d05e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d7452586cc29265607344b10abb6a5ab7ca0e0ca3880c9c523c6395d527a54c1daed5c5bddc080a9bf8043ce74729da228ade415f300656d09d27590451adf72c4f1ff6dfc55e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h483cf2bfc90281ed3cf81a19b1e2f92dae97307edaf3d2564de2995df91356cdc5821658af9def4e44a3c26c9cd235e4df045436cb29d1c73b89d95be3bbec6520106f7d2080cc62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47d2ab9164e7e209f6e4ea6aa789fb93db4a23b5e9c16ce666b83a0c89e7c4fc0a8ea99ff243a4912476eaf079c48a5443928ddf981f836f334cf0998f2ac6c76549d25563e1b38a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha70b4307f6f85e3580b6da04e9bbfdb7dcbe0cd220c3d60a1b3690b46da4c966e79bc05f7d424dcece4f59599f22b03c87b67af8ced386cd334a7ee9da4ce5412f89f6d73b7b01ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95abfb44f3c4ec5964e1c6e8cd5fba2540894d852a0aac1b8336563d0a37b0f5eac61ff1bbde860d423837ea700e8a8037ea1cd011a9902d0efd247d5ab36b3db5290b0044f913e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h746dfed3e00cdaf3cf5e73843a861b57690060b53bf852f814f63803c8fd590adb093a86cefdf8f555e97d5edff61112cf619b6924763641f02cca4374ea738ae3596faf73a32e3c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1a21f01c67a51a887118636da89e976c620de57e4e18d5eb9887f730e8d601824b538e1e9699c1af50e825acdccc7de5ec299c9a9a6d33b8446a924e08f013c25633ff99acffbd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3702acf4cde872978ed5a4fe9eb08fabc9b8fa6785eab1e98c7f3c865dc5fa8bbc6a4250b82b95042a9aa8cf7f3c48b9e4155394b9e1ca7ea6fee962463edbd063bd40b58549b1f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5da6ab23637ec143e4e5720d89064a67d3b4d63bb42111496289044919e290deb51315a87abba53e3e9ebd7b033f796682066b6ae72ccad18bebed4358928ea53389b4c10c6e767b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfb28271b71cba66f2268ea86891988ad0ebf89aa80afcb375e7992a742f13793c385f475f091a1f47b9b4f080d9ffe9034440d4e5ca069193c6292bd736265373b110ba130baeca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccab2de9be614a41d354c77a31991333cd5ec1cd48920fbb241491afb51f2ebe00bbdcf37ef757073f403b52ffb628b18f21452e9dc9183efa7b1ca7d08592bfd3ec43465fa16e43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h721362d2a0cabfd5e002690dbc55067fb080640900f4b6ed43472654912ad4db248fc72ef7bbbd6ac449889a85d857e708c6087cbb0b3279ea7839b491fbe2420fdd628911caf25b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b357e343ac9dd1a155c2f98ee55713ed6c4b6e4db4e5f1e51bac88b88bd80833c80ea933088483f20a945d07d8aa2560603b3e23013162f6d77b766bc35e70db5af5a31cf296197;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c157804ba1d0a90a7ed5b9d5726efb130fe33685b5fa76812ac056dbea565eb7c514738962aa597d0c28c1fda75e09c684647f64ba748e2d03def2bbd8736834a6b1e058414357f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8176cea4636156b17a438003077ffcd384b7977c726acb0f5604ad1b14652faf8f76783722665d8d54a1d5ff710a8c26f7a5a3d43f1de330c7ce462b90b751be8469a6e934a4cd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c663e21bf26225548ef789b74f3805366eafecd32cb881faef255378abf3f7ea452e0086756b9b8c0f32c0197985cd3439fc686cea3ea8cf759cac4c87092e801412410ce12f5cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b5e1664a46641140fc6e3ac91fe7f38dd8efcf6d9d8ba86f69715e08074e65aeec62ce0b8c7837eab7b79c70837757d7552c600d01974ed1b5b3f451a553d1de59a5741ef53ca9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7ffba8ad7b209b6a39a01371d3291d7da6c2656dbdf0ebb42692a15fd8ffc0010529c93cc66894a914d4ab6d43fc9ab753e4e19b054e93889878ae69f2fa685bf9f4a92782f2b96;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he41087a46ab3b306f731d30848c363849ee43d0d1d620f253515f5349b0e887f288ac8e9a806b300cb13607183f65c49bbaccf93e8688de33e1e598ec3bf7844075152b4b5e762ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h507c1806d890753e204bf4ba221b68e3a66be2d55b510db0f12d416fc9934cb3c19d67b8a02fe23b853c364d144f457a2192f73b8a0f25c497fc82c6faf24d79168b15ba12133970;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e12645ba893077c1988944495c62a7a1966ee0102ff453285041b9474e5e7d65e28e96f84d43756fdbb706c55640e77ea75b1ff90c6401f8ed9d0b44361765e0c3d7d405d3d9e55;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a438f6d0911a626a67da25b426ec6be09194b26ca369cfdf7479612cf67488178561ecad27d82fad7fa5fc81812f60337c5403ee8eb5eec6b2d6e1ca9a0338953c77ff484c31fa2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haba88d6eb800150bf84d2f2d71f5939445f21da6a9367b3ed03e83c4046abea041885994d78aba6109cc9726b09369daff0c7f15ccb5c76e7818551c80c8bb3b299951c618663a9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9416aa658216d6ea44f56a36c588893efff7de6e48fc37e538d25485bf4d28423d7a287fbd434946c6d2473eea379c88844ebd027f98aa6bd890cad2b03deabf5a0a931317d0317;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc97d6a0d48363296b3c64ee89ea9c0ae7a6a9ecd0a66d756b75873f99687db1097562cc4b6a6bc1e7f932ebac1e5f0c35bca45502b0d9ef4b0590b7814207bedacf5fadb1d1b4c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e93c0e7a8ea64081f2b046ee2ec59c8be58078c422b7396ccaf6e9f06ca626feeb5ce81412cbe2dc64be059a5a1ea948c2f8dc4504d29653b84e65bdee25c2a39e3d8a4e7463b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb8f201c8f4c3ea4578e9d15d7b43cc208b237759c5dba0877612878393d34b6cc2c161a6f16c721c42e5a1d3cf92e92ad48ec1983bb5610e60f515171b0437fb4a81a20fce4f411;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c15aa9fcafe3ce3293f24267649b7e5b921b7f939e8bec33a1dd08b6f7c40c68ad441cdc18a60a92045f7a452fcece994feb5e224e6aa69006a74a8364af8a7852e4f062552af26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0cbc7d42b04f1c98b04be3fa9caab7df08ca6d21cc21942ff30ad3ce8888f7aa8b3880903713a4b0bf05cf4efbd3f3b2e26c3a25f0ab1a0ae95bdfe55b6f34c3eafebc6bfb08a23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6033ab7a5c7669dd78b3cf506fb25f8f285d79e57b62b89686a3988412d698d6a4068e6d8eefe270700010ceac8c161c3a88fe8799dc85f778b5e397038634e4103a288e5a4e9ee0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc492cf6ce33bb6f5f2c892ec72dd04d93588574925892a370de781efcc92736ae43397db24ff0fcb49c37eedfab49aae6c4e1d35ff14072efb3627677e4583c9ba07e5893f45bf69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6b16ce8cf5944d6493a3aba52f4ac510b3641faed101bfa9b1f274807919feae3f989d618721734d85b23e20b755e5728d62b5fc3c343a0e5fed8c5c287b8c3682aa4cfdae042ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c62bc85acc7a6fdb8557efa321453bd588e7b73254ecd64b49f46705d8a64b03c524a28b9d53f93d0b35378e626a0f9d014eaad298f2c857b315c0842362608357859b17c37c5d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc48898c10622e77bcac0bac18ce8f6923e81b27c39e05de6a02aa4aef08e9b76a03c52806109d3e60a4347c6dd5e9e81fbc87efbd0416c746ad7296115415e61f90e41329d9b9765;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd03c822c048ff182d4fc5ea4698ddb2559ea1ca098a0df175a8840c9872dd105bd1094674ac0aecacef236ae4a9e434e9f2302928f3c8292137bd4ab9c5ee096554ef54b12da9000;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2139e1affab0e40e330da50ff72b90f58d0a91da8162047bcc54b9aced2ca3725c2aa6bc4e15b97397a8eac3c588062b03af7bbcaf278d2beae15f76db178c8fcc191b1fb95142e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e60a5c9df8ad37f9d9c75b448af0ada571cb708741bd279afa76dfe13ce81c318ecb85a1c31acde5f57ca00a3ccad0884c3c9ba7dc6b9d2cfc6ee2201e019fed88cef54032ca0aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haef9c9e5fae87024ea2adfd84690ee76bc23c728102079cf590e875e33751cd4f1cf98b73f93b46cc0bfffae89e76e77fe6d39239f43b95dc553087f13d27229c6a8752109821654;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2d703dc97cf555c5254cfeaf7f7a3fd3562e2332a943583d1b9142676f4c310cfdb3296b49857439ce50316166a16e5b407772d10703e6b58c265da3d918eba9a6bb0ad6a46f6b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea9ae6d3cd79881dc8f5dc4f4198daa52ae9844b820c48c846a236bf13127a3e784ce7a7fa5a53eed5bf3ff35b651eea40f02239d021097bf8c1cd9cb5cddebeb3b70b17ccb9125;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8df312d38d6e705a6e3d0c1226142610634ea0602adc1aa253bac08f676fed38cf1aa7b0299ace6aa50a338100cf81736985da6ab6842141165c1c9b340245f28e4ad5b57ad555f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43edc185284248d4590c1b450ef954aa51556e7ce1d1066731307456b7d99ac670e391e216c9a31beee59951d3d1e09b94cfdce51f38a08825eef0e9bfb4a9c45b41e451d8e27b90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefbcad955202007386d025c340d524d02ce8f8385cc279c85010e3944f340d0b4b96505ec37ee4e36c72881b3be26735c79568f6bb32fec02b2c9f41a1fa65b49b8b9a86ecd029e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5580e6de834280796729b79aa5fd118327b2afcc20603b6199958cd825f3c4b65ab981380de24475a8a9f5d08c96af046faa4250501b739a4db8e1be0a3016d8d9da3de5553f808;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15bdaee1a2940e963f9f80af6ba0f0587c8531f16dbcea44752b269910cf07490cc9582cf5ffd3a49a6a15ed0b938221fb951cd5f9cb1dae5b3845f0369ff1ed1d87dbcda42125f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13ba0a1c63cb31fd2f1de198e04ee97822770a4575e1dde931ecf972f9dc280c43558f3773769c2189637ee9b54f3b1be949a969fc5490fc214cfc164d8ea8560bd060e4f3ebeb68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3e77d0cfbc08d08d246a0026ecd975840d0c99c6e568554ad2d6ebb56a62a6a2430473248eb64f4490793d9877475f12e5fefe14d3a00cbb33fa982d48d6fb231396b15f07ba680;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f32cfbc62e651226bfc4174908dced870e0b796e5405bca6d38bee504341ad4062d30111dd504ed7cff9becca0c8bf8f06db7edaab58fca92ff1fb8694d700089f8ee97e9bcfd88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36198f079cdd9e9d849ee034f714725a37c6423f062f70a6d55a20e75d287ec2957525b183ad6bf610bf67453ab4d6b6b9d642f6be4960f60b536db51d4b90c41d5fcfed14a6d97e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf7bf7f406c484695cf507f51612f1e515a875cee104acacca6755f133ceb8f01f466289bd456c6b8d6f389e5727475f47dbcfdffb5c448501f5a64d975b45956e2a460b55f44824;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf323b0971bb34be61f61035f59f3a60b68f8d9db671879b10b2da6a4a1676b855b92b77e9617f5bc59f656eaffd5fb64f06490865cda757e229841e5c26e012fa48ed542307111b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee33decfff6bcb6af678e9bd6fe6296d835c7544831596d4689729d518514130fdf1ab51c9a53018c9652bc56a6268a3e48e84c1bfd04750d85107f343d861992e61514dd002e669;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d3fdeb9502d24d06e094b1cef6454bea70684fe0c27fb87f875968fd8bc7d75572a913c9561f3ab59a4749b1a809566e3899716090f91bda4d9be919ac4ba199fc8c837d44ce451;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a8493262052b6eeaed63704889bb55d0e594562527f684e8c014edf4d49cd1a1d51992310796c4770347cc2399c882b47af1900cb36db402da440d1c9f62cf6f8ecf64678f2a326;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd0fee8dc8dc5b7ac1131151b96209303a4e22c6e7fdef7272cb68dc7e2cb19abfcb9a490d30a0f2440a32a6c3e9cf0f1bcddb73f9c6848f41dc36d91bf2c5426da4f0464ce62587;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18c0d8d456666877fbb4193a0efcfb7114a83392b64a59d5ccf3b292ee0adb06b0250af3184ca980ef1ae5d6c42f6bdce449b6b470d11eaa976b1bc525c617fb835f8590df778fd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4630f8a32fd96fac230ccff855e59f9161049233604a805ac7ce66f7975c3b0f221448540089baa47700ae5a9f1dece9c5c20a09dc85e666461b2c2b8e73eb7a604120da507d12a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf22a188e2bfb656a972aeaef9bce9a03a712a923f0b4165522de1aed72a9270e63014efe5e9ac28a20efb3a3a9ae1cd472a4567b3b7c461c1fe7520cb7cfec38779c3e238e5237d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc6934606cb4c59f2e1021de6e547ab6231e9d2b50951163ff4a4bbb50b3c65414aae710a3fb158095ed6a01c4c4c627062899d1746954627d3e7903f6253cd22abf02af7d2b5f0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb685d0f00d9099a6f23b80851bce53f214363058131487a538a8721f9423d9b7a3657630709bc17ae615df0aa7ae21bee36fbb709ea8709e365a87ef31ca75366d83c2e873a8bcf1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h748e59ab8f7b9b9428dd7e8ae753b563e1f6a3a8f84edd52ba544aa9f303dbe5b0ae8cbac7c40378e174b76de9cd5f8c2155415e146d059d9a45883fef5af9c8ee43dd257da3f4e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f3373ffc2331bcf838cb220b938d16b03a52d711d05fb0ff72357c0cddbb6f583354f215afcad8c3e8ccd57387e1070728ae468eed942286a0aa2e088d483e9f12b421c1ec5df45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfea5b7df4ae10f80a3b926351d7d45f85467da3bbd690bc4812251454cc06bd79a5de3c695062bfeeebb2682cb63167dbde45b77b0bd56821986b944bc6bc4f72600dc5f21f9887d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab6a35e9abe811462497d3f1fce0f9b82e99548dc9067ffa20c536f156647c981913bba170a4677082a40d06d27281041cc07cbc2c73143a084f28405c302716dfc3fca0be94a014;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6b6a78779ab0f8915ed18564f863387a5b152b09b4b4f003caacbe3375f0dff95f7d07a0685d2e7507b0ac1178f519a0e01e5873bc6fb71f45f050a5fa9fde100deade35b0536f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25851d77678a1279e834eeae2aad90b94f9e47cbc5498eb55cf9139893dad911eca7fce1f0c56fc02589d456fa20bd2c53948eb023b3a50fa2d8b715e6d05728dd874844b9d17fc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8da7e7b81863912c9ee0f3a8694a5ba650b8636176fe3945ff369c1c31108bacadfb216b405b7ce094508ea381cbd2e5944a72d992e7ee5384f04089f4752e2c88c1e172db5379b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb57a7251d7431398399dcf8ff05ac2b40e99deb0cb7316c0a109ba2ee22451222ac0fb42c02b41bc885b1b0fa833fc0b6726690d573599912dda19a728cf8dea961327b795c871b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcafedc86a19bb0a5c18d9d3e30ba0b93c92ea986baeda420a44333da0ce1f6bba5aa89a51bf50cf2942da9e0f569c551b4653ca7369cd41728db09f86769c3df54e9387076da57bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43f7c6ef1a96dc85066e6c3acd63a81bae28ea2ccb34a8254aff42109c1644ff3f5abfb41efa5f63b118149ff099a542e15b4b1b9818db74393c6ff854ed5538443af067b2b5254f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48506e1dde6975869a43db3fca569424423a7cd717578c723d9ed85d66ea03a2fecdc95fae5c4999dde01671a2fd4a9f8f02694689234f251333cfb9dbcac5ab7fc83f32bcc4c714;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25ae971e632c1944b694174cc8b1311741c4ae5f652d260e0a0398fc0ea280c19b6c541add0c0f04006e9718c499128bb0d2cfe4619fc2c5129ceb2b6ebd06c7cc95e0ac496d8537;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef017ab59f9716013d588426144bffef4d768c75dc8008ec4b9d406bef96c13440274f89955cf3518ebef9565f4a2b8e1d9a6ec96cee9f673af81ce714520429432f27cedb066f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89a1c90b156c31d0a9081ad39257a9e97ee28fed3a58ce285cad63eca23307ecd02446dc90876006c9b690a88af9528207c1fb69f5dfe7e181633b5c5a07e97aa9a2c7f79f43ce3d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9282b157f7dc17b0f4aa7cb41fa256b0a4d942c0fdbe9edfaa56c3884f89eff3aa1565448ba47f5e88bd56e52e0c1475b5228b2d95269bd0ca900dfa6594a1cb22a990f0b1cffed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1774729e4a571dad29c12a88781a1a68a7baea7d6094d119c68c04d43b5a3e93ee0bf9f3977dbc96caa583d70aa724bed33fd7513a66882e5f6ccabebab44c90af1528258d8d35e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc77724d8562abc7ab564f34aa8faee30b546edd84b2e3e677104426e5842f18d01e45f12f988c5b50a7dafe1d9f806840c20b49e7ce24033e5b4e6ab08f8cb71bab82406bed499c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2ba5eecc6f6cd059219e41bf57060b65e7a0482c0051dc0badb8d0424acd92edf2d2c1746fabfa75aa16fe712f504c5621253fc2364e28020646a9c374049e65494ddec1ab65f95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd095e1337bc97624c6aaac3925f35a0bec1a3efe985f8ff465b3f2d964e5fa2f8fd526ecd85a56550a264ec8c30ef19e7ec05d85e013f0ce1766f8e9d5b7490d8947b3793d5f4741;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70908f8f59f6c99dea01e349feb2e52b696a2f2976e2987b9eba02cd24b3e5b74806994282d6506dcc90a860e9538ea6c4e611bf9de201c1301c5aed1a7bd88e54b32eb53259c126;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ee22ae8a073948f6bfbbb5cc3f979b7445b51c6c88e1a18bc3b0c6b7fb214cec8a81dd1a48ea895dba5d197e6e78807de893993488da603387984431651f735fddbeb390abdabc3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19e70132d52927c028fea3e7a3667cf13cdccc470b00fddbab0885c22caab96c17c171d82355874e33e6e2758a4b91cea4dba7262030f755e1d122f85255b2d84e70b6c2ea33fb54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h128e14844737b46bce69bfb119acc34af4c0a3825f31ab9a6f848e8394c7239a9459729ebb4b4462a52ee1380b91fcb11edc90f1b68d15daf40e9c560e5b352bd1fb9c8b2ad0bac4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1f72ea7868d80b29aec65165b9b64cd52050ed72e44ad1128f6deb4e6d99bac898c6c9b8138478de1316256546710d2359d4da15cafe7acecdfae43d26011992f85738bf8bd19a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h835e26653b05ddcbf741ea41a48e954c2b359ef3043817e4b1b269e59511fb0f27ded324a7eb321b2ca5d605bfd183e43357771808e09c7e94bb45bce6115787f0dcbf49057346ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77a013258d10d314733f68988faa1d842a1fa8a0e1a76bb8a862b3dbe6079c628af615fc42897cf84260c165dd98bbf265f89c9a1814398c65f2dd21f84394b887ac1056d1b301fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93036d4831b49b892a6a4fd3043b7e83c4a3b1449c61d8532a5ed5b03af267524e4ba078fc458d57f587aad9df350c31d079f19b345e9bd63048a0f2aa9135ee0ef0d5c5c3e5f73a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8ab752fc4f6858977cbb4f5fb093df40bc589b06c895839562649c13913c0021a9eda5d55d789ec3a489265e4893d2c44ebb3278c1e33e34633e3712c86775ced0236de14465459;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6f32816deab57fee7b1fd6b091eab2abdfe41979fba54c7f48dbca88cd4e41da5604704ef493a8e6e4ce0d6639e6e5f7d9939c23111bb7a900d063fcc21697f47797f750d9d5149;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc31c55f54a2b2d12a7eab3e626cccca012461631a8f1d3f25603f8a28ea4a57dcb5a89ff5826668b013b01fbcf457c6461eb869279b87e819ad0cc39d11f01fce236718bbe89e54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a73a55d9715c074e2eacdfda3c3b38540da95b4dc0b5670db431a1b556d494a3ab6b2bf2011f8e52c785e2f55a9f298f31fc3bb0faa0ab702e9b42b660d27fc2290c69915eaee28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f8ce8048e491cbc5e5d00c24c26d8e30586a80330deb3a13208c10db81141bf79da3b531863000f1bd5ff29bb63be988f9baa9a70a649cbaf2bf75e6fac421143f520f15fa567a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb51d5a958a745e234101c512d27066d34c9f0bec73cd8beef5f30941e0acfca8c98e6968aade51df7fcfc6552fc663445748fc6968a3971185df514705e03456126b9ce4a984ddf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49586ebb25cd6b22f3261b0abe649d6a2079fb879cf10f6d6a39ff9dcb6a713c76dafb929860a5ee6b2d38f60e5d055e3762852ee16db2e27c0aa29ab18b656a895bfed99f0e924e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24a48e880b7789d324e25c2b081eb1462a614633d124f6b6437af1a0f302d00617d9eb8619ebe02ee1ac39a8fb61c63fc2fc0c24245553b01e025588bbca006c5bd125bda5cd4350;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd49c3e0ff3ecffd95ef4770201383f9c551971a79392d9241ad266624a3c0b7b0b37c6c3d13f9d5bf9b255a87c4d878dca954429657690c0e93f79cdc89e2e1410c15190bf36cb24;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h993d2161ee55c717f9522331a5bfc28a491ad1e85568d7186ae835f6c49204b41a255662261f6a516ecd5d609d4b66ac0763f719cc4d22bab5040e471c79c2712db2951ab905642f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d2b7159082352cc2321b9b4ccbc5eed65ac40f880d9fc80a675ea7baa67cfc7c5cdb8d81ad0b9a5eb810e70f47a2e395f155e2bda3d932c39d617091dd82d955121d1afb237b3f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aa80cee1b43306b1db3b1ae9375e80b3be9f9564a2dc94f5d927c55d678db4868300b2f558d24683d429cd58296e21f04aadc95c79ce84ad57963af0db2b176a73ac1e25023fcc1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb28c466ba6bda64a449239b0f1b29418898741b1651023bc03ca36f395f26427edbbb874670887e7785f84e6a835b0bbe9590e33db9e12088c8a75babdfafa850a42ae02567a124e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2e3f53dd8c86a6611d1a13ef667b1455854eaa843ad1822435fb7b5e1538b7c28553e7bd6580c302ac4bf847d79feab8aaed1d50518002ec5c4581bd2ec1473927b035f1976d930;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68e65fc3dfe4c8f7c0691ff32438eaacb2716e960d838aff67f01a05e1bfcd35e27085110762b75a30e310786418922d9a6a015e2752c1aca1e461257696e3cdae8198c3c2f8e324;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a12bdddf4cc30d2238d4b5d184cee17415fa940955de803cfe5f8b07c4df78c43be2278bfb8992698f182e619b0b8778790bafeca59b39f41788bd60dc0b019403b81014332c633;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f63f134438a41a749ee5517a9d43fc02e61f652c421638efdac072c78ae58ec23ba3c05a6f2bc021d8bb66c638f75bb9239c41ab49cf07f6a0e1a859285b04591d0f975d0df4a04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cb4a8af044a8ab77f9279728200322cc6a23cd40f196c4cfc7f790215f4818b3275fbe43de578372de25b12c5e02836c6b05fbe5ab45bce5e292bef97b630f1b3e5cd5516f19f23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34edce4b73282dd1dba9de9e16b3a7e38a6d25f6920dcb566412500c2aca126228061cf1c9bac495e7c5bb1596a3638d5c4aacc5a3ef90db2aafba97cef017b22991d553d380ae8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc856986c4451eed8d4c9fe6d781e4198ba61ca1c8247e3464862ebb5ffda150811dd3556b5cb632cac6a88524aadd51415813a02de075605fce866becd32abecd87b4bab39c7821;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h993a1771837bb84d00b266eb454a5d01f6c78fe5ed459e17f9ecbaaa25bb278894c82d856260354cc26c19e0cf51cba47938c9bddfa46638a8255efc47d67e772c08e6e45aa510e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab48b5ebe336c2a22b39efa72fbb8e0d7edf8c7b5701c8b1f65b622c397627afb3c1c0da617718094cb3a5d20bbbffa226b7968552b83d675a87050a5c68f0f319504286fafa44b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dad01be71521435b1fe10af3b09f190bee2eeefdbeedd7469c005b37bc308b907e9e59775343a59ac6e1cf876a1f2ad63a96dca23d87d688144bd9b929bdb1a8df57637fbd37091;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cf3b8c40f43612f6a5b344cd7e54aff25cff7a21ac7f64e4511e331ff078c5b88c125efaf94044338df4092bf5c30d797146b9f53bd1461156df740620584aada2ac3df749900a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15c6e28638577c359ef2c66230945d58abac50d36f2eba3b03842ef637d22d805e999f20930786e8da6e22c7c0a520f7aef141ea40d413755c43be6fb19b9940e257ea3b9ab9077a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16da34b2bd8aa612e967f09b079dc4a0d4962267095240db75f1f0ac6ec283421ff2c859af7e70ff96792d034b8fbb22e5730d6adbd26c0d1c0e09b9610c99bd393a7c5b6aebf516;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c666ec7bf0e31246e31dea92cd3a5999cbda1bf40f7e70c1551b87d66a5acfdcd7b80108bebdbc009929967c51e35a36ca6350b607b34bd8948edfaf2de44dfc3161822acaf9841;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd827233240cf19ae9847e9cc2396621f893332bdfba05fde8724a916d8c28fb9a0bf9ba1165c79b711536028b8c63c451c21aacf19685bbcbd2760a9675eb2f424391bd9e5cebfb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68b53cff0710889537921fa868780dcd5af9e4d670455018bff12062f97a545a778b2b36b1ee03af390206ab1672764719c37eef6cc121822de5e2efd468b76db84486b37504b414;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d418e45cacece451bd930d80468a4aa56afe9b4659ea309accd067b7273abda3ff88a4f212d6c3631c5836130461564ee5718b98f98e4f60029fe5aed564084ea18273e9a15b541;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7ea887a09647d6ea489f47a3f5607bab6bf86668d77ee367901d83b92b805f47b55bb20adc5b9435296d6dfe8aff5455227956098116e7494dad8ad4b053db2906bff00be380cde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc11c7c37bad80d112af264736e102596b0bb38e5686629cf2ab0f659aa214ca3ce9287c8363817b1e0f666c3510521dafbc21520537d975a8a76195e8fb3d01cd243860e2b9269aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ebe5016bfb0ae1445608ab23e12d02c084785c19c2bf2dca39c49b1df0056ff020d31329690795f69fdac566bb0a7673f45b4fe0adf72da3a9275161a9e6c69cc810f4254dca781;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d06b0413652da489770eaef5f651475b6b448babbd1f600a80c8ac910fd76c0d5f8a456b8f96e6c7adcf24502669a649c3cb97efe60c970ba690ea6cb877a1d845c54d9be74deb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39be9f373fdee84bb1edcf597e60c14fdc49cb7a39142d7c1a29fe761d87d2e5e0f92745d93afbfe96dd3696440c7cf99bc579f2329f0d17b70d5fb2fbcdaceb6abbb313e7e43c6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a9104ff1126ab20388b4c1129eaef50e0819059b0cc4f7309dfedbfe8fd3be482e91883c209c31da2a839f991b848e721a4ce9c7ebf28e5b0eed97f704401b2dbcd2eb95285b313;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3387f0a7d72956d6362565150a06c1d2f115f4c210c3540cb24d40f8c5a557ad7ddfc1ba9a34001907640df2e22cdb450297cbab6e6b70295c6ea728458f504f83d581d8f3aa1f99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b681719a82153ab396536c610634111a222cdce77fd8f38fa16771f2645b560db8941720cf22f3ee6dd096d0c53b5bd0cc41a75899a4a94f1f673fa75d5e87db68d814ad7c4c685;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a83f0ad97fe2b4e88de0c516e5e6b0f1779e69b07c614182201bba0f9f8894ec20fb4ef36c4e51dc5cc470272ba2a4bc6b77944a0dc73ac5877571c2bb3a3e320d2a9a5a7c240b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd95b2c74b091efe06a2f1affb1283704eb86d734f22665f4d0d5d482f7bca984f64fc810497fa7cc3cea91dc9202a81bb83afb5db44a5bb1c0ca9c5291b1351cee7107dccbc89fef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf58ac42714b5ccb61809be49b31f1fa4650f2b5e2c54298e5399713eef85b44578b90ca3ffecf1f54f8962b4e92b53474d9d56a028d73b734ff6f01cd4efb59accc4c5b6b1fddb08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2ca18fa4951f2d7ffbe194273a5d01dc1b99de57820c9ce19be8a576115eb3bad9ffdd706db54d7d60042bf7002ab695ce593833272157e086520b3fbaa156ca712251826c33966;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1264e1ffc79c7ffc9f24697293eb50cdec9f683bd77bfa5ea77c49f69f40eb3259457b448aae2071a060cced6afd8b380a55d60c9ad8a8a4c5556851fe7c37c8036b11e8c577a0be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcac648cdcaa99bea1e42df82cb33144cb7f70563ddf630899b0e95a4fdb0f2eb712fe3d446600cedacf4edb1f5275db4f8c7a960416241f40711b2627a65419007d7dd786e81b91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3097aa88a15f77f94a0e27fb45f5a4f4dfac510ed720c4b94b65014056bcabc4fb0c867c563573181909a03eaeb4402e20f31825d8be5a2376a68e7d3946dbe8c93d59b6011f4a74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf02dec2f2de7a4878eab4ffdbc56c0c23659fa2bd4fa73a6e40392f1e220cc7ec7e8d64ad2b602d17e6c2491b5fdbd449f7484eaef85b8263c12e2cc7589f6ef14785b3eda724fec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h712c030fe5d01734dca9312d1159613024390accd6152657b4bcb01e34502638c7b1a91af8b8df328b7eff9f890acdec6e9b250f8a2176625b773817a1b19ea8069ce82f146e72ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8090e7026dadc45303ca46e6fdff1fdaae4a083948d446ac073de890b1c54a6f4b90072cecc6d4c812e4515d1371e38588dab25657bcd4475aaa82691d6a2e8f54c3259aa04f001;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33d3ee16246fb60b2a5b9a940209fc648b581d8f2941c7b3755f4d207c5d8a0b10817227af9c875ef455bf02392fe44b669adfde52de34f3c771a37fa2976f2aa1372cb3924a1123;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9f624202023a609b0c7737d839696cc34000eabb0c49698270e267f58ff71c2f4ff4635070a26f5ea3d5d7e0c3a6fedd6d770aab1fc1f12301e714130589e5e263a60c7c485a165;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d39aaea517a2c5fff7f7c802b80e223e398130ea9d37613e99e8808d03313ec115b9a8c4f62c412fcaf9b50fc53368afc1998d4e53331d995a99fc0cacd69b7a58e07eb6e4d252f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42394c6d6184985cdadca10f27a70de3bf7a1468f8fe865e0f1c5ba92e73e744dd7874c6b2458baf420de56ddcaa9ff2f3391065f1648f26153bfd651ee03896ad9d3ffc1e24cc49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd49105e6efc157d2c5add0a9d32d4d420d7784b9a803a35bff59898ebfe11aa0042f13b83295ba072dc5aafada5649006d055f1c2f509dad8c82a4d4acf46bea794b59858973a052;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5a2730839e0659ed077abc9cd9b90549d8a5ad0662d0722efd6a43e3d87e5ffabaaa0fbbfb19ce5702fb2e34a7b06fdffd77413302902d1b0dfbe309e1c26cb23b03076c54fda09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9004b8f2f231f7c944bdd29146b75b0743264f58a29043bff65883465f81150d34f24a23096f80098111266183297b60a868cc43bdc1b885694fade927aa5e1631d408245dea7991;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52fe92562f6b54c3f6c6bfb07bee78df6c6f95fa927b3204adb0e5dd820819d6a154b97648d3fa6612493804a29de6469d4934360c111f5741872ac650efe75963f4ad8ebc956f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h286693bbf41c6d9a3f14478e14f944c5788b928c5a04a67ca9e4dd6d1ccaa78195b76c61bb215495640e60967902b7f4f403ef270e1f17036c0ac2c07c7f4c337abdb00868239022;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c023578ceacde870fd8e6ba397ff5b42587d3d46340fcd8ef3cbcab751bd8483f55c4b32f9428335658282a31aa9d5b62c5ae7eab9b2d91063edfcc9721b46baac912a6d39f5b5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac418a8ccef11ba117eb20dd2ee4f53d866d4de4870599b18601bb005371fc6523fc95f2ce9085630fc9218a0480e8e5ac21b04fc99f6954f5b484c5e0768c676d04777077509370;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36eda6d1e9341b09cb6cbe220425ac63fa6dfdc3535720ecc2a4838017b2275e844a69cba7fbf9e860882c6b5be9ec0dfa3e6ba8ab1ad4b3208a0b76948a8679327f69b965cac06b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha391f2b37145790798c2da6bca38e4b31ad041245e3b0b1b3161c358ee132583ccc0dd50dbbb18d08514ad705e1ae49dc6f5a3b2cdbf50fa9520fdf94f7b6e14c100c46b6cc0f16a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he42e39c03f4c8b416947800dcc19fc35518e193d4471195b87a57ae7055bab91c901322f195303e09830f3b9acc58202d8430d2210d76ecf5c092cfb2047b2fb0b70c5f403b7665;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd092e208cdc7f6a7b053d62e9d07f7253cfe3248e060211eaf4433a8fc43629dcd41236df3393b06434c814696bbb86007514931fac521120eba0da138256f45b5a3133400bd4023;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he03def0c2e2a9e8132ca2cf7d795459a13bd6a6aecbaf7bbcf5882fea5fc4dff8fb088a399c51eaf36e7691ae19a87f958285c9d860f5d7eef460d24a9bffaab9222527fa33f40a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef4866b864b8b5a48f9d5734b1c4048c8a21292190c93d04f9252c45d2f6654b5b58f1c11dacd251746bee26b73f3b7ae09c41ad55b255f70930be800b95b95e099eaabe48cec35f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha26d6d871adbbc05d27342269068a6adc6f0e9ae2b8cdf1d89d50cf58c3ce5c7f319fbc2b72b7dab483e507c59fc6e8ff8f0daabfe8ca0e58d987f4933a60af52c6d6cb7fa062916;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68d408f56a37f817f21cf8fc01ac9a3f0897a9b0226af19ba13261f14f5af51b4739b53b363f53820da43732557f828f8de155fa7c70ab8b4d8235b9c4bc9314d96309b5c99cb130;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8774a0f6787b3bd15940e9c3be5654303a555b1922697597527d48bdad01a43c07114c7cbb322760e31cc2040ce7f30032fe22da11a5c735fe93d4d8dca53686149c8e44b01f881b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f714da862dc284707856a5fdc66df1c092b192c3d41115201f1da5d4fe3f2cf4f4e46ae5c72c3f7f4fc7b5e0dde258a3ef84b538fc4ccb507b62644d3355ea6fc2f64484a5c0834;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d73eca7c5e2850b04e4e7c9b284afa430856f5a81c444acd609fe37031a351c9b728f5225db2043615b5b8bec41c7b8decc3873faf01c8e3a3a6c4857b36ebe6f0b573896612564;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefa6112a5d5c9c9d69a2f2fea950692ce55d1a0b32a186a757c7fc1d37879f8aa40cc9eb7eb68243a57eb6d2feb8f28fd82e34baec5941d72c947eebef08ae20fca45bd9c46ae7e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7822448507904ca78919159fb3470f36200248adee477431d707647ed0be51f5570e93b55581abd1afbe21e6e5b31caed792924612f2d378304d1df6ea10b7dc9fddd6426d09583f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78af24c1a06d05dc6fdb322fa55ae8b57ad8bcbbde93df60d3031b69c71374597d5ce0797ee5853c498d2c088c1517473f5d08f4dc5584629cc856a06ed538e949091ed8dfea8df1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h811f0f27b10109957ce2d0f053c3cb3ed77a797cf6329cfa539813caa1c58e0216ac5d47608237eacd16c0a8bee150c2e88c35d2c36b97475572e2a2e993f9742b5d41ff9a801760;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6be00ce63a046ae6f5f4e8a36847539e22174661db423911a84ab9c9bd8b4284e2101321148b3a750d2157d61b801301237c3acd2c973997303d477733c4b939aa1e892fd2ca36a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10281dfa7231baf6961ef0f1bd0deaafa1ffb3ec443d003184b1348759696ca148cbc7916621a723c7340ba3d5ac04255fe2b5e901a34d0feeec2a20c6e28c729e035aa5b3c6bc8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h406f0eb8b19fcd62dfa6cb5ea98929cb3476c3c4b59fed120af5794683fd7cbc5a89f05e91d67c64cf2b7ac268d049e800580d38368ae94266fcd8442d7a1fd35703edd27a6be3c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf00b87b33c670c7c78cf1d608385ef84ab7535cf92ce98d7c98a11b803d80828489f2cad47dfe6a23a2536c632cfd441406859d6ba99be5eec634b607cbaf70f68b0dc886dd1713;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee96e35ded0a632453ed49409cfaa6f423130b631938dd109d86dc1541a6ca11d0ad26ff2a7031a9b01ed4ffcfbadad3ffb0a48729c85b0993f120468f8f2406095dd0bc535b850;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7ce72b249103533357138fc23cb3e6f29607a4eb21fada37028b9bcb43b13016559b03af138353887094d14dfbfbd4284553101e34d66f88918cc361af7d2881751e83853ea3ecd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ce20ed3cc5df65306afe03bea7068175bd429383d14024754f89125c9a6f69f2b56cec0c92f7e57be48e2fef519f60d48ee6fb5fd406050b67c95fbf21d643046e2d31ba0a61c9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb07bb38c24c329e615929b1a35d36bf584b3dee113ddcf82061f364a96525306cf68cb81929ea39bebad12e4f13153b0f7e9adfef7a5b267dc14378ea2b2f2dda01d936e1ec74c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69edaa94fd01b5c843e8636add810e79b58d4ac978a067751148a999e198c0358ada2827809f6b93c3c954f070fef4772672072ec888ccc63644edce498b151b2b623ef60b5c9030;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27880362ae69ff09066e74984d6833f4442fe11deaa9625ca861a53107802f6c4c461468c6f1220867d2ad301aabf0276939c9233e69c5d57e1ab9b8f018d958efd1f38007c9a8fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d9f5820af9b4f5f480668a96bdbd21ba4faeddc60a41c0bc15cc6fad04769f0b29c78bef3c111c363c385ae6a187e52004b99055a1ab1609a00a867f2aad164ca8866951740d70e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80c2934672034441a81f7eafefe1979042a80cf7a9d295be84895a9645e28846fcddbebff4dd3c2d618256a479f1ebd53ef2166061b9256f548b8a988695b8a47b43157d31ab1b52;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h671249772da2a085d0e4ed268fae6d25445c5bccb03db5df0f9cd44e96aa017b87df032d03de63c71dc1883abf6fbd1e6c2c41b298dc725d1582a94fe5daab87d5c7a35cdd733007;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h335a9ffa28da1539b996b18e600e93854a50b6e97fefcf08cf173f939583f31789847599a87888dd93533147eda2ecee6ba1b60e4c72198ce6f49c000c20b2ef765f4e7ed67c93e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3720940d6e8419be8dd9ddced4acb5ceb61dd04536558bfc30dbaa904e422a0d40d15aa132b1131c7c0e8e2b9c8ad1959d4b96637b7e455bf21f8d7b93906f22dd48cc6d0d2dad8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ceccf105cb720d18ddb2e319fc13dc4f6117b5376ada85df041ab9dc4fa5b9bb8e56a5446a0751784de014d72c7d3bcedfa59c3c3c16c4d408b37d3c9c7fb2e3df3aa216fc95f6d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f87219a1b1d82525203f1cd4a5fb16a71f90f5590263e51221b13cb8084338b8fefe06872971f1cf2b7d9fad8ed64169ea4caa6add9580aa378d5beafe8f7adc2c715bff9a00acf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29aebbf97de376bc8d7e8e4f2d87209fdac3ea207ad4cd559b20ae394c91262fb3d33cc33a864a3647edd2f41d40e829d5d3b785af3f30cffdf7d3829e14f118b7d0c1bdc059e4c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c0c40daac0ae47e738de99390fdf7b5b4d4e618d2d3c44276a12f569a6c61db95f25e34082f7cff905773ead9a21e5bcd67e6bc137b9ad7991692a2def40da9630d292f2c733f79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bc654cc179ff039a5ed0342276e6cfdb4b098e8600163504d6686bcc2427ed3a317c5e31edb22fd8eb23e748480044cbbd09c135cf140c72f43821a8666c2558471c6f1467ce73f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h507453523466c48a6067ea843dd9ab5a9d015bc147699ce475a4fbb7d657e8cd7ddf559da1c0f21297e3fd202c3abec7ae192a9f1683af16db3e4d11e4da844b312052f4696e60f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88a7d01b61960d278b3fe4047c7b0d11dd563d194c5755e584dd558e900cc9e22c38da51f877fd1a8a6fd739eec8145d1a0d7d82f00f0140b995f60ab2dc8414ba203d0d1133adef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86c83af9b17ab392292bd4d93ef2f144fc392c45eabf04e994b966b343ca392c26c9b56440f1fcae3c3376df5fd3c6796e3e2665d010e1446acacbc55da53fe12f838f4dcc8513e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93c370f6cffd6846fedf0144ff0b2c55c8e47ffed5c59a5899dfa1156df54a02b6f44ea25c88caa54ae08bfdd65bc5e3a180804041b712154313081e271b7d2615d30257afb521d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa9edc16e29835ec725c63cabd9850f1bab566b257b6ec2009bbd0df020f9de3c8a60d2da5739120a8a3d6334e8ff98187c8485e467415f976761aa3fb8a74dd64a6f8c7b3233623;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha932077025cb9d3739a079f725cf33d307c23f4559057517672e3ef5045cc4f3425b127120fe135d48288c9fe7fd2cc507c135e978ba8c7ff5e61581650909a45cd388cfe6f22a65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16e27c09b2095f1a0dc10cbb8bd3510ffe4ab86cda4cdf8af1ff2655210aa0749e7d0415a1514b7bca2db8dce4ed918b858f3a4a74435e1bc809eafa4d28e852afd2d7b5b5acfcf1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha20a053059c6e47a6458135e4ab4dff0227ce25ff0a58fd77dfa23cface4d6ce172f3736a7414b21edcec72646d50031349e90a147d5552695e0621aabb784e9b0ec41c23aa48e05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3307332152ee6c2f69f51c368bc258dba79869804b4f9cd7cef612aca2a3849afba88d229b245a14424e4f4511412fce9e377d1dba957898698926fb6b8f692ff7449ba26fb1fdaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h204541462999bc36da909a709def10a9e7a0785b2221b80bdc84ba772739b2b245222aeb77f93a42b07ec3339df665feac7c71e2eb49c0811707c2006c9e86434dd93fe55742abf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb28aabe82ac022896392ca27e2b5a2854eca4c4de1866a7c40069f786828f01ea798087a93ef621d3058deef249910f0bae84b445301c002ee6da4f17d491a6af14350fce2b4753e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2880229ba281f4dd00b95254aa5aca4f9c92e2be5994682fa8fac8eea082c62fa508806f0d4fb25fc817e5cf9e7ec9d5a90f5c652c5889a204329619231f4cc54502e5ca41ada72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h999f788f97544b3940e992564b05e844f0eb7b3e1f3b1ef1c046e0e58699149dd65a0e52868e7454e07c8004f1aa91a3c3bd69884512c5948797b6f122b561b0f9825bdb5e0a7ab5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3eae89e9a4bbe9c0ae808e8bfccb3e9322df929030ccdce56477ff35f856a12823017960aa9000041c15797ed4ba9aee9221acfddbaf4a38bdc1b506914e45becd6fadc595bc545;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d09ead29d8a16f1c9e57ce28d251267476e60f5cd22345b87c2780a48d35a7b7a2e07a1fd23fd7071029c5c71c65c62b12d3bee9f309824e176cf10ba78b7704154fa53479a0534;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h315e26d4ba2a11da860a1532b15927e005417f792f092c072138f869a0ee03feeed9589f9d35989f469f1b46de43e9761abf70288c89fb15c51a39003d0c56fb1cf913258b8555e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h637e8e8156147bab3f98a79680674e111bd70ef91059c28ba41a312f1c2a27990bccb78cd7f5f590a775ab59b2b994a66bc5e1ff5955d36281bf3025fc86924694b95847baa4dbc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc859babf6ae2bc1de9010103e477dee0f76ab3f5c06700ccd0a033a3d14d1eefdb4611f4389a0390086c67026e90b0da838cf7bda271a5facfaf2cba40ab4b22a3a52166b1487a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84258f654f0741e70752c80bfed3eecfddbb4381cbb36d7b22bbe04dff3422e1bd855ec4a827c6e736f8a762617e7b8435a66094ac581adba407c50e4c7d196fa67cc5a6057bf5e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33fac4cb83aa3398ed6123f7356b48fec1e5fa1272b504ada83d6673c73551f6bde8af2404aa8d46bacf5efdfb35af359edb63f6428018c6bf9c0489d9ef27243bc75d5910130166;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb663b495b30c1d6d666e68f41929afe75279999f7f2c03ba41a2b74cb45d4597803b00798532b950d1ec41b36d7abf1ac6c68f2577d8deecf06424c779672ddd6d53cd3aa863a0b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c8caef68f1fca18c2f0c1bca329c4abbcda301d88d88cd8679ab960c528f6a22ba60a0285cc4b34a8aacc72d556bd27ac52b39be30f24ea11a488665e3e93bef83bab060feb735a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ac119bc0df2acb082d927968e4bc3c0580ebf9efca5245fd573eb6df897756911d7db307b818e29c2a3bec2508629b2fae28a0ebfe2219676c9656931d31ffec2d88452c007f2cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fb76adc7b8f9b8c43ed780dceefc08c44561e188c5299ae7ccc71009110b47a70dc34f4feae7d4f6a9c5ca20d533ca8556ae1f7ae8c52a4f5546cc7c42d068428b68922d28c611c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65566f5429fda99d23104a89a82cc3a267dda08c918efbb25f84648d06be299e4052612a2b92ad19fce1d78892e9150b743e3e995ffb514330d4df94a361e904cf8653cde795c13a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc79ffce9397b30f9596e3ea4a478c7cd5de9b29d7c4a0827dfe2646f6d7e50b82a85548d89b2d93e8c0bb76752ebfa271cefd6277bba39aaaf64a924546dff6eb1c74e3b1c6f6743;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd8d098b90a6e458eda7f60c3dc75fc0ba2e5b83edb8eaed21f2a5ac15447607535c9f0af2d467566599524a8f05cbe9830f4ffae1d2c0ab33b6d2bd1e383d1d58cd40e45cda03e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h145da539a3e5598382212652297731a3773c2b88b926f43997d1dbc3e11b029eed274f1d5bf8f6fb3b5c98b2731a366564cd71b45d461a186b11d4de438d82c5a0ca78d939364996;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a05965b2e25c35fe029e65363acef6006be0f0300431cfb8f870588968cb5ec6e60a59c0fb6abad625ca22670971e981054b68d447eff94dfe2f735d0e0e853fa1dbca3752f3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcd8e00955722659daadb1bde0b373f5b7f3008c3e05f3fc484125c9467b395199e4a19d2f9b2b6f40c77dd0bffd5462bdd42b09a23759d2b630ae1451422d7d7acd3927eaf5904f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb955690a9c96908a6c3bd1a164b359751b2bfca9a1d95aa91c5fc9b597dd259c0ea465c56484e041589bc4cc332f2875c2fae9ad603cf286df9b108c1e27ad1d9c7c415c885e2311;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee447ba5e71a36633b662325ce26084016ed8310d6ceeacc060aa58728023e8315ced48146c7afa670f0c59016916664968bf50eca020e2a03cd849d3e5c9a4f1a907ecfe8d9c93c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9776db9a8598bb1198495d57f8ab7364430a9fb8b9a6ab2cd3e9037ad99afd95a3e9921e70a5e1805283ad10e066c7889228e07d9a36542ab72acb6b05f2a0cd4b42f01f137e9bd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d8b1aa6aec20c585a3004876156dacdd444d0150c53c9ecd34e68507085c0f989a609205f3b1f524cf1a78e0177e99d3f1a9f0db719308ed3482ecd7bfa709d14cbb97ddab81e7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha94afdcec6a6485dc9dce5431a15681693eea7fa5c5a5458f70b9d0dc2db93346b548195af8408912124e650cb221ab685f95e42f1b5f52abee789ede8b18e031ef198ce55c06fa7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f8afb6e94a8abde84d45e79f63426db868b447f7c141199ec339d5d8866942341c250a1acdaf7b3f3337167a7af9fc18b7e5d782e50af6f8945cdb865a0691eab7d2472fe38b196;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc928aa84c2169eb031a92122dd3d07e08a181091887d4eef8e8958c2db359bc663f746ecc41431b3011f406516dfab6e09e15599894a0721561fd935ea79effa887af04d8328042b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e719c7963c83324bc05ea421d6d867c5bed860e817b3746eda94f1f9f1626fba0d261f3f917dabd1966abef05627f08a099cb79984cd607834660c24b2e2b69b9b6a914e1ad6bf3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3166e1a20ee518c16878ea4c86848a641ec781b8c6d38ea7f2753c2b558b9ce6d2c1205036045cd27b6f3a2b07e235ec52702d0830547c66c41703f0094799d5649698013cb3715b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ae426ca38f8c174ddaa377fb6cf3732c6d30d98865f3227b6ae5c65b1be2a7e75720924f521ce56126be16db69c5560add3bf60c7f0a177faf4bdecc8834eeb6c3cf3887b5826eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h183f434fda4b2d2797794740a6071113c5503558812aebe3805a9eb972ca67a6e9cd35728eb339270e815bc63ba3d217a9094b9943244a03db958f8f811242812ba053292e5d5e9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc19fad1bd1c8ad400442014a95494829240405fed05e94aa919707683f0f0bfbf33dc06b3d7975437df2f151b6ca68df864a28dc34f636bebf99f21c7448fb7eb7c839f0632c8e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd35b0fa79291afe47084399ada646c8f25baaad96f9ef454d269de86b9f70f642a0c132ddb3a301c474f1c579d2882102a7229241a2a29e5bdbefa1b03699b77341e7213243a0cc5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7efda3e82a7944f4dc635614b050d3f9060629d29806fd3c94ad266170c9d80599b112d63d002aacc0aceaf96536469a6d9b5e23c0d58b8f2d69d9034f399ddafcc5358a2567d76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ef37af051ab8c0fcf25e1658845677740d32b18a0a31d9d6d638110176ee7e21e6196777f71a49e971f3b24be6a664994447e2d1e4493815e8a95ca0c9857416eef9254e189d3a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2e37838febff516774bee285d4d7d1bb07793d42fad58f9a5f2a4ebbc82e585dd2d583f1c93b38246c90d5b26ab87f05ee0515bda0eb788ffdf9555d3a8e7368eb61d9119d10631;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e6ca73146d7db2d2bb25e423494ab184693fe20d57049924d195ee4a422b3429cbd968321e0c407f1203c26eb5fe7165c48f11fe164c98651f5a007ff547e317962b6ea34e14cdf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he80a83ed993d4e3928835b1978b7fdb345ce040f2f725caedc91c631dee0fa4847423d2c9df77a658bc078eee5df13dc812288e1c3f6c355fc28cf3d9bd767129079a248a9497e0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h604511412e80155c39fa7bfd1082a8db3e736ad1945c6dbbe9acbbf3f0be92c8181169a0f91cdd47c4d91e5cd8925f10987c05ce884a0890d509e1cb922e4d1f3bc1be2f615f30fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2d2b76c1cce9f9d92c05c331da3386c4a3733caf7845a0d58730b58cbc5252b52c4cb3cec2f2f392e14859cc2b56ccacbb6c48933dfc3d94d145b792c8992c0f1cf2721a75309f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha01a80a24c6b1ddaf0279e60b9fd21faa1841fa951f03b658a0de50fe0b4009bb8747b1ec1c1f4c8873f0683ceb281f2b511209be5d2424547a3e21347bec0f8f4d4cc3293fe6f39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d389fb390f4cb4f77ad034d940d49d421fc4efb2af9f5aa6b9e765b473fd3123251c20b4724253500f41d973d3e372cac4f9f3c3967bd4fb5abae4dfe0e8ef5f517973c168f8a36;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h870da14456da9ac1894cef1142cbf04a29abcbd6aa01f9cc7c26e911ae70e3eecc0bdc6f61f9e77b9af6dbaf7ecbfe467550893505a5410c08fd9d88b11bc2ba8428c51cb4fc62b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h433027364c706a88ada7e62b501f3f51d3b49c1ec7679fa72a3c8592f4fa165cda6d8d1127d61d37cda43eb1ba959f8a20dfc856ea8e91166ad8b8254a347a0195bf9615fdd302a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45c52493ea946e1c3b3c1a034f60cb6ad3ccd54e6b3005fbf52d1b41006e0ce192466dd8352c40a13726dce82499a498d858be431b8a4a31edbe2ab148361511ad6234dfd7321ee7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5adf70f6d6288440f399049cca5046daa56c6bb8678342fdf3cd48f2ec8cb7f03e0bf1da3a4b8e2ea2e60c726efc23e3cd5f3131c6563f63a6804e1fc7f5baed6adea5acc7be44c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a47bd566ee259a9a4063f4495a367ff8bc250aa9ca91541489c92b98df8cfd2eba913ab3160ac6e2b96e443b07227f4ce313f4db94ff747dd2ada531b293a565d114c41c175989b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5afad6c78d2935b59627bd189cc3dd9f3a31fc4cbf8c1587704a5fdd059f1f9995be4f8bbf7faa7db6a5015efb26b5910ac496b6ed7b4af279c54e3b28c84ace1b8d83ec893301e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e62c72ebe6d4aa2ec96ce7fe2cba93339ee022c877a58c83d9fbe58ee91330f15b7bc6b4fa9a872f45f4b3d55d8480107321d7b59ff8373cddb0388c0848a0f755fabf065d0856c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7966347c1d7103889fe491f2ef5a03763f428aee49bdf7d3ccc01caa83d86f9f79c8fc625ad1a1e559a866c393060cffbd1757a73c982877d1e6f89789034db43cce2abe66629d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha25a6fbf96cbeafe98f08d1aed2ece56572d431f765c9646dd977ee08f065584308b0ffe77b9d0a03895dd8b9311cd4df3e89a93c6d500c05acdcf8caf5b7e5ccd7933d4f6148b03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ac721a044d8d8b4bfd5cc1a6721c8fac43cb42db65224b64cdd2052d540ca54d299d21ad56ea32b5b604d2c82a3d26edac742608f2e6ca21de381fdcb7cd4c64fdf0f7d34171d98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb88ea206b2dbabe478a6fb40ec0136f377076be7913716fe5c8f7b5561f1b069e5e0c9cf8827e518506b442289f93814960f4b3c85cfcf1206ccea2c72d2f78067a458a970d72947;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb036c387b1307f4d5dbc871a04f972f3f35678c1db612fb0c0832e5e9f9703d76cf2f1725efb5cc2b7076d55c960d0b1230721579034baf1cd64af06b9f6f147ecf6c965fc210bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c8ff523f9227552439915c8446670fbceb496c31a80ff855a7e7a96ac73b459b273f0a1fb4b504ee7b25f50f54c16258d363a448be0b36e760dca77af106b1369b9c0de95ce0895;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd9c3b0e15dd8882552e84646f4853cd93fd2de365db987bde64960e569fc253b426cef97c1b07d7c3a63d49931483c00b264990526e2f0bea348325137a856e83f5c470a7285a30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f95ddaaf206a107ce577cf4d5e5673d8a460322a83ff56dd109a7e805c30eac1ad94723c4d43176cb8a5479632515f94960ece5245944da9d2b32083abd0a88787d73103891689c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he07bb8b43cb56a3bbe36e5f3c12344251ed8907bdd6f64a1828eed06827e5fec5fae4a01d7f1e71c80a9a7868cfa7e2e8594474ce0fdcc636acb26d6ab4d151579ba24661c4c1e6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27fe7589de131f53e6958602b56c205dd4b6ed680dd8cb1130fc48ab4a4a097e4f70df49bc112cbd855c76eaddc8739b8a918334ec375285bc19ce18fbf321ca0a67cbbace0d1d67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39863204a4958d2c2b8969830538a0855df04347b13568ed99ab770d02ed582ca2174666d8e376a67253520f212bc5df37c166bfad6728fcf2ae9272ddd8f6a583245222514de40e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc1d7a0574a641b32cd5a4b49d2fba40207e00cde9faed47902dcfa7055cb987b315af14005ef704887308ccf4045b540ae0abfb0f4a93f23f69e4e06d19db60d0fb00780dfba47e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14a9f6aff4c6a178546ce1dae2ba94e0f8cef2439902bf543fe30b6a2a66aa93ec36cb8f8bd16ae5ea8082bd8a250a085f5f834b314f29676442cd788f2445ac944abc5604e00c43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4e14df86f58756071ebdef40816e571fc41437f4050a491158669a2f79bdcf007bb0d66dde1863ddce78f170a27e25a8900d2ef083347d50f51df5ac65cdbd41b93bdd8c4e81ae2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17079f21ec9bf213ff519cdf4b2d1d0a4e60963e5e17e64dbe53016d7518a46e28f5c252304ff47a98dc291b667e4b52043d548d5d9d869660e70072cb7c7a537f0e048e00f39dca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h988b741ceecfbffff745dd028f1f3e63974334f6a0a5ce261f118b7fc4d4bc71013b882f21122941ef6649adb9513fb89b9e9bd6d422abaee0b509c16b56f8b6560e75b2e6ba14ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2aefd83d071e19993f9eaaad54c2ba39b5117d28e143e55d6add3dfb78d8fe29f4e8de32b8eb9613b69d9e98213cd5ed0f0ea3caf0db1574b33f1b94f00d75a03f56538a34776db4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h539704d0727727220253ee91ab2d9b0b2e819ce121fdb67ae1360a69c0a0d353d4b5b52cb9a250d856d1d17dddb1178978471b53585156bf69b4ee2643c29b33d503577a4ba9f30c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ce0178a688a4a988cc07c2880fc327444a3e9d4c4751718a92f3dd45b9eb4f01d163e1f5bccc969099777b3e6844f8388e82961725afd92f72c330fb6f613a74cf25d17d0a919e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef30c6c1212a449aad37561ebfde3e74aa9298b1dd9682b8d5c9286b3a96bfc0ba6493cb0b884942035539029beeda5536c768aaf13e555717c9de6a4dcbadb567541819e65d0228;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf085e7389d960f799b33b2628ada62e1c9cdef597721ff97a4d879bf0131c2603a5a5f9cf941ec0cfe0119ca6c4392fadc1a0279b78e727896af9a5a446e2ab71227b048126fba3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7aeb35d8cdc85db2fd88cac2a621a2e454c0a8a1844ce2a8833b8b8b6a5e485fdab66f4ab8d3d40b8375892303a4b90b748a796198741fbf78bfab71e0837de4b4d73217ff8eff70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6042978d7b6e07cb283bf580b20b506e2baaf2a07b1eecf63a15bf008242994a39c849c50c4f3d95fad97dfaf3b8f419040ae288a32b3cd80f4296f524bcd4c8fc6bf028e768e2a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec73891f5fe6abf32cff246c90227b5ca8ea5fb9442f066ce04c5f148af358a1a67752160c4c74d70e61023c8d1d2afe54d2751f57cedfd4f0a1a094b5d170bd96c9727f05dc0914;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f912e8b2ca201114ab22bafab2d0a67c1a65b0b059148a99095c742327f06edaa94b905eee07003e8901356c961b1b1d49b991039c81b25eb50b305d91a139e0e2cdf12813c48c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h659028aaeb7c040e455d799ce3687ee96809cb8b1c5d6adc9adc3f36fb71f134ea15b2e21e20d308ee76b56543f2abc7559b6dd5333d54b5b67bc5d5bd50ee959c80bdedc5a16241;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7938dabd24ff104726848f5a656ad3a62cc069563204a8768eba17d055111ec0380e7884e4dc10a58fa065889ea54deadf9c93ae81efbe50e5aee5e9cab8715b149bdedb7dde5ccd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h632868e338d15421c9a7ccda2226aac48df5e54a2fa0acecf225b4e07df3915a8d6022ae984c21835da8a7a96c7848f019f7b29e2e0c79615e7bba956a32d427b3671e50213c631;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9737485b1fc6d4158fa9d36821fa62aebef5d3c3fde447ee5614e4b3cfdea0be896a9a0ae6f9dceefd19305c7d860f17177bd817ca7b41afd91122088f4e47bb7391621ae716baf9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26419e476c9cf1aeba6c0d509646a2b98366c4fc67feaa0d9472ea67d29c393c35c7c78b432dd40e02aee736d505d2a3cf77c4fa3fab75a79a5ea29ecbb4ddfe080de5d279982150;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h655b91e31d26ec1b8f4ec20c90f5a65eb51f814dff60c83936bd83d298c4d27cbaa772ce4cb6b05afcbe2e6a2f35912ccf40002f7894a72469b63df68b0706a7377d6b4955f86ef5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79c9989410cc1784ed6bf65dd8fe35e6c389c21e8de349f16af0a3f9a24c5b6361e5ba66a23624ed4eb33a87e3d17b4dce91c06ab08d9d094ff4bbe7275f6d682fab275408c76af8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h749102878f3ac66a9edc2b6391c0c7432b99570451ec4a7080a7c8300bb2f72264bc88ce72983b17cbe9f50637b77e5abf9384f3e5710fc2872d17cef94c021de304d66644a0dbc5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he23178323b7292378b937b59e8d22c458abaa2a01eb31876f5e337884af4c7a84e53bdcb14b3e1666763611afac8fb3e31a75d76ce5f51e3ed128418beb63f8c20503683d5d272da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58b98f989f68a142cde5ef3be75b68576fb2a5ab8ea19ddf8aae1fd55b513c542cf45f5fc842e2d4573f5e4b5e73caa732f56db67491440464cae889cbe90776999176c62d3b99ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c3b840f2dd4769e47f00360bb5e861484d5c28d66daa29192c3cc1c6bc5ed40a7813450fcd922a6499b11bad846d968a5ab2f627d0e53bd2a878d6c96d25a4e179574114d385590;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f0ebd0b61303bba26f4d8c8b420329d1d6e631767082a848d7fea8a090b1c836947130005d204eea64587584578a139ad38e52b7fe670e3340cd19e2a92274b3274c51b809c1f41;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ee1801afb38294b2176d23637b1dfbac871eade6c9bcae02a433d7404c209a19a27a578f11e016905160b3eb1dbd1a48685b977c06240ef1212f2aa58680f2ccff90f801adfd451;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h971abe33563550490e02400b59ce97cc3bf130168c0f9a7b94c51b880f8f6e7be59baae61450e60c235f6dc4af812878c9a2780e3b4a205d4bf5dbcd1237700ecc32c59690906fe3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bb81a0d29e9e18f6576994099d3c65b16e79e06683c7a49c3277af13f2b48e726f93e2e0b394f8fa23764a9185f82cb320bfc6b7893a106f1d5af1fda8b62fa888ee7a63c7c03f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc134c4428ad34153d9666136fc5cc903c7ff3c67f149c270ad14dcbf2b338c24599b6801eda05b5e20cd7cc18a4aed09fe1a66447cfcaf4d05c2c86bf60bb0a9ec24118c82f10231;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haea5fa1b1073b2457b4b71f21244c4f4b50891158bbcfd7fb5dd893766c40da61ffdf20b5a82f8c7f013878c9cd26cbbcc603606664508de21dd66839e361906c5b52eb9e8463723;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he504ea4fd2a414eda32940e201f0f490579f44e574c4a00cfae4b3beddd2703bb9df768ed0d80ebca7b6663e7ef25167b0873e5d92a468435807b32de5b8a376377b6af1020ee8ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9022edd941d22fd38c7f14740f18df995dbbf78ccba17ff86d8354673a47ab5b259dafde792337f6406e48bbe5b40e1d1bb542136a36bdf5947fd775812bb02a31a72f5414c5b3dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ed1d3805a4d664dd184ff0628b4ca794a4d684f4d6357eefb331037cad095c2fb14aa94326c0bd5fff1cb4409345ae10752e0d67a3df52fb65695337f707efe2bea21f680be32cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h312bb45b267f34e0bea4d63618159c45359e5a5989fd6578bbe8b93afbfc17f9c146edf6764ec9255e32e6fa3a9583e146154a2740d28894b23a5566929d9aec5b0ed140b043cf23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haac8045cd7fa578a81af5b8da3e65795464f1cdb330730324907fa5c57582ad72fbc6a92e2f92fd083701c75866f97d83da687c325dfc72c17ae6c44068f487e620934a1526e07ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f4a44695eee0d8c72a84f4ffbfa5cc1de4c85a6c9183aec5f37559c334aa41825323ea4296894e50157bc0d2dfe67b650624c36a4789e99ca4bcf68f1a9a09bf4b2361170493426;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h911cf0c7cdd46b92d0b88adf0d30b6bfa8b56c924692b7cee498769d75d071ef274efc07a4d33a40a20c57a1c2eb46a98bc81993eaba8d2872cd2587c55f138ab522038d14d2ca4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf12fddfb01a4f6b92449a3d978d0114dea6ab8d1534c75f16c48e008c3202c619530f618d46f48caccaf422b992219c3a9403b91b7a058d9fbea98fa3fa816e2c453f0c3f69a6a8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc12fc39567fb7a158f94f71f0933289019960f2b0cbf8d934086a4f1a831fd06212aacf04e2b7122e20dc5b3f1ba83b00caccc74ba6336a8d36473d28751990b812ad01e799209a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24b584c70650fd230a398280eb9bb2968a07a9b2202ceece23c2d8281a4374c21a230595f0d7f608a920eb9fa388a00d01a4d8d271b991d095166a188716321280be96769284ddc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18300fc5e8485aa2aa69662002566c4d1a11ed9d6828355f2c5d794bfaf33f346606ca570ac5db880bbfbea5d986b76797fa19b12b85ab46bc16ad3758c9a94b2e66ac26a20c87d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e9ff8827f4fbb66a79d0ea8962cd91a91029bfc54a9f5028b333765784f519e9193ea081a6bb52dda3bf58f2295429161c4a0804afd1f51105884fedb4c3bc38d8e8d0a6aa1b211;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6778cd3d78b82073029ca175de5b9e7b3ee5d18e08ef683fdb8ff4b1f48de8f7637a493cab9ba9607cf69e259d7d7bffa7da784d4306c109e8eb30a364ee2780b7bdb47793c4390b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h384d2dc6a832842b58850347f662e266aafedebffd8e441d73cd69d6e087249b88baf670f37493d6cb1364383650382d9c235aea9863021dda4780a19e6a956a556e576fbac901a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ba067196cb392575639cca4bba579603a187c81a12d60f6fce904a69f7bb1e060f1b928a481d4865a794c2f71e714ff81c95c7855097238195f802e321f81b90a6f28097cc5750b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2531a77af453ef22eae18b2a069a834a394f47a545d972307cae9cb2dcc459a572088231c966525de68c73182d4f718155c130f28405a6a32f8be2efecf92b2c227499ecee53fd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc724fde6e59d423b98b7df5cfc199f42422c6dff540c731b40fbb7575689d8f966b17c357c9c72e3da41cd2f24fbf7ef86f2e9bb4f998aa8db70704e573a41be49ecbabc3f45fa33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc541dc0d4c96dba75e8e325c8aecafe027e27f91bdf26cdf082648126b55b15e524f95048141d225c05795799b348518a0c656ffe964d0f6d692ee587ca46a75425c4fda855ac4b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2e3bb7607a15d13ba2e0448254b4a51248768ddc05b5c794db976944bfafc54491692c2245316c5032758faaadc7979993eaa38b49a7b8cff7b8eaa1a38b8dcda36219580b299b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf8e1ade15040bf556db9315dcb3243e94d2ddc9636829819cd8b2a29d8cbc43ad76956204a25b02dccaa3dd9ec18963278ed2b99978391681954c69d6715b028f0c8f3efece5f4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3abc5191824e66d6f95459e658b97aeaf6285614c1b739aad3b54bf594297675416061894838f07b23f1e3cb7cc54b12d2adf4f34b56833d744e2df4d03b9eb1974ca8a0aac4a7df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h337faf5570d6094209836fa3269c432e04ff735fca0ddff4345136e049151bda06b28321be99148e6b826a34e4d601a62bc91afde8e692312e2049ec6cfec4724e3fd0d0c50b5259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa5ee0cf409d3cddd26afefc12a580395c2be7e0dc70d344445283b9446136d412541aec62407fc9f6372a1b578d186b9af20fe1f9570c9550fae0cbb5d96da00eaf7263e250d8f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83505d25ab989878feca9c9fedc2b7e291d6fb6af8fb1fdeb451e5e8c35cafac5f750d3217adf1c44c7b5afe242f2b0dd10615fc757d43d1d7fb1fb370b03e5a936163c7bd94f0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc83e4c9b26a9b743c44f3b0aa90f694e11cf9de32ee5e7cdef168f33efa2d165893f05381309eb0a0e506371d7bf74536137d3961e9718a05944b22ab3ac79728ec54a0bedee5d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccb8749054dd5a2a97feb4cc88693a89d3916f1e15d381737638bfe5709bddf9ca242976534326b903b0bc6636605caefbbf5889b658e2ef420b9fd809bfaf1cde3b0f2ba87a847d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64c6f7953dbeba352b7b48b226743877a49e6763c1448036447dd9c9d733777e8d88f68c268ddc4120e127c993c41095e313cd106f0752bef76824c15d9a4f87b1c435ef68c54b77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c59f7bcd8df096b4ed336e49ba2de2b6ba8e92748b94c03c67aae28676960fbc406cce1e5c10314669d4586c367e9631cef5cf244ded09c9a9d1517dbff99d1985a3c10645f7b6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c6f593a104377356a690a405d4b4ba234e196932ba9c1207dee7a92616ee855c8e4224f2bf7149e7109602a6f71d3543596d601297c3bb084cb1c4bfe5e088399de8b161e767338;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61df4ac35b05a82c71f7806db3a137675f1aa8adedd24ae05b5663f2f99611b85311c289c0c09fcd6770de1ca86cdc32393d0f08a63c3ae384103fb82400d543d53929692bafffe3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc982348977a306a5adc1cba23daaa90b21e028713f7c3f4880474345bf1c2027f16bd1a138076e99b0622a2807548cf94c6c58d0194c118bfbbc34a779f384b23269920a656cb387;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbff5a87d3820da8989c25e281a959f6409717d2a5c0564552dadaa18b234207b0a0250af17f4ae02334c55aa0bdf95e8063560036512e9836b64f060d3b02f322617c2b53c7e989;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddba0dcbe9881d686925d05c31bbf023b2cd0c4d10254d1d128e4637f2cc17e32119d522438ed9ae289173c4dec3648fd3b77c430681b74067df5ce3d49b0bbb5674ad973a0ee4dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24af88fb8d6f86418e10a349a2574fc3b264978101af955af8e05174d1c38c5ea56067bbd5f18f5ca8b1aa1bf1032b59dbb767521521f4d3b90fbbd1883eff1ab2a61c8e658f5ae0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48cea7611f69acc3cb5c2d2667e4af752a944d7dce26d1159a74356cef3977ffe06d9a255cedce22c5b99a49cbf5f3a71502ad98c7b44e4949a20f8b6aef9f4b29f586ae6b3763aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9e8f079b6d2a0bd019f204d92397c9b0200bb81bd5164f79ac46760787f7ff38ef563fcfe4b46e702f85e60cb123787bd2a519cbfc66b0c3ee2cce754fe2ab1a56cbe66f4357b18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19c064ad87f332d57a416b742c91817e9180c89bb90d093e44d3a95433a29cd4d17a94b7485a76cba7cb6b669f2846d1ada5420474b4e82e16eed9e55bd5344f124e4c31a11b85c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1a387a2fa3feff18e930d2d0476853b13a86d955124dd110d8ddf7bb864f0d9d8bd4df9992a769cb79dda1e250ca5e6dbf0cf90c9af61b60c4edd8491794ef5509ee0594d75cfb4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f2f082e061d4480c1fe42c76baee987dc8de937d6226849f8a035d81aa9b66802b208440c2b74c60c209db339183b85ba321089b6056af55b0017587d59bb95f6eb576214537c9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89f04ac4cb3fa91439b068964f981204f3803448bba4b63a94f08bc39b9e7c9a6a9ee0938f2d1ef2b09e00c7f0c9afc3701a3a6fb421b0e0a52a44a814ca4341606d3e87c9540bdc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6117bd8956008387bdc73be2915d22d863a9f9caf68eb613ce5ad9ac966cbfc9a82c38ae6ec31b494de39e0c24dcbb28b710a68925e1dd7ca304fd064756631b5ceff1719d9a3cb4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9e9fa5170fac5dbdaff78f84a46c07c24f83358245c7c010a6a7545ae284a24ee0c7584560a32f8de47c4ce23a3ebdb5aa5eeeab770276739ee0d3a8503bcafa8e762c68af06fd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h420f9282c77605c02a23e85d21387fb42ed2963558f21b7c6e007d1e5b336657b67ed347240df23b564265b8e5aa13844d0ffe922a08db8d00eb840661269ffbc89a911aaeb9403e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa662b02f338a57c4ab074f9a8555b6dc3ee94e39c42d7d33e8ce4290a811ede060241a098e02f61afc8d4ced76c02648367e51d2069b129664447ca185d2b296bae6eff8115a87c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e5d2f9bfd509a0edbbbe3b150ce829bc259bb30a654f7b1548019a7a32fd490cea86345059851567c8247d95c2c33a6e51d8bf648fc991aa8789d31cb78f9a73877155bf410dacf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12ba6b2f6c58080c04720aa2bb9173e91cea026dd9b0c792f07714e4ddd106be4ded1dcf21d205a96e376ee8e0ce974bcbf615fae921835dc59336c86fef0d20c4fd4175d1f63115;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b5850ece67e1accb7765ecc0f4e6e63a5e4a4b973b783e61a17ffdd1d65b590abf46bee2ef43eb598d25d198a23dd39fec9c93ab0fef343d3f7780753fc79672fd27ee07e6ab833;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb349df537551f57b1aa30fc56a643507e33c67f47e5a7f92e7d332f083c5baf49723cd2286a0fdff742e87231eaf5b0e404e9e0b1bfcf0e0103689ff191118fa2b64a5dff855cd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91efe2d471b22dfb43a3fd957539caf852410b17ca9a4005789aa86e144116b4c732df78375dc66b684a142d536c99fd49518ab3ba75b00b28bf3bead15bc934f1a47b6078630365;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd83d0f378432655f4ba6ac5850b55e28892ada20d5f4311dca19b95ea95b9b4ec706d9493b5526b1592c0584769830bb9f1e493e98f27e7b21093b389447613d5cdb9c8cb54d819;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb82fa2fa2c8038b3b9d2139dd2ca3e807252cbfdd31d4cec2a534c254e9b966b0d1dc2dce37a85200d59f287301c9d0892569058c120964a69785edd9bb636ea520ad51081bed15e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0c4ded5f852e230c9be6ab49f38d150183174f967321fdd674149af1847f1f7614f49b1bae6634f3c02bc2968a3e92c228afddb18efb72ec4ed0d081e491e7040a7aa7883dfc9d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac292a5cb1e89a6339c95fa34dfbd67c7e26ab6d480e2882aadda6cbf18dc961394a80898d287c559307d3ab842a86cddc04caef93f19001005b049d3d93025f1551d69ffd941dfd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0ef75401e70a98bc83b854dc76c18fe04a8006c78bb23247008c5dfc322f439db4bb88dead0f9b9e0cdef2acbd8e779a6472510a677bf1c19559e2569986ce1a995fb51fadfea2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h427462e82e78ec837d0904cc42704150ff301719bfd9433a6691ede94530b72673af0c34a049e379030d3a438fe57c72ffdb0e571ce31f7bce6d7746b511cfc0fc5a374ba8dcb469;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d1a5aa02cf1300a6f9e8b7546217c7134ebb706e5b6ea25348c490a7c831f0c9271a2d93ffa4d67bf261886e71c4b8e3142eb434726e260a0a9dd51057fc185ba221eef9c556aec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h268692c0c7e3bab9db3d78c629e48a3eb92dc12b7b6769c019ec6c0a35fc58fa071bab59d54d0b3305b2ce1488271ca18c1cd05b97cc0a8919e2aeee15f27cb51724699bfc9324ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcacd9a72e3fb192ddb37d96f4d44119629a30aee88a13ca91a049d4e5213189c55abe35d66e68f6ddbc82847ed6c7eb8da0956bbeff803e29e0e5a02257c4ca2fb8d296702baae5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1619770599c2c9d08247f2922f6b1613d5a917da6de2b21d0eae2c15f993c7e27991e76bac808c5fe7a7f82b1ddd7a51e7eb010a154828a37e089702a41c3a212480083f6dfbb28d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd34b0ca8e36d0979efc17e6c7eb75a68319c2ee902d27790a736e3c2f627983ec754133b3219762f68d8ac6a4c2a3417527955257652bd666bc923335e2bb4a00dd808fcca8be73a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4c1b911b0d81e4d331b8f4c26177c85924597889fff5d2423d49a982bbbc95e13c7de6a0d608de8597110e989b1de5a495bd006d5afa493780ba655fc473845e5f5ec599afc660a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe2749f3a54a1641cf6cee4708f927b3dcdd3f62097b892fe6c0bb1eab49325013c39806bfdcd8b18d1fe129c59bb4744f088d6ae3e086e39e2108286ca84a86db0e55d53368517c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h693a1079b323c6128277ff8577bf932569b884befd72042f8b4a9c7aa5f1caa7dfe778d7813e58895771651580ab1c8f833e49252422cb21c739091640179a9ab2f6cc8264bf5eb7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h382e55bfaeb06a4c4b133c6082826b9cd5b92dfe9f2bf0dcceec17a524627c2f39d7d588b0c837a31e0f893d60de5582a7f3e45e098afc943b9fa7534ecd0b3869a91232f2ad381;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc059ad9856d0d6c8500f7fcb1e3bd830970b01d2734f375533723aed20de377cac8e46db9f7bfe08af1602d09bf475acd6a02d02391cbb7c20e3cbcc547f48bc84a91612d9332e03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab50129d382e78b8b162785bd45b073f8f944c68f82889fc7bf3311073ba8c19cafa063734a7e0ca3a62949ea6822a551b855f4e60c4adf9a9b590874faef93923ab78e8820566c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed63f5542d0fb2c04bcaf6b904f4857a1f15aaf6cb9122cd98f7cf59aae6dffb56ee0cc69f9cf7c3acf830ee91fab81c12d6214b5098ca5d6ee778a39fe78fddf5933893709dbd95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf90ce65d5f082365db562a33f7abb08622e02f9456117c42d94c48b81974979fecb43197c5379ec1f2c48058f7a64a1e4dcaefe650961f622595e6a4f1ac94fd0e270f7fd4006057;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa83e289e464758e1c340bcb01a2e58fb571297495b0599d06741a30546d70335bc21a715fe9d9500b2e3d212abee1f675997522682edc003bc61b70d12f730a3a44c7cc697b3a6d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a921de974c192a4e0641ab08e6d46996a11e4c3191b20f58ff9742b01bf1a9d0793cdb7e2756fd6cbe84d3ff354e89dde63848827d0c9dee7c190373f57ecc69354b0fa3adc5446;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be788033357ba1a404255abaa2b0e824828929087165b4d91af9859197244c299534bf76b86990d6075fe7e9751c3c10a4fb2f4ddca3130f8b8a0c5fed15ea9e1857193c5c6c7f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc783213a48db3b02a3dd739da1ca27242bb2c17c2a18783feeae6e1cd94b15ad055579b85b608e0cb305d8362e5a637619fe5b6021c3b2ecfbeb8a882828ff68889240785e28397;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc88cd9acc021b22cc4f2a6a4fa208af3301dcf8e602da2130f8771e7ca3a1c16b345c75795477f527c4bf57f19793d7c1c5ef1cc2ca5ae3ea1bcc33bb2cd2e0d92f5597acf5f4fa3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb5259d8c4136ee6b6642398eb8fdb990917543e0ffe535fee00cbb63b578a03c35fc115e73112a1e435d8ba36817b4a317a213cc64c0642ad7caf8943fdc7548f80da856454e016;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h317f19eea784819317be509aaa7e03503820f67dc6e8310b11c129320611d87cfb56d72b88d765358e8042afb7816c79834007a8fa2614e926f6a1e6ef4df36fd61d4cd479e22273;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d3fa611762c8f27909e240ee9b7d1e55ac77cd01346d79e0c6b84f7adfd7e621bebdf519c246aebc3a2be18f97ed368e23ad470752592e66774d65165252b92d843e4c04bc980a9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8063a044c2660ed9821c62d4dba4b971f54ff3ab4a9eed6f6601443493e2e425d83313870d5bb17e72e8db986419da7c97e093caeac210eb14ffb2b0aa7c2eeac878244041ff80a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h616db379bbbc58ed3ff51cbf0aea8d1f1a5937e5159787a64df15fd1ffcbc3e9d4ba4cf2bbcf80e12ff0c9151a5e47905d5767997eee457cc3006d4f1fce834e4569db20a9acf934;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b651709dc1d7d52ebac913c12ab5e95609c815fe9dbc740e760557efeb99c0bd63bd922a2047943f4a351f7f14fd3affdfad61a3c490dfdddd128b27805f28adbac5d5d15c7a725;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h722e2233c535fecb419abeab403bbdc69ce1505d7d24f14ff89bbb4daf607f81e322076b3b5d61b5443a60222387c15d7e0c04b9e5f11914a199c2a6c8fe4633b029542e7ffcbf31;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcf219485d2d61d7bc5e4720f0351cbbaf7f18edb60bdb012bba1d5e7ee1e3d75f022cdb70fc60af51e0c36e1b4b5e6514d07e44f5bd3f2d2b5bc89655236aa3b35c755b92191c4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd24af7057363773a192e1542465cde25fb6656fefa6039523833219d12f6fdf091d49875b94922063e914483a2444f0a2001874a5e11eb2ac0b99d136055a8c6c9c0dbc041a3406;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd39b234cde1f41c742b3adcec8abb66db442a154923bf7a5f2bf597a6c97b212f4b3dbe1976f2ed8119a4e3af1a1ffe1cd4523a9abea77b61950a96db8c9a71d84497293d9c7b969;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedcddcb966944c4cb573e190120ce004ecf097934603960921cbd5215ece47b335248a0982501976d0b65940cb3bdd9eb6d5c6f1623d76e9ef447628aa2d0416580b8b458f754f37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d18f0add0d2e67ee974f2b6f8c45bde35105e27f4b86e5845d60359ae3301d3795447732aca06288b0ef10faf419593bfe2c5306a079e5646b36daee82e23cb5d1a2896ff0e8cc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22e203ff6416ebf9b3358b9be34356025e2524f180e2b554d5807bf1d81cc2090746697a2795a0efb4a133047a4ea2b2109e1030b9cc6a5b2cac882df3f3f3e52cd0abba88b86cab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e5dca156336d20f2487828cddc3c9d572126dcb5dad1c614b27705d5941813a54f6c672ec049b5be3dd20b31c2b834e2859ef0d290f90198f07ad6e2b820a16931aa2eb75930322;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h185df44f09c94f6b0a029667dfd7c666b0e3f547f33eb2db36b0e7b465ef66ba18add87e29b88f696b89f3b0cedc0fa4704a082d592ab6daca2406236a6f4c84323c52ba721b72b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5602c6733212043c7cf4deecc91b072c6e84c39f4bed657009e330e5961c499d7b49b3c8bfeccbd44e2df54df87ffa30d458f02ff09efee17884ee820f41f0abf5756bfa3469cd5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70265a2caa7c950ec54575dbfc5e7413f7b8b3cde12dcfb3d8576fbf5cafdd2f7dfbcffd8c65ef34c92481b73cc573c8f61c16893a280cb4744d6cb70296c4e3ea0cc45b76c46603;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf52c99f90d9438aac8dc2ffd0af300d86d5b6e4ab35b29a7840375341c334e18e5833833a2027c61dc23e501d11a120165d77f07267130307dafdcc2d926237c22ee14ef2e1f62b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33ead8d3bdd16292e4734d1f698c8d3f186550aa73c1c9d0b869ee031751b11c8042c8bde12ac2a681e843dc95bae8ce99a51a72c21e357e7783e8a1f6ffc863ccf9beaac2755230;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56c3fa00c54d068830f39269dfc6b5881329c93809a4cfc744e2755f19a3eb7fbd1ace054634e451307c94b1fb7bacf68f0ed0c0171ec43283495d17defd84c96e8c58444a888414;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha66c873d45dfa1a34e966c9d4312310472545b9e9efbaf9b97a8b5a99fbdeed79c4adf584dac8a84e90dbe696f693ab1f4218f9a5a60ef67be099cb10a5c3fa7eb650fe0b4a21136;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53086045fb957fe730a39bbc151f429cbe8154fe5ea2415ba271c2b17665ff6b6c5f15083815a267ac84c25a3bed76158fcfe00478f1ec95baa58b5ead5b6b1ce51a0f5ed0d0e4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h562ee8ca4db0cb1cdb17c17a60cbb629d53291d90c6285360b864f1374e63b2683923a6fe08fddec9a6737c2d4e231b3fc9aa8868a932c65e7d8f8ab5f1067b7366d3400b37aced7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee851dc74fd29f7e783c74584e78a9ae8a49775688195ed442756becccfa7647212dcc695fa358adf9e061bc4e7865af43bec7a234216cda9332290969baa687540f2ef503fe7961;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe83fed9ed19e7f8c3ea65cfb368e89231c54011927bf3f7c429e2991cbb290a02eb8598f73a85d60c0b9ae17a7923805ac85f3edd29261ce9c5efc86005999b1c6f83710cc41f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbbf82dda0f4c4504a1bb5230104e36eed34d22249d0151c77be44b6949591243ff041e1027165d443b0e7fd1a2c9430300abd16890d40159a980a80f94fd2cf9c0e190fcec3449e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0e8d4a068f490c7f32f9009a34729c233813dd16fbafef685c2c91387c6d501c8e8d54f8aa94fcbbbb9d66d5b7ed926ed32c013f1f4066615c036a5a60e0f221e94949e4ac0d9a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha95918006c0f8909d985b1b7d08eaff517b00613858306d0ef3861be090f1fba0c7c18255aaa932ab920e7b935d8dcf2793f53850074174c962b5ed45353014a6338ba26274e0711;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ef753e891faec1b040072be58751383fc72340fe8cee6fcae9c1656ed2852c94182c354fe8827972ab5d8d5012adfce464dff6ccd61de975e0911f8acb641b4e05e50eb17b3001;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf01242576dff3f59c4f7739dc4eaa44820b7dd85e6d9855e95d2608f21739069a85e1f5348352ed78a921eaadbc0c53c71232d8967e33ed10351859c4cdd21d2e7034ee83639cd34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57d181771121261b47a087a0e35cd762ec294b0180c3a38aa1f3b1fd4e94a4e6b7ae4d22876a3d369d476e303cc450ef5bcb2014d59cdbd8b6d65337f49d3872063c622849263b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5d2d042b36e66be2389297a8d08aa556d8a30cfde75bd1b3a6222b689e1bde42513d68dd6d94f81de29826ac9d372051ebdfa8ef7cee0c7836808be9ccc3e187752d4277b92b594;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa45de72ca344c919d69da8be67a1ed3c9f714b5019a36b3c1d5ce9af9beb0cc080006e1b7892b86eb50a0a4c19de20b42e07c68d9e40a31ed2ca509e562a1620e3b892fee17f0b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13363a9f2086bb18ac05634b027c6bbc8726e928ec18553b813f72d9818d51104fd9b1e7910ecb02eeec6d209b6cdbd0341d73f9186e3582f066c1b7684fbc4937978ec8af83c941;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc49ed4ed6f814dab2b5a8a60372a61959799b6980f9c9615f0351da6dbd7bd551b5fabd08f5aeb3173e9051ae89dd1eeb63b300a6124c7e77347f49457e8a725eac86d8d09817b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h176d6e04df6cb985d68d07f87ca8b9d999551921cec00c6e1670547e917ac17fdb994b8790dea55deee4609ea801f7d9029ce70db9f6aea5d8ea0b6b584802ceb7119e0894718942;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ca02685cccf8193c8a680fab8f8a3aa4c85dee043da1e7d583905e475b48c27d5e31bb3d6d049bd91ad597e6ad201513fd035843b5f6cede50d09eecece0be21c854fc8173c43c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43a4d94cf3605fa293c043b35f353e2ffa4dddd306ac8590ad84ee8b8a3992c4e32312cbdf55bceae32bc8efb0264c460b43981a8ccfc3bb5d94bfbb9ea74ed4008cc7d01f72c7c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h961e4baea5c1bb1b92a09fdeab15ef36a646a0de24d5a3d8d0e6e1cc7fe7a83460538954d8e366ab7c1c35bfa96d43da1e66895c64dbf06646d118b35b7317368d3f0870b9f2405e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab3e7cb8c4c569bbdb8dd7e82df13f1e2fda6f056ee04966f194c8ca8143bfd804747d192aa62645915793f895015cd2b804040daea262bbbb05d7d96d3ca37c1eefbc6be6441e17;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf38bef5b1a4c05468b3ddfdf2e8b158a2a76b3df9dcada264f2830c18ea325b248f469982f495d3efc1b169df5700bb8f5b7e4d2d902e814f82af2d7c8a424be1a68be0f23a4a5fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23425425ceee532035b611d26c91c78f10b3731386c83d08d3c6dc3586c2c22eee05fa2bd1e68c1cd54713b7df07e73651e5660e7bd3c7a3fa3ed6a6766fabd8acf636aaecd9dc42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf08496e35908a0f6dc798ac31752ffcd0ea03af3bff0ed205e471978ce0b390c3237aa99918ad5003833350847b74999343e49e874db9053bfcad959799334ba10ca3d387c67df62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c5baabd59db619f854ed15a21f6814ca0b746a3683516adee5a48250735099cdbb8485228933a0857ec87544fe111934aa9d232ff77bd7ab135a42943c96becaacc9f9f8169d87f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16b22580a34410f51ab02173814cfd7b42947ad36102ef2acb2be4f25e4dff01249a1a5053bbdeb8c59148260a06f5deb5d509a1cf8c7f3beff53ba0b61394934a663950e23ef3ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h203122311235e1dcf6f9c4a9cce1bc25fc506f7aefd6cde4226fada6116a80d59df2efc7d1d5bdc56f7a55d276b118d3a4b91fd9f0c00e29bb2ab188d7ffee9ab39434ab9d5c52ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefaaa2641bffbb3a5a8722b05a4852891f5b059d50db839c73076197c02550d5355447b2c20eeb772803ebe71e5a304024df2c886bc86f65a0460b82647d3a3a2d063ffdb0f2b96e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bbe57c9ada96563b2391c302dc600a06d9b0150fc7954eae87d8067b65f6cc7f4aef51f4fb70adf62dab9a55c2636dd197998da3a2e87109d753b22f943a71eea02de4282ad6dcd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d64d75b5426b9361f207115c88410de64239b2659a8bfb613fe778b7d64f594e87ff5eb9450a0f20c10876e23370b13ee6052e904f7ea00171fca51b4cfbff9b76914f406b59d89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h848f0ef7d7ce78ca86c915a28c40dac9487f5860d409c8ed9a2776169ae9f5b77f276447cbf6616c160244807568b5f65fa9cb091542fc0c9a66b042df7d7abcb2f48ed0728dc32;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d356df1baf8c782dd76f558e8e00b9e043d945e3ce9988067530edefac193800f978dcb766f04a3eee5ab77e91f233ff7116217f997d673151a9eef177895ffc1af6d54db67dc3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h361a9f54fb1584ee05dd21082a6c1bf73c122af760efca394ca2a72356c32ff97acc82c8df2f9f2915ae000145eda09c324d4e0d519f4da59e276f4a1db0d39f43ff81449281df2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ded45324971c03e451ecb87bfc393029e0e910604d28fb461d16ceb815757bce7cd80e7075bad3dc7f0c43a24153412ba0dc10a4b0e13ed2609f811bafd8173e3f30ee9350dd02c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he922ee483762d9566b14d3c0439065a7b7636a65261d0e524a798a2be9652a4b8cae89ccfdeb15aea265ee12dcaf68dfd17711357271314c2b89a19af662dfa206835b269c19d8ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27d7961e7e8b0b5ac0e078b3017a6135a88dad8ad4c46ef67deacddc4f203966bfa3b4c45f4941dab69d85c4f4a7a64312730c482637034435753f1583a8db300bebe0904d996793;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf33ee26d851f4dd60549c14dd47e37cb5dfdb7396e340cb7d50e8535687db8ab68e1972771b245542f84a3b43187a9723acef0e6d83f00f2bd165c0e7526d06aec8f71fe19447e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a0996aab213ecca436efa84a8329ad638942d02224472feccda04ec1e2bff6d2eebfb67a8a5cb73f6b0b08e9258bb0bc4c774dac9c09e401bae12a8bbf8592704947ce4f41a2083;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3579ba7b553712010aa407c9b702cc0145b5f7d7239b530ecc32b7f06715b6c01bd7a4a1a1833bd65a176fba6f140c0fb732270842912d4274ab5f1ebc1de9d27ad378671367c86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5327a45b4ccbc99e8217f9d62d60674c96cb1ce7e3c313cb2f8b0ef3debbe0245602430c9f7b025155e294d7f1f68d41d247f0352b351a39ec2e567343c0f4c7de10926bf10e76b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1201964ccd27193b69ef74065c085d8ab5dda2bf1b1a51873779558869545d16cc5c47e81a40481040a42ce97f5cfe5e0bc062fb78d24186e25c934ac25734bd55423e67c96a486d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4ef694319f10fca2a3ff7d5157e5382f5771bede81a2d972a0262c2379f12ef3b2b581ef293cb83c7de8e22c61e38460936ed5e7f2ffe7fc5b2ca420b2c774e6066ce3e8a0a6e11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha307f91a116d4e249adaaa2b0a6377ec3eefe15f8e9345ba5bd4438b8a8de4f740af16b0b34b6ffbdf46994defd7ad2f8a9dcbdef87993729197aa05300b6841b0e032a053d0e408;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3c5adb2bd3fab0a02152b542266b45c46e599fc997cb42e448a54c03f0bef4bf324e0121bc4c328f5043e03aff40f97b60d7a5ff5cb6fdc8de8e115f7fa08a13441479e79b4ea9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12733c42e61775438c98a4968b7ac55d661c3f48ecfe59b7f8ed9ca444df3c32627f1ec46d76488dbfb642a15bf210f64c2435901e4c547e2bdc07f2e92dec03f7618f7f7a22e680;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda98edf99be70f83d3c6585f8ec4e2b00777b39fd0fa3df4d8b5d3914613764c4b9face9fbf21b91359287815042ed4d7cde1ed64d107279b10739990fd095e1adf049aa06d10295;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69c9a4672e805ece7bb1a09cf5f4a3a6a81e9d3fcdab78191c19b5704a99339457ec460c626924b0d887d70e868754f9afb5737c7a9ba0d400c4bc34644439bfcaa2ae3ac0342567;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffa3a4082de698466e77594e61901d0adb0e510cd8a9364001523c141b19585d7921e8ee87e9f650e9834a821c0c6be4ff8de2d9c24840634a0ae4038f8ce655c44a3f6c60449964;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f05a4e991c59a6bb07b47517e71737dd32eb0e8e7904a1ef13cec5755a66edfc7f415729752677bd9deb31fb05b60fe5a95eba742b06ccb3dcb6dd53748e1c80a484517e9d33dc0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fee50bf99eb2390d25a27169c3cdbc53fc0a5f1edb4b8a3dc75733124b288ed0de708089ba27998de4639ef33e4e424d51485b21d935f54a5df35db4c0ba0a3c19e5d57860034ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h520b9eb6e2d488b43af7563eba682f1730ab1ddfdd0ba279403e583feff3623dff7d311cdc64106ca5b6dbb730efc681dff0ee95aee4f9b33519fa9fc46e9e5d58aaefd865ab4a65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha82e2cbd438d9579f0d3377c9e54e5769fb9b5b583602422eca31fc7e02f4c3ebb5ffbd8ed38b1cbebd5ad8cd460792d5de12a406ba6b99e1d7c9b5f2724bf34f3959d703064420a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca32d039f454b2b757962180701216a18e31a13d398338c96d3b9882b7400d47e47891fe986d189b38b9e45fb8e7aff58cfddcf75d7a58b58de86b8597f16436f53cc458f4fba90c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecd04671ee493a98debe4823d3580ab7850246054b0b33d52e33f32b5ecd35be6d2e253afd18c995cfdb7477d6923b2bb6ec04c92aaa23d13f83224dda532363a8e3ed2634874eca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb99502848e423e4d7ed1f31ef12ba9fc9242990f4cce239f0b7923412cb25a25aedf40b7883c045be191bf489ee7d3c652fccceef1f05011286eb97aa32056645db01dfbf209f30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3e908cde332a0a29ae0f0f9cf4056f0270056dae68f11f920d74b24763c223feaabcbcf852bd13595763026323ec3f97cc9a0e393e38cc686ba7242510eea2c9e91ec1375b8110;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74d2af05f3ac0a8486f2f3549067fa634de6ae12db8935ae204f21262d12edc8b39ee1b07d0d291366e38f4a8b2b33cad02fccdfd3348cfaff7bd866883706aeaf0bbcae652e0015;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h362a096c839134a381f97ad6416f91546cb876e8114d954a6c518b4480bbc1a338ce21555fb35c29b008525bf1381fa897648e3b955d9574d28ea7f9493c04c9cb276d7bd3f57909;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6b5ddd896c551afa8f2693a70c93e97ed651159677abb18078146169689db7f49c0d257383e00e53b9e6ca460410c8d486616530a44815283aac1879c8212c4f248479dcf873c94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92a6d2adac7192614a57fc3f8222fd5763c7712fd6f8392b9cc7eebc56d1445ab57e9dfe5b07a5a2a6189c2ab11a308c33d2421abb1e9c190dd9e242e388b77107faffa8764b7f5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha36d27578f2788a7dc49f766d5d5d4d7571b4dbd87d43dd1861b04e6f1bf67bcd26e69c622696299aafdb010779a8946dc8ced9b81706f5544e624208213ad3aaa410fa9ecb74889;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha366b5acceffcb0c7d68dfbe1b75d2852e4bbc4f1007c27799a1ad5f7dc3563bd56a63aacf7d8d444de34989bc1e9fef6f8f66778eb029b5767d977687e9c7e1d1a5a96de51595e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2368ffc698040acaeb08a8f9a7627a4c264ce33f04c6e360dbf97b470fde7fa0500f658ea8f2226472feed7942e78cef3201d62b6cd2bff1f1816b94f29fd97d95303c404a2a7369;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0eceef522f767a9d1d8ace619892636e580025ae6950457f97ff5b4e30fd9f8d31535fe0b679511c8b16371ee0cfff503b5f04eec4e0d73f8d551d2eda30ba2a5860d2c28df9a49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc0dfbec845df9ef3ff66ba7a61a3d748344e6c435db7820571edc158205097483d6da918b8e4e9883cd5c341ad586ea1d901daada4fa5b128e93b764d6a2845e1679103ca192d7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cd9bf5e6afd87b37774f860ed5dcf28c3844b520b464f79599ab9d012fdc16d058ee821e17e8b8119c1c6b4e332729db8ecb262235fd3b2bc543fb33898e5e17a2ebd2bb66dc5ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58ed0a6a3095cac8e8c54018620e10c62b4920d6432ac8c3b70b4c2d7bec1fca83e5dfcfe4220dee55133ac15c9a0dc68db255a48b7230f3b1076dec2e8113f3b87ef5aec8a56627;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bfd55dc7573f0f8897908f32b8c52ad6f6f68374322e5dc1dc2198910dc8e5139150945c43deafc1ee4bb7f6b1e9b1d74f2775bfc5c4e34172be6895d31e995bac7aa14c18af5b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29c51278d5b847a1fab25f0dc925b71c59db70bd336f5149bf08e3ceb21d8e24a50ac48cc48979d26211f62aa8fabeffc7e95fc0cda15b2c3a45f2a64457af1c655e87e3df13f97d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32e57c5f0b8abde79ac09fe6723279df0d83302cdac041b7dd0b498ff3780ac478ccee2a3df49ad35af11ef2b209359a133567f6fd7e0a253281034fdd5c8edd585d3530c69ef570;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d6be658a6fd31e70b2a50d5843bd3ce138db6d06b6c01f0c722a9ed2e45cb1cfd7985405163196c35d2aed75b29e99a6a3b5aa1645c930c0cb879692008317769cdd3213d1e0eb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h778dc129d6a3d86cf31065accd5e0a41ff86a2afffd9fa266d948ba923bc44334352f5922a0479254921260af1cc8ed30d3b648a7dd2a973237057a37bc68a2e556b88fec17caf51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e5793789246051d9c0543afb05af15ab536717324f10a6ff50c83271e3c852d17c8687f0fe44879c4288afe7f8cfd1c5b74abd370f441b5883bcc0ccefb162c21f9578428eed277;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ac3af16f00de62e7a2f09d5d3688c3dd2ff824b5a610bdeeb6b9fd30b8cbd5d01e3cd7d078faa2f50aec6b93128010a83b2ef054807598d765667da2151562d4e4e1572af115fb0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34742551f7e0fc50fa68171f8b003c29fc7d8a6074b13ae77194ac86c51397e8e8695240f51ed10bb79c3a8701023ddc752204c71050643db2bb8113e32cd5ef9c24bc7549b3234;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h505168271ed1898eeeef81257959e57e8b12721d99a086c2fa159b691a0815be7f06c7c362209ba1dff485df99dfdbc720efaad08241c827cedf96e27e4c3ba26a3c84d1290bf112;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e91c0a0cb9572b2311ec184dfd7ce0b2123a3822556b46df710e3afeea6640d2901ded09fad30fa698339bc3e9c4201680893061fc47ef48882d8b371012a471ea4f41dd9df03e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3becd5da5e931af5ae599fb82906c08973f04a1eced29d00b594933779c5253ff82d38fd16f48a49ca81c41531dcfe9748cdc9d8f05f3afd573640e2204899ab4671c49ffac9b731;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f71c1110ffb88a4195162202fb535fc0b2a60d4653820dd506c58d1de00c68ff9d589e005bd97c5cee84a992e9d35ccc4b0dcc1eaeaccdfbeb3607f181af93841bed35c99402e1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef3f61c2430b94758b05320292a94c12b52a960bf8ac883f9fc065b705bc856cedfa1803acad2b37bb0c452c19c459fb7fd887b51b347a29426ccaee7338ae31cb95bdd7a43b76ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0126c179cc11675cce7c4d431b4dca57670899979616291d59ef716f6cb562ab4d8aa78e036f7d85522f10f9ec43c4ec500d78b45b9cd6ce26cb9ef7fbfe3318ed5abf40163e7f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aa20f03666963e94fa102f69a64dea1ab797f152635e94da52e493447e1317e087ab08929dbf00878401dbd16f82663520c1cd67b63e1416cdc306a7477e29af9919516054969b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76e615a37eece6e47d039c373568c169481299982068bc97de8867090549530fdf79bd7b993e03fa0e268d2990e2551ee4ae843294d28bf59fd638d1f3b96d44d1d2b496a559393f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfaa56866ccbfc600651d4154610cf64c7b03a750c5d1f6e024d3231039e565bf8dbc58ea101113c12bb98661a84aca78c561275b812919f87e99dbae0f28c37a36d60d8531f9195;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ef201af118c80af8630df0247b59fbc59224e8a01cfb47908156650756031f287607cd2f684db13b5a7dd7219567ce9120d32e3173ca1d9ec0abf839b9c6a91e6b30ad796a159a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53afcec817722467b8786b09b347209df65c3b34180512c3b2e37b4e222ee4cd8f7a38d004c2dbd81c7a3249c1aee19a7ed54f91715d21b0fa56f25f735c565565e4768840593fe8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he29632a6c3a312608d1c1c052af6ae24fbdca631987fe99ae27fc017383ec423cd16796d00c5ea01f908319d15d01e3039df4b90d1d5900634db54cacf2c8b9de4392c873d87be14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcc79a01ebb8ee73573f0a5bacb6bebfe8e01ce5e1a3ea415d385673b94e1727e95ed0bf4b9a36997b9748b4a4b139efed37eefa94b0a8e2d9b343541b225cc56adcf29b1989d7d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d1a9cd822f6cedefb7160b9cadf9536f6773a5250457803d364948ab245b503bff9ca7039fc92cdb4fbd95d78cd68f547fd06bd2cb787588662ef5c3561035369d544dab5f1c1a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bd8888818a53680487f452fe841b761a7025a738a1d856d79165a7bf38fe5e87fd915c36ca8f8012ea0a2f885f76110a96026e68aa95dd9cf1addc9dcc9920329a7fdeb0be196a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h326a6cf50c21491975f92dc6581fc4c55a4cdf52462482d643f089701a83d7617d550fd32e77fb0bc708a9cf9da693ec8eb8e0da3abac4535f31370226f4caadf1b46ce7bec4e551;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9170dd227d3f4766251e4464814411fe32af2bf2cb4c7d91834331b69c8d8fe11a3d09794597d6f72d2244cc82cf9c442d71cf988b2fd9fd7b46084146b758a9e76dda04bfc43018;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h919d0f302559da1624e7d8b0d8368ab49c2a4a4c627eb5e3567155771aaf5971739d571a26e75e2aaf4a84329be748b5795f03fbd36e1368f73609e2822c5c4b55ef0eadd33a0106;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dd5ceb769462af29acd63d4c70c7b1e0d7452facd64a5bba6673ff888a839316a05b79c4c947beb743f42111a0d3eee93bd19ea2de42aa75e161ae8d6765caccfb5c7195a090a5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc633f138bd1536165a81735a008ffb8660408a2ac861b68ed075348ac9df403e1083488af64d4e3fcd16d1eaf0144545415e5660f41f022fbbcdedef34b7ba0948c550a64c0918f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha736ff77955b19495afff01b3eefe6314a4d19d1e63519ae2a59ee36efbd2f4eb782976393df9a55658b61c53e5c931f46346266aeab0f3d3e5553c23f347f3c812480fcfc8d5461;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce65f1d9e6ea4578b458f7f777752e1e690ab47d9909a35ec785e86d0c211f58c7803f68d828f7437b4db5b834a1dda35a4428ea46e3b84eaa45a2de34c1cafd625c028e0813a4d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9f7347d063b7600d4b330a9af08db3c31db229f2f4c824750c2895b2bb584012ca60b312cfddc67fc500ad14e1765b1dabfecaf140d0528eb9b494de20e4a39bfaa16b0955135f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9f044acd8fd3dfb1f30793e4c18e692adbc9d00945419c4d4eaefdafd0eef8f5e105ec07dc45562e627a7d98ac9ead03f1b4529c8f5350b429010a35df46496193968a918a51aa1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2e936dd70ab85e5e9b1cb4c846f27c0b98192ecc8b6a6c6b2ea4a2d705c63f3944560c0f18518e866e557bbb05fb5221bd82ac4f1dca0c36bf6574bcad6dbeb451b7ce0def0012e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44bf970163cfc50506da5bdb3df8446b8b77c93efc1d85266cc26fea131142ea5ec3bf6c076bd092d5b89de16f1cbee4af00089c20ac316da78b830ebe068b7c2394bc52bd72716b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9545047847bca24f8aa4b16135f7f864b8d5ce715a22d04b3711d32a3eb1f7954afcb45f5b670d6a98865e80edb03a3d94807f70de180436a7cd6d08e58af07427994d9a9a25237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9126bab87f5fc5580c3802287c7e2ff8df3d25a4bec6b7c6d4f7423fa92fd564284c0bef88ed4159ccf81a7f45a2f1a81c77248e34617d46f7a9a17372f7c83433af3fc2ce41848a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b5a13fb778e1c267edf4692f73997e1dd2187dd8150b662529580bac8ed512962a2e436fca9fc26ada7bc9711f5e84df25c1eed47221ac8dd79f658d5457de5a99c4d8080648189;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf269b81bedc4349b2a6cbae38dc348cce9b01a84a9fa115cecdbf135e7b4f23cef505c24b014eff5271b95bdc45f10d7c0625113a3469120eb25c751d1873cd75238fae2be944e28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97706fd68c588cb30fe03ff57283373a2f772876e5c594b350561af66bb6575405624596818c12c269a0f797b40ac1f7b48fa7d3dc9c5cecec323ddef4102a678c33c984f18679ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66cd06155dec5aa78f15d9b6482c01bc57e4499da9fb06e67382bada856b287c092908b75b842d0c5dd31c622ec0c9f7623bfca8ea7bdab0ff3d769a678ccd2364860ee97501b39f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73ab31ce80927b86583043c3e5f722ab32c197b2f53f9ca87d07bd9f1f59717f068247605e2e58df41d8c42906d7724995b3482a8d08131d46272d068727462095a905861ca3da05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h671f9151d05bf5743e8e8c34be327d3c1d1d3922b1db6f19a29e508cdf15cee68643ae2432bebbe6799c6b51d774d1eec7ed687adc82f9c9174f5be30e0064788d408b4797f590b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53e12f2004281e7ef6bb81207169d8b878ead6b5f70ff0014ba36575bf32be106fc7d5499a16b725d93f0d46242907fe0f54cba927d94fcd70f2ae8cb806c374af2b76979a7da1f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3f94faba2fb5a9211a3bfa78ae57c0b894a209821da027207196d5f16fb9d391f46e84c26872d9de9d6c194f49794a3cac0b353dad0c38e554f289c63ca2c5bb72433c8ed525a6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19cba58d5648e6658ee3b01354180798a61e73b7e4a1d79b241a8e54b6d140ffce2fd3429ccafa16f31404a2aabd185411adfab87b7ca85431c3c57bf05c5a3226460dce23eaf42e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc5e2d0e89307a7585ecc0b95cd937af3163abedcda1d561d637da1cb9c0ed023b55b2f7b08d2eec266bf8deccd7fe5e9f9fb18f5af759e25c54e145b95c7ee99f257491b18cc67a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8789b3a8432dd535adffa5364da132aa108894b8908639480f67adb2f14e139b2dee64836912e037047100fdb031f6f06186e36a4d83f3f4cbdf60214285770d27510f5eb2a83517;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d57adc5cc14e9beefc33fb3c2cc310dc63417b2b00d55e2b42fd2248cd834b5f510d93959ae4a82beb22e6d489f6f80afcc8b016b342c7da064949a6dc7e948a1bebb6f2a85b5b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h749ba1038d7aa83ae199ecd53aea8ba391f2e45837f05d1fc12da97638b4370a00712c1ec09ed20b3b9a63ff1d6af07c6de07783fa4745885f2bb9f9b3ecc9c68d6a2597c2f80f22;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he54811e23075f22c16ac225f1e560199a947bcfaff8ce0bd1adaf319b26c3da642523ed2ebd4a9eb9dbe0db1175ae72b0e00339d06ce682e24a7a240fb92218cb04462d05f06cddd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb444d30dd6ad49073544c16f1e524df72951ceeb9ec45c2aa85fc75dd28479701ce9ddcf042bebebd3a269f57f8dabab4639839ed39e1eb47e5ea77dbddd1acdd9bd39b4cde62c74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e50e97c06d14836ead1b51feb920824e5f4a317cf62dc03814976cb6273b5e9ff1b03f203ceee644f92f2e9d6f95741875ecf5d7b7d1ab329d7e2ab8a53a057ebfe70d81d4be219;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57cdd71cdac285a466305bf70ad9bb4dab1fc192e737ef65a3fff4a90e0b386ac22fb2721dda9dde4a97e63b9ea08cdee358d60db514bba3438370ba2bb6b72332002f826dd38594;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90e30aa9d806ea3f603bd6a5c1bdd06ee318416861d9cd339b83f40a091b9305906da8a43f6e690bc18d6cb871c3c2a717ed2d73ff1e5df022317d9597993c034b84ff00c38f566e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fb505cf62bdbaf67ffd5d97680a1432d5bc16e68668a9a3d8f8036f5d6d13b971a001096a7547f3cd1dbfe8b74cb8d8cc0ac21815e62474acdebcdc43a205f23f43e9c007efff56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce5ec8b54220403940f57b772d99177b9e4e0a1d3d53ef87e94b065476999dcb7fbfac2cb7693932ffd4b462cb6cc005dec5bb8c3bab54267362909ec6d7c23e5d483268666175bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd09f45bd74857b4c59cffa0bbffff9d6e4188a264eb4bda9e456949a0764f0ada0019ee9cd793894cf1398cae09caae4afde46a80e474aa99e9deeaef24d98376e23942c094ed9f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2e306fcbdf1da03e9485d198d62699e66ed1871995232828f5bf29878a11cd3418e2752e5416d9875e36f7d526ddc11edea9a3e509dc202fe8d2a8f40ef3bfb045df47291c863ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45c999fa99eec37645ef908b290ac214a713706ba1b49da90d7963bbd139e0c00f3f85c654dfe79e4bb1d06039fc5b46a1c239ec85a08aa88b73c0bed4b9fea179097eb5017df960;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h423aa0c8f32f5bacb16f236ef49f9bd6641ab8b5c2524bca9d5f579b558887e8000a6e554b7fb53fb627a819431229cf673f078491c8d026cf8d3d0e666d2df00fe653ce715cdb12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd908745b2e7032ee248676e2e9bfa787cd0c370f7b9c531ee3deead6d7d8fc5d38928aa5c098727cfc707cb8d239350137c574144e598cefc5bf4323f130d3a38df7c675007d3d4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb071e7e8f1c5dccfd99fdceb91905b5f9b95ae6a2478e554ba95cdaefa4ccdb7a87b8e444b5f10e09f202756cba37436610753a6e8fd8e5bf93a3a445213f5799b8134b7411320fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b73c0e0640feae43a4c64e61abb8e2f10f7120878e60f3049d5a2a0c95c156b39400b1686cc71c5cc812cbaf647a7c201236b2dc2a61fc26f6af79cd346dafea09c22b1d584110;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he695d8587f21ed6ac1db2e0657a3ccae1c93d997b569b276a57e1c71fe6ecef7464b9aede0654e2960ef6e1f3b6f6b33415bdb70de8332df91c5e8d3f1855d75f215f39b0a3ee3d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1db923af3382fd9ac9ee733c4460d120aac84381bd3b3fae38396cc5d9d541a45e2e86c0131abf2f833f36aeb70159ee9d68c5c6b27d63c42d13f611270e2a1e264ec5d738687a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf6df590e31c8e320559c8bc014669dd46ef4ddced5fbde8d1da5f1783326189000819762a4c35da4e8b11ec4713b22f384eb148fe32566558f523c4730232428dc29451e9c5fb71;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab8a6211111d73f148f02a6baca5b93894b3b11df31a042dcaf93d2792fe66cc768dbd3c99ddef64e8ec2c85e2262e8f177dced11ced15f5deb99ee45ecb61e66938e7ae67d279;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h644abcc25792d0cbfb7701e86c7b88a5b3e6831461a8df9b895bbf6e9b523a7438d5fe98858f417458a508342180cab3b07fa3627edc8206e769d6ce811c773fec03fd111f2bc9b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h781ce1384b78a3e93dac8e6969020746f4fc1110a7bef7dd58f08bdec9993b059d179c90e6ff021c9187eb183dd88be0343e0b150e8f0af5711bc4a9ef7371aacf2a3f95e0239a38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he11878620a1ce67e6f05669a24f0901732b6d62b117ade6b985b0c99bee9bc0fb7f7d558418045395fb96ccce12b9a523c07ae9e1d02018fc57c2c6759187aa62c0c98e98710f884;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb577ef8fe6ff0e10fc89b0fc67e9d018b37ed1e1ebb1dbd1900088c06e306ffd2abf2b0ec6a15db419c06759eb7e7fc38f8b016eabbc1bfe2edaae84da6b128a793a40159de5af28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fa6aa7c1d1b654a30abd4e6439c288150745e5319f06e197f31ba3c601f2820a1898c595e86073c1ef375303205178d341ea3708f40ef9e8ba4487274fb2b378bd622ececc03dbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h719de517808f31644b58dc134400b47c39117bbf6ec9a22e9bea93023eed06db5147b6be80775e18ba17ea8db929a622308ef44cb276043508d4a0c616f4b8a54cacee7a3b336912;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e299bb908b94d18a6a547c99b932c77fc8f52a16973c9433d55f1b20c3bb7d7bc340571819106d9263e825bb68148515d194d95ed5a7c66b1c52d2a2c0104fc7fd931b1387877b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48c75033a6328106e155dd8eb54a4f4a63d3a8565c193b52dd0bc303acf57c3edce88a5000e294e785f9feb33ff716ffbb129704e7055191d36919855b7a3d3e40d85b3a7f5a259a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb705661e9b20bf7f466ec30b830cfc661f7b48e41960a457ba67cc7aab90a34c4b5e77177b254624483537d920b256b467c10a402720be82534d9cacd80388ce066480e9d4fb4d02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0e7f24a2fa558282d3b2354f1e7407f50f75174f81d3592ec92c74d7d6daed43b12f423736be28cbe0f7f57885f39f1ae2f4d7ee5774045c98b909955a811921471f72be8a69b05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d2e63c7b1abd0c1d30037654ec29b49da61a2e9db4750ece3aa3d8e280f1b19770024fecc136f40a86d28652d5dd1d1c6998fc33ee6d38b6c3026abb426c92663a8c83c3f66d768;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h264871a6baeca770f006f3cf8fcc12f047f30e0a96f794e2093867921198f00932a7f220c3c65f60d00f3b926af905db645fc6cbfbb9a14eaf4ae1004082d3573ecd8785353dbd5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h868010f2952bccdb495b3cf42a4bc8bf5c8ccdb55cf93a85a75d40a03210449760bcbfd05453909db7de4a1afd8898a3be4008612009677c254306b2abb8eab247d0fbbada547e67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3216eedebd2bc0dcfd1326b0f545c74aee20413877c4ca27f55e7c76f85bcfd0eeb447708a6d9e65b57c6062971304ac4b13bca09681741017f988907c26f09bb9d2c7d9d187a31;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d6dafb4f6bff47a4ce935410ea947339c888215d8550e850c450e85291b0ef44535ac2665f8193602210323547e1d3c6c166822931d575b766bc22a1fe184cf80dacd8b538c74c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had67a4bf7dd0414c27f447d8534a7dd858ad85100582c1696cb903e6c72a9d8c1bbc0f549a6207f25f641f18d737af13554cd55a642dde0d007c63425633ba5cbdb601a74f4b6f3c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8f2a90b2db6c2426a28c3feefc90a7765d1fe63739b45e55f21d52999fcd2e723a7ec28151ca29095832b72b0a8a27d4bdfebbc2d0c1ef6e14e40ade73d690c0663045a785d054b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7235a221d57912ec1e01ef5919e2085cc37062a85c60962bdc9c7171de7aa54e260485300600e69525ac316635f5863330c232b081483583e78646a453c296eb3e5b7e31fd052b0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h335f3590758dd880e130f1f025232de7b07f95443adae6d91b498b36cc5186d1cd01dbc8f3d6e230249105a7a1cc719ab2273519e192e4f34720eea90e5f4760c13895726f6d9ba7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heabefe28904423050e4c1a50909407bdd848e0615214b33f30bc79eb35e3b024df86543c0eec6c91bd26e3d512bd2f2eeed02e050ff834db7e5dceb9ed6c56247540bb9b380a8461;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8e158b9eaea3df88ec070a93fed1ca686a5451bd336db5597b96f9ee87d3395bda93dfebb4a4100e286e4b2002833adf77652b4428e510d9c6a27bf455a7bb267853c07952622b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5775c75fb800661c1c76968f66ba5c02c774212c6fa8fdb2daf3ca933bc3ed3d77963ec4ebf5e9228397d4a8234015cb68517598f614eeb33d1d7f14007430f426feb231f1a87269;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a99b2b9f2597eedf066bc2432d265c12b307a1d8b6fb5b3ce538950d0753dcafa9b9858d87c9f60268d94cb2f5112572141b22a9d4555805036fae626089afa394a4bd0d1ad24df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6ff95e3887370da4b546ae42d0e9cec5c5abff2e78d0fe7e35849820606aeb83f70a40f97db97db32cbef0f44451c10f3a5edf818e1200df41c836244a408763214b21f3eeb53b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1424930c6476858abb5ffa771942b898ecaa3261aa09660ee9511bd29d5f0c9637079a255620316f0cb25c89206a42604859830d08cb5ff2338d8151e0153a31d3698e30393f846;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h963a703bdab269f291e8b047c66e86f317362bb2f13374571ba1df8f589947121dd912e83f32d088fcc2885a3d1ef31f6ed7279b95312cd2e71ff2cc0363af0766c877ca746485b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59bea286ec240440906ab2a019d7dbd1921069282ea3dd51db1eaa0aed806b05ad36915c4b0fa0848479a4535ad10a9708790fea2c86875394b87d1d490423eed6db089d0c95772c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50eb2aba2fb847cb996141546969e78a45ae3869212c59aff3e5d9878d2e96a57f1f705df0c3007c3977e1be2e9734dd1445de310abf7bbf78ac8bb77383835f438fe412cec47efa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff8121f23463cba329283ff6ce5c785b115acff365dbd15505d91899c411e581bf133a5883c77ba180ee61b19ea779081039837001bd8e07437bbdb8f4a59fce85a897e87e93de8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc008dc18b7224faa139e2bc4f0669df61d63a3234997db142f6e9426d0f29725eec3903462fae70606ce56e47bc5b42287e13f56c2b07eba0b07f43ac9a0838726539da2d4b8964;
        #1
        $finish();
    end
endmodule
