module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    compressor_CLA54_64 compressor_CLA54_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
        src32 <= 54'h0;
        src33 <= 54'h0;
        src34 <= 54'h0;
        src35 <= 54'h0;
        src36 <= 54'h0;
        src37 <= 54'h0;
        src38 <= 54'h0;
        src39 <= 54'h0;
        src40 <= 54'h0;
        src41 <= 54'h0;
        src42 <= 54'h0;
        src43 <= 54'h0;
        src44 <= 54'h0;
        src45 <= 54'h0;
        src46 <= 54'h0;
        src47 <= 54'h0;
        src48 <= 54'h0;
        src49 <= 54'h0;
        src50 <= 54'h0;
        src51 <= 54'h0;
        src52 <= 54'h0;
        src53 <= 54'h0;
        src54 <= 54'h0;
        src55 <= 54'h0;
        src56 <= 54'h0;
        src57 <= 54'h0;
        src58 <= 54'h0;
        src59 <= 54'h0;
        src60 <= 54'h0;
        src61 <= 54'h0;
        src62 <= 54'h0;
        src63 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA54_64(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    input [53:0]src32,
    input [53:0]src33,
    input [53:0]src34,
    input [53:0]src35,
    input [53:0]src36,
    input [53:0]src37,
    input [53:0]src38,
    input [53:0]src39,
    input [53:0]src40,
    input [53:0]src41,
    input [53:0]src42,
    input [53:0]src43,
    input [53:0]src44,
    input [53:0]src45,
    input [53:0]src46,
    input [53:0]src47,
    input [53:0]src48,
    input [53:0]src49,
    input [53:0]src50,
    input [53:0]src51,
    input [53:0]src52,
    input [53:0]src53,
    input [53:0]src54,
    input [53:0]src55,
    input [53:0]src56,
    input [53:0]src57,
    input [53:0]src58,
    input [53:0]src59,
    input [53:0]src60,
    input [53:0]src61,
    input [53:0]src62,
    input [53:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [0:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [0:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [0:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], 1'h0, comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], 1'h0, comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      input wire [53:0] src32,
      input wire [53:0] src33,
      input wire [53:0] src34,
      input wire [53:0] src35,
      input wire [53:0] src36,
      input wire [53:0] src37,
      input wire [53:0] src38,
      input wire [53:0] src39,
      input wire [53:0] src40,
      input wire [53:0] src41,
      input wire [53:0] src42,
      input wire [53:0] src43,
      input wire [53:0] src44,
      input wire [53:0] src45,
      input wire [53:0] src46,
      input wire [53:0] src47,
      input wire [53:0] src48,
      input wire [53:0] src49,
      input wire [53:0] src50,
      input wire [53:0] src51,
      input wire [53:0] src52,
      input wire [53:0] src53,
      input wire [53:0] src54,
      input wire [53:0] src55,
      input wire [53:0] src56,
      input wire [53:0] src57,
      input wire [53:0] src58,
      input wire [53:0] src59,
      input wire [53:0] src60,
      input wire [53:0] src61,
      input wire [53:0] src62,
      input wire [53:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [0:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [0:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [0:0] dst68,
      output wire [0:0] dst69);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [53:0] stage0_32;
   wire [53:0] stage0_33;
   wire [53:0] stage0_34;
   wire [53:0] stage0_35;
   wire [53:0] stage0_36;
   wire [53:0] stage0_37;
   wire [53:0] stage0_38;
   wire [53:0] stage0_39;
   wire [53:0] stage0_40;
   wire [53:0] stage0_41;
   wire [53:0] stage0_42;
   wire [53:0] stage0_43;
   wire [53:0] stage0_44;
   wire [53:0] stage0_45;
   wire [53:0] stage0_46;
   wire [53:0] stage0_47;
   wire [53:0] stage0_48;
   wire [53:0] stage0_49;
   wire [53:0] stage0_50;
   wire [53:0] stage0_51;
   wire [53:0] stage0_52;
   wire [53:0] stage0_53;
   wire [53:0] stage0_54;
   wire [53:0] stage0_55;
   wire [53:0] stage0_56;
   wire [53:0] stage0_57;
   wire [53:0] stage0_58;
   wire [53:0] stage0_59;
   wire [53:0] stage0_60;
   wire [53:0] stage0_61;
   wire [53:0] stage0_62;
   wire [53:0] stage0_63;
   wire [16:0] stage1_0;
   wire [19:0] stage1_1;
   wire [24:0] stage1_2;
   wire [23:0] stage1_3;
   wire [32:0] stage1_4;
   wire [35:0] stage1_5;
   wire [18:0] stage1_6;
   wire [24:0] stage1_7;
   wire [30:0] stage1_8;
   wire [17:0] stage1_9;
   wire [25:0] stage1_10;
   wire [28:0] stage1_11;
   wire [20:0] stage1_12;
   wire [29:0] stage1_13;
   wire [23:0] stage1_14;
   wire [42:0] stage1_15;
   wire [23:0] stage1_16;
   wire [17:0] stage1_17;
   wire [33:0] stage1_18;
   wire [20:0] stage1_19;
   wire [19:0] stage1_20;
   wire [25:0] stage1_21;
   wire [22:0] stage1_22;
   wire [21:0] stage1_23;
   wire [31:0] stage1_24;
   wire [24:0] stage1_25;
   wire [31:0] stage1_26;
   wire [23:0] stage1_27;
   wire [17:0] stage1_28;
   wire [25:0] stage1_29;
   wire [34:0] stage1_30;
   wire [33:0] stage1_31;
   wire [18:0] stage1_32;
   wire [45:0] stage1_33;
   wire [18:0] stage1_34;
   wire [27:0] stage1_35;
   wire [33:0] stage1_36;
   wire [24:0] stage1_37;
   wire [23:0] stage1_38;
   wire [30:0] stage1_39;
   wire [38:0] stage1_40;
   wire [19:0] stage1_41;
   wire [20:0] stage1_42;
   wire [22:0] stage1_43;
   wire [21:0] stage1_44;
   wire [31:0] stage1_45;
   wire [29:0] stage1_46;
   wire [33:0] stage1_47;
   wire [17:0] stage1_48;
   wire [23:0] stage1_49;
   wire [42:0] stage1_50;
   wire [47:0] stage1_51;
   wire [21:0] stage1_52;
   wire [40:0] stage1_53;
   wire [16:0] stage1_54;
   wire [37:0] stage1_55;
   wire [20:0] stage1_56;
   wire [40:0] stage1_57;
   wire [14:0] stage1_58;
   wire [34:0] stage1_59;
   wire [22:0] stage1_60;
   wire [20:0] stage1_61;
   wire [23:0] stage1_62;
   wire [34:0] stage1_63;
   wire [13:0] stage1_64;
   wire [5:0] stage1_65;
   wire [5:0] stage2_0;
   wire [6:0] stage2_1;
   wire [13:0] stage2_2;
   wire [8:0] stage2_3;
   wire [22:0] stage2_4;
   wire [9:0] stage2_5;
   wire [10:0] stage2_6;
   wire [12:0] stage2_7;
   wire [10:0] stage2_8;
   wire [19:0] stage2_9;
   wire [9:0] stage2_10;
   wire [12:0] stage2_11;
   wire [9:0] stage2_12;
   wire [9:0] stage2_13;
   wire [14:0] stage2_14;
   wire [13:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [19:0] stage2_18;
   wire [8:0] stage2_19;
   wire [8:0] stage2_20;
   wire [21:0] stage2_21;
   wire [10:0] stage2_22;
   wire [20:0] stage2_23;
   wire [9:0] stage2_24;
   wire [12:0] stage2_25;
   wire [18:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [9:0] stage2_30;
   wire [16:0] stage2_31;
   wire [11:0] stage2_32;
   wire [15:0] stage2_33;
   wire [15:0] stage2_34;
   wire [10:0] stage2_35;
   wire [18:0] stage2_36;
   wire [16:0] stage2_37;
   wire [12:0] stage2_38;
   wire [16:0] stage2_39;
   wire [11:0] stage2_40;
   wire [12:0] stage2_41;
   wire [13:0] stage2_42;
   wire [9:0] stage2_43;
   wire [14:0] stage2_44;
   wire [11:0] stage2_45;
   wire [17:0] stage2_46;
   wire [21:0] stage2_47;
   wire [12:0] stage2_48;
   wire [17:0] stage2_49;
   wire [10:0] stage2_50;
   wire [16:0] stage2_51;
   wire [18:0] stage2_52;
   wire [12:0] stage2_53;
   wire [14:0] stage2_54;
   wire [18:0] stage2_55;
   wire [12:0] stage2_56;
   wire [12:0] stage2_57;
   wire [17:0] stage2_58;
   wire [12:0] stage2_59;
   wire [12:0] stage2_60;
   wire [11:0] stage2_61;
   wire [17:0] stage2_62;
   wire [16:0] stage2_63;
   wire [5:0] stage2_64;
   wire [9:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [4:0] stage3_2;
   wire [5:0] stage3_3;
   wire [14:0] stage3_4;
   wire [8:0] stage3_5;
   wire [4:0] stage3_6;
   wire [13:0] stage3_7;
   wire [6:0] stage3_8;
   wire [10:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [4:0] stage3_12;
   wire [7:0] stage3_13;
   wire [3:0] stage3_14;
   wire [5:0] stage3_15;
   wire [5:0] stage3_16;
   wire [7:0] stage3_17;
   wire [5:0] stage3_18;
   wire [7:0] stage3_19;
   wire [4:0] stage3_20;
   wire [6:0] stage3_21;
   wire [6:0] stage3_22;
   wire [4:0] stage3_23;
   wire [5:0] stage3_24;
   wire [7:0] stage3_25;
   wire [5:0] stage3_26;
   wire [4:0] stage3_27;
   wire [4:0] stage3_28;
   wire [11:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [14:0] stage3_33;
   wire [8:0] stage3_34;
   wire [3:0] stage3_35;
   wire [5:0] stage3_36;
   wire [6:0] stage3_37;
   wire [6:0] stage3_38;
   wire [5:0] stage3_39;
   wire [6:0] stage3_40;
   wire [6:0] stage3_41;
   wire [5:0] stage3_42;
   wire [7:0] stage3_43;
   wire [7:0] stage3_44;
   wire [4:0] stage3_45;
   wire [5:0] stage3_46;
   wire [8:0] stage3_47;
   wire [12:0] stage3_48;
   wire [5:0] stage3_49;
   wire [10:0] stage3_50;
   wire [7:0] stage3_51;
   wire [10:0] stage3_52;
   wire [6:0] stage3_53;
   wire [5:0] stage3_54;
   wire [5:0] stage3_55;
   wire [10:0] stage3_56;
   wire [7:0] stage3_57;
   wire [3:0] stage3_58;
   wire [13:0] stage3_59;
   wire [5:0] stage3_60;
   wire [9:0] stage3_61;
   wire [3:0] stage3_62;
   wire [9:0] stage3_63;
   wire [4:0] stage3_64;
   wire [6:0] stage3_65;
   wire [5:0] stage3_66;
   wire [0:0] stage3_67;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [0:0] stage4_2;
   wire [1:0] stage4_3;
   wire [5:0] stage4_4;
   wire [2:0] stage4_5;
   wire [3:0] stage4_6;
   wire [5:0] stage4_7;
   wire [3:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [3:0] stage4_11;
   wire [3:0] stage4_12;
   wire [1:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [6:0] stage4_18;
   wire [2:0] stage4_19;
   wire [2:0] stage4_20;
   wire [3:0] stage4_21;
   wire [1:0] stage4_22;
   wire [2:0] stage4_23;
   wire [2:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [5:0] stage4_27;
   wire [0:0] stage4_28;
   wire [5:0] stage4_29;
   wire [2:0] stage4_30;
   wire [1:0] stage4_31;
   wire [2:0] stage4_32;
   wire [5:0] stage4_33;
   wire [2:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [5:0] stage4_37;
   wire [6:0] stage4_38;
   wire [0:0] stage4_39;
   wire [2:0] stage4_40;
   wire [2:0] stage4_41;
   wire [2:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [1:0] stage4_45;
   wire [2:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [2:0] stage4_49;
   wire [3:0] stage4_50;
   wire [4:0] stage4_51;
   wire [3:0] stage4_52;
   wire [2:0] stage4_53;
   wire [2:0] stage4_54;
   wire [3:0] stage4_55;
   wire [5:0] stage4_56;
   wire [2:0] stage4_57;
   wire [2:0] stage4_58;
   wire [5:0] stage4_59;
   wire [2:0] stage4_60;
   wire [5:0] stage4_61;
   wire [2:0] stage4_62;
   wire [5:0] stage4_63;
   wire [2:0] stage4_64;
   wire [2:0] stage4_65;
   wire [2:0] stage4_66;
   wire [2:0] stage4_67;
   wire [0:0] stage4_68;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [1:0] stage5_3;
   wire [0:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [0:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [1:0] stage5_67;
   wire [0:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc7_3 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc17 (
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc18 (
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc19 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[18]}
   );
   gpc615_5 gpc20 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_5[19]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[4],stage1_6[6],stage1_5[11],stage1_4[19]}
   );
   gpc615_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_5[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[5],stage1_6[7],stage1_5[12],stage1_4[20]}
   );
   gpc615_5 gpc22 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[21]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[6],stage1_6[8],stage1_5[13],stage1_4[21]}
   );
   gpc615_5 gpc23 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39]},
      {stage0_5[22]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[7],stage1_6[9],stage1_5[14],stage1_4[22]}
   );
   gpc615_5 gpc24 (
      {stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_5[23]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[8],stage1_6[10],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc25 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[6],stage1_7[9],stage1_6[11],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[7],stage1_7[10],stage1_6[12],stage1_5[17]}
   );
   gpc615_5 gpc27 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40]},
      {stage0_7[12]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[8],stage1_7[11],stage1_6[13]}
   );
   gpc615_5 gpc28 (
      {stage0_6[41], stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45]},
      {stage0_7[13]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[3],stage1_8[9],stage1_7[12],stage1_6[14]}
   );
   gpc615_5 gpc29 (
      {stage0_6[46], stage0_6[47], stage0_6[48], stage0_6[49], stage0_6[50]},
      {stage0_7[14]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[4],stage1_8[10],stage1_7[13],stage1_6[15]}
   );
   gpc606_5 gpc30 (
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[5],stage1_8[11],stage1_7[14]}
   );
   gpc606_5 gpc31 (
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[6],stage1_8[12],stage1_7[15]}
   );
   gpc606_5 gpc32 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31], stage0_7[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[7],stage1_8[13],stage1_7[16]}
   );
   gpc606_5 gpc33 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37], stage0_7[38]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[8],stage1_8[14],stage1_7[17]}
   );
   gpc615_5 gpc34 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43]},
      {stage0_8[18]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[7],stage1_9[9],stage1_8[15],stage1_7[18]}
   );
   gpc615_5 gpc35 (
      {stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48]},
      {stage0_8[19]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[8],stage1_9[10],stage1_8[16],stage1_7[19]}
   );
   gpc606_5 gpc36 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[6],stage1_10[9],stage1_9[11],stage1_8[17]}
   );
   gpc606_5 gpc37 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[7],stage1_10[10],stage1_9[12],stage1_8[18]}
   );
   gpc606_5 gpc38 (
      {stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[8],stage1_10[11],stage1_9[13],stage1_8[19]}
   );
   gpc606_5 gpc39 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[9],stage1_10[12],stage1_9[14],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[4],stage1_11[10],stage1_10[13],stage1_9[15]}
   );
   gpc606_5 gpc41 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[5],stage1_11[11],stage1_10[14],stage1_9[16]}
   );
   gpc606_5 gpc42 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[6],stage1_11[12],stage1_10[15],stage1_9[17]}
   );
   gpc615_5 gpc43 (
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28]},
      {stage0_11[18]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[7],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc44 (
      {stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage0_11[19]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[8],stage1_11[14],stage1_10[17]}
   );
   gpc615_5 gpc45 (
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38]},
      {stage0_11[20]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[9],stage1_11[15],stage1_10[18]}
   );
   gpc615_5 gpc46 (
      {stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_11[21]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[10],stage1_11[16],stage1_10[19]}
   );
   gpc615_5 gpc47 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[22]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[7],stage1_12[11],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc48 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[30]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[5],stage1_13[8],stage1_12[12],stage1_11[18]}
   );
   gpc615_5 gpc49 (
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_12[31]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[6],stage1_13[9],stage1_12[13],stage1_11[19]}
   );
   gpc615_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37]},
      {stage0_12[32]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[7],stage1_13[10],stage1_12[14],stage1_11[20]}
   );
   gpc615_5 gpc51 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[33]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[8],stage1_13[11],stage1_12[15],stage1_11[21]}
   );
   gpc615_5 gpc52 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[34]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[9],stage1_13[12],stage1_12[16],stage1_11[22]}
   );
   gpc606_5 gpc53 (
      {stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[5],stage1_14[10],stage1_13[13],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[6],stage1_14[11],stage1_13[14],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[7],stage1_14[12],stage1_13[15],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[8],stage1_14[13],stage1_13[16]}
   );
   gpc606_5 gpc57 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[9],stage1_14[14],stage1_13[17]}
   );
   gpc606_5 gpc58 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[2],stage1_16[5],stage1_15[10],stage1_14[15]}
   );
   gpc606_5 gpc59 (
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[3],stage1_16[6],stage1_15[11],stage1_14[16]}
   );
   gpc606_5 gpc60 (
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[4],stage1_16[7],stage1_15[12],stage1_14[17]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[12]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[5],stage1_16[8],stage1_15[13],stage1_14[18]}
   );
   gpc615_5 gpc62 (
      {stage0_14[41], stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45]},
      {stage0_15[13]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[6],stage1_16[9],stage1_15[14],stage1_14[19]}
   );
   gpc615_5 gpc63 (
      {stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[14]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[7],stage1_16[10],stage1_15[15],stage1_14[20]}
   );
   gpc615_5 gpc64 (
      {stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18], stage0_15[19]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[8],stage1_16[11],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[9],stage1_16[12],stage1_15[17]}
   );
   gpc615_5 gpc66 (
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage0_16[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[8],stage1_17[10],stage1_16[13],stage1_15[18]}
   );
   gpc606_5 gpc67 (
      {stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[3],stage1_18[9],stage1_17[11],stage1_16[14]}
   );
   gpc606_5 gpc68 (
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[4],stage1_18[10],stage1_17[12]}
   );
   gpc606_5 gpc69 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[2],stage1_19[5],stage1_18[11],stage1_17[13]}
   );
   gpc606_5 gpc70 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[3],stage1_19[6],stage1_18[12],stage1_17[14]}
   );
   gpc606_5 gpc71 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[4],stage1_19[7],stage1_18[13],stage1_17[15]}
   );
   gpc606_5 gpc72 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[5],stage1_19[8],stage1_18[14],stage1_17[16]}
   );
   gpc606_5 gpc73 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[6],stage1_19[9],stage1_18[15],stage1_17[17]}
   );
   gpc606_5 gpc74 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[6],stage1_20[7],stage1_19[10],stage1_18[16]}
   );
   gpc606_5 gpc75 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[7],stage1_20[8],stage1_19[11],stage1_18[17]}
   );
   gpc606_5 gpc76 (
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[8],stage1_20[9],stage1_19[12],stage1_18[18]}
   );
   gpc606_5 gpc77 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[9],stage1_20[10],stage1_19[13],stage1_18[19]}
   );
   gpc606_5 gpc78 (
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[10],stage1_20[11],stage1_19[14],stage1_18[20]}
   );
   gpc606_5 gpc79 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[11],stage1_20[12],stage1_19[15],stage1_18[21]}
   );
   gpc606_5 gpc80 (
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[6],stage1_21[12],stage1_20[13],stage1_19[16]}
   );
   gpc615_5 gpc81 (
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46]},
      {stage0_20[36]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[7],stage1_21[13],stage1_20[14],stage1_19[17]}
   );
   gpc615_5 gpc82 (
      {stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51]},
      {stage0_20[37]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[8],stage1_21[14],stage1_20[15],stage1_19[18]}
   );
   gpc615_5 gpc83 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[18]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[3],stage1_22[9],stage1_21[15],stage1_20[16]}
   );
   gpc615_5 gpc84 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[4],stage1_22[10],stage1_21[16],stage1_20[17]}
   );
   gpc615_5 gpc85 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[20]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[5],stage1_22[11],stage1_21[17],stage1_20[18]}
   );
   gpc606_5 gpc86 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[3],stage1_23[6],stage1_22[12],stage1_21[18]}
   );
   gpc606_5 gpc87 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[4],stage1_23[7],stage1_22[13],stage1_21[19]}
   );
   gpc606_5 gpc88 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[5],stage1_23[8],stage1_22[14],stage1_21[20]}
   );
   gpc606_5 gpc89 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[6],stage1_23[9],stage1_22[15],stage1_21[21]}
   );
   gpc606_5 gpc90 (
      {stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49], stage0_21[50]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[7],stage1_23[10],stage1_22[16],stage1_21[22]}
   );
   gpc606_5 gpc91 (
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[8],stage1_23[11],stage1_22[17]}
   );
   gpc606_5 gpc92 (
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[9],stage1_23[12],stage1_22[18]}
   );
   gpc606_5 gpc93 (
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[10],stage1_23[13],stage1_22[19]}
   );
   gpc606_5 gpc94 (
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[11],stage1_23[14],stage1_22[20]}
   );
   gpc606_5 gpc95 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[12],stage1_23[15],stage1_22[21]}
   );
   gpc606_5 gpc96 (
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[13],stage1_23[16],stage1_22[22]}
   );
   gpc615_5 gpc97 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34]},
      {stage0_24[36]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[6],stage1_25[11],stage1_24[14],stage1_23[17]}
   );
   gpc615_5 gpc98 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage0_24[37]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[7],stage1_25[12],stage1_24[15],stage1_23[18]}
   );
   gpc615_5 gpc99 (
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44]},
      {stage0_24[38]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[8],stage1_25[13],stage1_24[16],stage1_23[19]}
   );
   gpc615_5 gpc100 (
      {stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49]},
      {stage0_24[39]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[9],stage1_25[14],stage1_24[17],stage1_23[20]}
   );
   gpc615_5 gpc101 (
      {stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], 1'b0},
      {stage0_24[40]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[10],stage1_25[15],stage1_24[18],stage1_23[21]}
   );
   gpc606_5 gpc102 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[0],stage1_27[5],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc103 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[1],stage1_27[6],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc104 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[2],stage1_27[7],stage1_26[13],stage1_25[18]}
   );
   gpc2135_5 gpc105 (
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4]},
      {stage0_27[18], stage0_27[19], stage0_27[20]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1]},
      {stage1_30[0],stage1_29[3],stage1_28[3],stage1_27[8],stage1_26[14]}
   );
   gpc2135_5 gpc106 (
      {stage0_26[5], stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9]},
      {stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage0_28[1]},
      {stage0_29[2], stage0_29[3]},
      {stage1_30[1],stage1_29[4],stage1_28[4],stage1_27[9],stage1_26[15]}
   );
   gpc2135_5 gpc107 (
      {stage0_26[10], stage0_26[11], stage0_26[12], stage0_26[13], stage0_26[14]},
      {stage0_27[24], stage0_27[25], stage0_27[26]},
      {stage0_28[2]},
      {stage0_29[4], stage0_29[5]},
      {stage1_30[2],stage1_29[5],stage1_28[5],stage1_27[10],stage1_26[16]}
   );
   gpc2135_5 gpc108 (
      {stage0_26[15], stage0_26[16], stage0_26[17], stage0_26[18], stage0_26[19]},
      {stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage0_28[3]},
      {stage0_29[6], stage0_29[7]},
      {stage1_30[3],stage1_29[6],stage1_28[6],stage1_27[11],stage1_26[17]}
   );
   gpc615_5 gpc109 (
      {stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24]},
      {stage0_27[30]},
      {stage0_28[4], stage0_28[5], stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9]},
      {stage1_30[4],stage1_29[7],stage1_28[7],stage1_27[12],stage1_26[18]}
   );
   gpc615_5 gpc110 (
      {stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage0_27[31]},
      {stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15]},
      {stage1_30[5],stage1_29[8],stage1_28[8],stage1_27[13],stage1_26[19]}
   );
   gpc615_5 gpc111 (
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34]},
      {stage0_27[32]},
      {stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage1_30[6],stage1_29[9],stage1_28[9],stage1_27[14],stage1_26[20]}
   );
   gpc615_5 gpc112 (
      {stage0_26[35], stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39]},
      {stage0_27[33]},
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27]},
      {stage1_30[7],stage1_29[10],stage1_28[10],stage1_27[15],stage1_26[21]}
   );
   gpc615_5 gpc113 (
      {stage0_26[40], stage0_26[41], stage0_26[42], stage0_26[43], stage0_26[44]},
      {stage0_27[34]},
      {stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33]},
      {stage1_30[8],stage1_29[11],stage1_28[11],stage1_27[16],stage1_26[22]}
   );
   gpc615_5 gpc114 (
      {stage0_27[35], stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39]},
      {stage0_28[34]},
      {stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13]},
      {stage1_31[0],stage1_30[9],stage1_29[12],stage1_28[12],stage1_27[17]}
   );
   gpc615_5 gpc115 (
      {stage0_27[40], stage0_27[41], stage0_27[42], stage0_27[43], stage0_27[44]},
      {stage0_28[35]},
      {stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19]},
      {stage1_31[1],stage1_30[10],stage1_29[13],stage1_28[13],stage1_27[18]}
   );
   gpc615_5 gpc116 (
      {stage0_27[45], stage0_27[46], stage0_27[47], stage0_27[48], stage0_27[49]},
      {stage0_28[36]},
      {stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25]},
      {stage1_31[2],stage1_30[11],stage1_29[14],stage1_28[14],stage1_27[19]}
   );
   gpc606_5 gpc117 (
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[3],stage1_30[12],stage1_29[15],stage1_28[15]}
   );
   gpc606_5 gpc118 (
      {stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[4],stage1_30[13],stage1_29[16],stage1_28[16]}
   );
   gpc606_5 gpc119 (
      {stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], 1'b0},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[5],stage1_30[14],stage1_29[17],stage1_28[17]}
   );
   gpc606_5 gpc120 (
      {stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[6],stage1_30[15],stage1_29[18]}
   );
   gpc606_5 gpc121 (
      {stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[7],stage1_30[16],stage1_29[19]}
   );
   gpc606_5 gpc122 (
      {stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[8],stage1_30[17],stage1_29[20]}
   );
   gpc606_5 gpc123 (
      {stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[9],stage1_30[18],stage1_29[21]}
   );
   gpc606_5 gpc124 (
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[4],stage1_32[7],stage1_31[10],stage1_30[19]}
   );
   gpc606_5 gpc125 (
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[5],stage1_32[8],stage1_31[11],stage1_30[20]}
   );
   gpc606_5 gpc126 (
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[6],stage1_32[9],stage1_31[12],stage1_30[21]}
   );
   gpc606_5 gpc127 (
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[7],stage1_32[10],stage1_31[13],stage1_30[22]}
   );
   gpc606_5 gpc128 (
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[4],stage1_33[8],stage1_32[11],stage1_31[14]}
   );
   gpc606_5 gpc129 (
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[5],stage1_33[9],stage1_32[12],stage1_31[15]}
   );
   gpc606_5 gpc130 (
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[10],stage1_32[13]}
   );
   gpc606_5 gpc131 (
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[11],stage1_32[14]}
   );
   gpc606_5 gpc132 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[12],stage1_32[15]}
   );
   gpc606_5 gpc133 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[13],stage1_32[16]}
   );
   gpc615_5 gpc134 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52]},
      {stage0_33[12]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[14],stage1_32[17]}
   );
   gpc606_5 gpc135 (
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[15]}
   );
   gpc606_5 gpc136 (
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[16]}
   );
   gpc117_4 gpc137 (
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35], stage0_34[36]},
      {stage0_35[12]},
      {stage0_36[0]},
      {stage1_37[2],stage1_36[7],stage1_35[9],stage1_34[13]}
   );
   gpc117_4 gpc138 (
      {stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41], stage0_34[42], stage0_34[43]},
      {stage0_35[13]},
      {stage0_36[1]},
      {stage1_37[3],stage1_36[8],stage1_35[10],stage1_34[14]}
   );
   gpc117_4 gpc139 (
      {stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47], stage0_34[48], stage0_34[49], stage0_34[50]},
      {stage0_35[14]},
      {stage0_36[2]},
      {stage1_37[4],stage1_36[9],stage1_35[11],stage1_34[15]}
   );
   gpc606_5 gpc140 (
      {stage0_35[15], stage0_35[16], stage0_35[17], stage0_35[18], stage0_35[19], stage0_35[20]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[0],stage1_37[5],stage1_36[10],stage1_35[12]}
   );
   gpc606_5 gpc141 (
      {stage0_35[21], stage0_35[22], stage0_35[23], stage0_35[24], stage0_35[25], stage0_35[26]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[1],stage1_37[6],stage1_36[11],stage1_35[13]}
   );
   gpc606_5 gpc142 (
      {stage0_35[27], stage0_35[28], stage0_35[29], stage0_35[30], stage0_35[31], stage0_35[32]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[2],stage1_37[7],stage1_36[12],stage1_35[14]}
   );
   gpc615_5 gpc143 (
      {stage0_35[33], stage0_35[34], stage0_35[35], stage0_35[36], stage0_35[37]},
      {stage0_36[3]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[3],stage1_37[8],stage1_36[13],stage1_35[15]}
   );
   gpc615_5 gpc144 (
      {stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41], stage0_35[42]},
      {stage0_36[4]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[4],stage1_37[9],stage1_36[14],stage1_35[16]}
   );
   gpc606_5 gpc145 (
      {stage0_36[5], stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[5],stage1_38[5],stage1_37[10],stage1_36[15]}
   );
   gpc606_5 gpc146 (
      {stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[6],stage1_38[6],stage1_37[11],stage1_36[16]}
   );
   gpc606_5 gpc147 (
      {stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[7],stage1_38[7],stage1_37[12],stage1_36[17]}
   );
   gpc606_5 gpc148 (
      {stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[8],stage1_38[8],stage1_37[13],stage1_36[18]}
   );
   gpc606_5 gpc149 (
      {stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[9],stage1_38[9],stage1_37[14],stage1_36[19]}
   );
   gpc606_5 gpc150 (
      {stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[10],stage1_38[10],stage1_37[15],stage1_36[20]}
   );
   gpc606_5 gpc151 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[11],stage1_38[11],stage1_37[16]}
   );
   gpc606_5 gpc152 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[12],stage1_38[12],stage1_37[17]}
   );
   gpc606_5 gpc153 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[13],stage1_38[13],stage1_37[18]}
   );
   gpc615_5 gpc154 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[18]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[3],stage1_40[9],stage1_39[14],stage1_38[14]}
   );
   gpc615_5 gpc155 (
      {stage0_38[41], stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45]},
      {stage0_39[19]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[4],stage1_40[10],stage1_39[15],stage1_38[15]}
   );
   gpc606_5 gpc156 (
      {stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23], stage0_39[24], stage0_39[25]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[2],stage1_41[5],stage1_40[11],stage1_39[16]}
   );
   gpc606_5 gpc157 (
      {stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29], stage0_39[30], stage0_39[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[3],stage1_41[6],stage1_40[12],stage1_39[17]}
   );
   gpc606_5 gpc158 (
      {stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35], stage0_39[36], stage0_39[37]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[4],stage1_41[7],stage1_40[13],stage1_39[18]}
   );
   gpc615_5 gpc159 (
      {stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41], stage0_39[42]},
      {stage0_40[12]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[5],stage1_41[8],stage1_40[14],stage1_39[19]}
   );
   gpc1406_5 gpc160 (
      {stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17], stage0_40[18]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[4],stage1_42[6],stage1_41[9],stage1_40[15]}
   );
   gpc615_5 gpc161 (
      {stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage0_41[24]},
      {stage0_42[4], stage0_42[5], stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9]},
      {stage1_44[1],stage1_43[5],stage1_42[7],stage1_41[10],stage1_40[16]}
   );
   gpc615_5 gpc162 (
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28]},
      {stage0_41[25]},
      {stage0_42[10], stage0_42[11], stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15]},
      {stage1_44[2],stage1_43[6],stage1_42[8],stage1_41[11],stage1_40[17]}
   );
   gpc615_5 gpc163 (
      {stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_41[26]},
      {stage0_42[16], stage0_42[17], stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21]},
      {stage1_44[3],stage1_43[7],stage1_42[9],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc164 (
      {stage0_41[27], stage0_41[28], stage0_41[29], stage0_41[30], stage0_41[31], stage0_41[32]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[4],stage1_43[8],stage1_42[10],stage1_41[13]}
   );
   gpc606_5 gpc165 (
      {stage0_41[33], stage0_41[34], stage0_41[35], stage0_41[36], stage0_41[37], stage0_41[38]},
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage1_45[1],stage1_44[5],stage1_43[9],stage1_42[11],stage1_41[14]}
   );
   gpc606_5 gpc166 (
      {stage0_41[39], stage0_41[40], stage0_41[41], stage0_41[42], stage0_41[43], stage0_41[44]},
      {stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17], stage0_43[18]},
      {stage1_45[2],stage1_44[6],stage1_43[10],stage1_42[12],stage1_41[15]}
   );
   gpc606_5 gpc167 (
      {stage0_41[45], stage0_41[46], stage0_41[47], stage0_41[48], stage0_41[49], stage0_41[50]},
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23], stage0_43[24]},
      {stage1_45[3],stage1_44[7],stage1_43[11],stage1_42[13],stage1_41[16]}
   );
   gpc606_5 gpc168 (
      {stage0_42[22], stage0_42[23], stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[4],stage1_44[8],stage1_43[12],stage1_42[14]}
   );
   gpc606_5 gpc169 (
      {stage0_42[28], stage0_42[29], stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[5],stage1_44[9],stage1_43[13],stage1_42[15]}
   );
   gpc606_5 gpc170 (
      {stage0_42[34], stage0_42[35], stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[6],stage1_44[10],stage1_43[14],stage1_42[16]}
   );
   gpc606_5 gpc171 (
      {stage0_42[40], stage0_42[41], stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[7],stage1_44[11],stage1_43[15],stage1_42[17]}
   );
   gpc606_5 gpc172 (
      {stage0_42[46], stage0_42[47], stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[8],stage1_44[12],stage1_43[16],stage1_42[18]}
   );
   gpc615_5 gpc173 (
      {stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage0_44[30]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[5],stage1_45[9],stage1_44[13],stage1_43[17]}
   );
   gpc615_5 gpc174 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[31]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[6],stage1_45[10],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc175 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[32]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[7],stage1_45[11],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc176 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[33]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[8],stage1_45[12],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc177 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[34]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[9],stage1_45[13],stage1_44[17],stage1_43[21]}
   );
   gpc615_5 gpc178 (
      {stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53], 1'b0},
      {stage0_44[35]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[10],stage1_45[14],stage1_44[18],stage1_43[22]}
   );
   gpc606_5 gpc179 (
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[6],stage1_46[11],stage1_45[15],stage1_44[19]}
   );
   gpc606_5 gpc180 (
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[7],stage1_46[12],stage1_45[16],stage1_44[20]}
   );
   gpc606_5 gpc181 (
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[8],stage1_46[13],stage1_45[17],stage1_44[21]}
   );
   gpc615_5 gpc182 (
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40]},
      {stage0_46[18]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[3],stage1_47[9],stage1_46[14],stage1_45[18]}
   );
   gpc615_5 gpc183 (
      {stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage0_47[6]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[1],stage1_48[4],stage1_47[10],stage1_46[15]}
   );
   gpc615_5 gpc184 (
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28]},
      {stage0_47[7]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[2],stage1_48[5],stage1_47[11],stage1_46[16]}
   );
   gpc615_5 gpc185 (
      {stage0_46[29], stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33]},
      {stage0_47[8]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[3],stage1_48[6],stage1_47[12],stage1_46[17]}
   );
   gpc615_5 gpc186 (
      {stage0_46[34], stage0_46[35], stage0_46[36], stage0_46[37], stage0_46[38]},
      {stage0_47[9]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[4],stage1_48[7],stage1_47[13],stage1_46[18]}
   );
   gpc615_5 gpc187 (
      {stage0_46[39], stage0_46[40], stage0_46[41], stage0_46[42], stage0_46[43]},
      {stage0_47[10]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[5],stage1_48[8],stage1_47[14],stage1_46[19]}
   );
   gpc615_5 gpc188 (
      {stage0_47[11], stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15]},
      {stage0_48[30]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[5],stage1_49[6],stage1_48[9],stage1_47[15]}
   );
   gpc615_5 gpc189 (
      {stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19], stage0_47[20]},
      {stage0_48[31]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[6],stage1_49[7],stage1_48[10],stage1_47[16]}
   );
   gpc615_5 gpc190 (
      {stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_48[32]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[7],stage1_49[8],stage1_48[11],stage1_47[17]}
   );
   gpc615_5 gpc191 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[33]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[8],stage1_49[9],stage1_48[12],stage1_47[18]}
   );
   gpc615_5 gpc192 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[34]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[9],stage1_49[10],stage1_48[13],stage1_47[19]}
   );
   gpc615_5 gpc193 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[35]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[10],stage1_49[11],stage1_48[14],stage1_47[20]}
   );
   gpc606_5 gpc194 (
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[11],stage1_49[12],stage1_48[15]}
   );
   gpc606_5 gpc195 (
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[12],stage1_49[13],stage1_48[16]}
   );
   gpc606_5 gpc196 (
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[13],stage1_49[14],stage1_48[17]}
   );
   gpc606_5 gpc197 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[3],stage1_51[9],stage1_50[14],stage1_49[15]}
   );
   gpc615_5 gpc198 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46]},
      {stage0_50[18]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[4],stage1_51[10],stage1_50[15],stage1_49[16]}
   );
   gpc615_5 gpc199 (
      {stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage0_51[12]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[2],stage1_52[5],stage1_51[11],stage1_50[16]}
   );
   gpc615_5 gpc200 (
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28]},
      {stage0_51[13]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[3],stage1_52[6],stage1_51[12],stage1_50[17]}
   );
   gpc606_5 gpc201 (
      {stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17], stage0_51[18], stage0_51[19]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[2],stage1_53[4],stage1_52[7],stage1_51[13]}
   );
   gpc615_5 gpc202 (
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16]},
      {stage0_53[6]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[1],stage1_54[3],stage1_53[5],stage1_52[8]}
   );
   gpc615_5 gpc203 (
      {stage0_52[17], stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21]},
      {stage0_53[7]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[2],stage1_54[4],stage1_53[6],stage1_52[9]}
   );
   gpc615_5 gpc204 (
      {stage0_52[22], stage0_52[23], stage0_52[24], stage0_52[25], stage0_52[26]},
      {stage0_53[8]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[3],stage1_54[5],stage1_53[7],stage1_52[10]}
   );
   gpc615_5 gpc205 (
      {stage0_52[27], stage0_52[28], stage0_52[29], stage0_52[30], stage0_52[31]},
      {stage0_53[9]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[4],stage1_54[6],stage1_53[8],stage1_52[11]}
   );
   gpc615_5 gpc206 (
      {stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35], stage0_52[36]},
      {stage0_53[10]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[5],stage1_54[7],stage1_53[9],stage1_52[12]}
   );
   gpc615_5 gpc207 (
      {stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_53[11]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[6],stage1_54[8],stage1_53[10],stage1_52[13]}
   );
   gpc615_5 gpc208 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46]},
      {stage0_53[12]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[7],stage1_54[9],stage1_53[11],stage1_52[14]}
   );
   gpc615_5 gpc209 (
      {stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage0_54[42]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[7],stage1_55[8],stage1_54[10],stage1_53[12]}
   );
   gpc615_5 gpc210 (
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22]},
      {stage0_54[43]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[8],stage1_55[9],stage1_54[11],stage1_53[13]}
   );
   gpc615_5 gpc211 (
      {stage0_53[23], stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27]},
      {stage0_54[44]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[9],stage1_55[10],stage1_54[12],stage1_53[14]}
   );
   gpc606_5 gpc212 (
      {stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48], stage0_54[49], stage0_54[50]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[3],stage1_56[10],stage1_55[11],stage1_54[13]}
   );
   gpc606_5 gpc213 (
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[1],stage1_57[4],stage1_56[11],stage1_55[12]}
   );
   gpc606_5 gpc214 (
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[2],stage1_57[5],stage1_56[12],stage1_55[13]}
   );
   gpc606_5 gpc215 (
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[2],stage1_58[3],stage1_57[6],stage1_56[13]}
   );
   gpc606_5 gpc216 (
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[3],stage1_58[4],stage1_57[7],stage1_56[14]}
   );
   gpc606_5 gpc217 (
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[4],stage1_58[5],stage1_57[8],stage1_56[15]}
   );
   gpc606_5 gpc218 (
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[5],stage1_58[6],stage1_57[9],stage1_56[16]}
   );
   gpc606_5 gpc219 (
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[6],stage1_58[7],stage1_57[10],stage1_56[17]}
   );
   gpc606_5 gpc220 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[7],stage1_58[8],stage1_57[11],stage1_56[18]}
   );
   gpc606_5 gpc221 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[8],stage1_58[9],stage1_57[12],stage1_56[19]}
   );
   gpc606_5 gpc222 (
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[9],stage1_58[10],stage1_57[13],stage1_56[20]}
   );
   gpc606_5 gpc223 (
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[8],stage1_59[10],stage1_58[11],stage1_57[14]}
   );
   gpc606_5 gpc224 (
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[9],stage1_59[11],stage1_58[12],stage1_57[15]}
   );
   gpc606_5 gpc225 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[10],stage1_59[12],stage1_58[13],stage1_57[16]}
   );
   gpc606_5 gpc226 (
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[3],stage1_60[11],stage1_59[13],stage1_58[14]}
   );
   gpc606_5 gpc227 (
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[1],stage1_61[4],stage1_60[12],stage1_59[14]}
   );
   gpc606_5 gpc228 (
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage1_63[1],stage1_62[2],stage1_61[5],stage1_60[13],stage1_59[15]}
   );
   gpc606_5 gpc229 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage1_63[2],stage1_62[3],stage1_61[6],stage1_60[14],stage1_59[16]}
   );
   gpc606_5 gpc230 (
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[3],stage1_62[4],stage1_61[7],stage1_60[15]}
   );
   gpc606_5 gpc231 (
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[4],stage1_62[5],stage1_61[8],stage1_60[16]}
   );
   gpc606_5 gpc232 (
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[5],stage1_62[6],stage1_61[9],stage1_60[17]}
   );
   gpc606_5 gpc233 (
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[6],stage1_62[7],stage1_61[10],stage1_60[18]}
   );
   gpc606_5 gpc234 (
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[7],stage1_62[8],stage1_61[11],stage1_60[19]}
   );
   gpc606_5 gpc235 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[8],stage1_62[9],stage1_61[12],stage1_60[20]}
   );
   gpc606_5 gpc236 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[9],stage1_62[10],stage1_61[13],stage1_60[21]}
   );
   gpc606_5 gpc237 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[10],stage1_62[11],stage1_61[14],stage1_60[22]}
   );
   gpc606_5 gpc238 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[8],stage1_63[11],stage1_62[12],stage1_61[15]}
   );
   gpc606_5 gpc239 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[9],stage1_63[12],stage1_62[13],stage1_61[16]}
   );
   gpc606_5 gpc240 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[10],stage1_63[13],stage1_62[14],stage1_61[17]}
   );
   gpc606_5 gpc241 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[11],stage1_63[14],stage1_62[15],stage1_61[18]}
   );
   gpc606_5 gpc242 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[12],stage1_63[15],stage1_62[16],stage1_61[19]}
   );
   gpc606_5 gpc243 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[13],stage1_63[16],stage1_62[17],stage1_61[20]}
   );
   gpc1_1 gpc244 (
      {stage0_0[46]},
      {stage1_0[9]}
   );
   gpc1_1 gpc245 (
      {stage0_0[47]},
      {stage1_0[10]}
   );
   gpc1_1 gpc246 (
      {stage0_0[48]},
      {stage1_0[11]}
   );
   gpc1_1 gpc247 (
      {stage0_0[49]},
      {stage1_0[12]}
   );
   gpc1_1 gpc248 (
      {stage0_0[50]},
      {stage1_0[13]}
   );
   gpc1_1 gpc249 (
      {stage0_0[51]},
      {stage1_0[14]}
   );
   gpc1_1 gpc250 (
      {stage0_0[52]},
      {stage1_0[15]}
   );
   gpc1_1 gpc251 (
      {stage0_0[53]},
      {stage1_0[16]}
   );
   gpc1_1 gpc252 (
      {stage0_1[48]},
      {stage1_1[14]}
   );
   gpc1_1 gpc253 (
      {stage0_1[49]},
      {stage1_1[15]}
   );
   gpc1_1 gpc254 (
      {stage0_1[50]},
      {stage1_1[16]}
   );
   gpc1_1 gpc255 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc256 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc257 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc258 (
      {stage0_2[45]},
      {stage1_2[16]}
   );
   gpc1_1 gpc259 (
      {stage0_2[46]},
      {stage1_2[17]}
   );
   gpc1_1 gpc260 (
      {stage0_2[47]},
      {stage1_2[18]}
   );
   gpc1_1 gpc261 (
      {stage0_2[48]},
      {stage1_2[19]}
   );
   gpc1_1 gpc262 (
      {stage0_2[49]},
      {stage1_2[20]}
   );
   gpc1_1 gpc263 (
      {stage0_2[50]},
      {stage1_2[21]}
   );
   gpc1_1 gpc264 (
      {stage0_2[51]},
      {stage1_2[22]}
   );
   gpc1_1 gpc265 (
      {stage0_2[52]},
      {stage1_2[23]}
   );
   gpc1_1 gpc266 (
      {stage0_2[53]},
      {stage1_2[24]}
   );
   gpc1_1 gpc267 (
      {stage0_3[48]},
      {stage1_3[18]}
   );
   gpc1_1 gpc268 (
      {stage0_3[49]},
      {stage1_3[19]}
   );
   gpc1_1 gpc269 (
      {stage0_3[50]},
      {stage1_3[20]}
   );
   gpc1_1 gpc270 (
      {stage0_3[51]},
      {stage1_3[21]}
   );
   gpc1_1 gpc271 (
      {stage0_3[52]},
      {stage1_3[22]}
   );
   gpc1_1 gpc272 (
      {stage0_3[53]},
      {stage1_3[23]}
   );
   gpc1_1 gpc273 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc274 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc275 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc276 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc277 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc278 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc279 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc280 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc281 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc282 (
      {stage0_5[36]},
      {stage1_5[18]}
   );
   gpc1_1 gpc283 (
      {stage0_5[37]},
      {stage1_5[19]}
   );
   gpc1_1 gpc284 (
      {stage0_5[38]},
      {stage1_5[20]}
   );
   gpc1_1 gpc285 (
      {stage0_5[39]},
      {stage1_5[21]}
   );
   gpc1_1 gpc286 (
      {stage0_5[40]},
      {stage1_5[22]}
   );
   gpc1_1 gpc287 (
      {stage0_5[41]},
      {stage1_5[23]}
   );
   gpc1_1 gpc288 (
      {stage0_5[42]},
      {stage1_5[24]}
   );
   gpc1_1 gpc289 (
      {stage0_5[43]},
      {stage1_5[25]}
   );
   gpc1_1 gpc290 (
      {stage0_5[44]},
      {stage1_5[26]}
   );
   gpc1_1 gpc291 (
      {stage0_5[45]},
      {stage1_5[27]}
   );
   gpc1_1 gpc292 (
      {stage0_5[46]},
      {stage1_5[28]}
   );
   gpc1_1 gpc293 (
      {stage0_5[47]},
      {stage1_5[29]}
   );
   gpc1_1 gpc294 (
      {stage0_5[48]},
      {stage1_5[30]}
   );
   gpc1_1 gpc295 (
      {stage0_5[49]},
      {stage1_5[31]}
   );
   gpc1_1 gpc296 (
      {stage0_5[50]},
      {stage1_5[32]}
   );
   gpc1_1 gpc297 (
      {stage0_5[51]},
      {stage1_5[33]}
   );
   gpc1_1 gpc298 (
      {stage0_5[52]},
      {stage1_5[34]}
   );
   gpc1_1 gpc299 (
      {stage0_5[53]},
      {stage1_5[35]}
   );
   gpc1_1 gpc300 (
      {stage0_6[51]},
      {stage1_6[16]}
   );
   gpc1_1 gpc301 (
      {stage0_6[52]},
      {stage1_6[17]}
   );
   gpc1_1 gpc302 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc303 (
      {stage0_7[49]},
      {stage1_7[20]}
   );
   gpc1_1 gpc304 (
      {stage0_7[50]},
      {stage1_7[21]}
   );
   gpc1_1 gpc305 (
      {stage0_7[51]},
      {stage1_7[22]}
   );
   gpc1_1 gpc306 (
      {stage0_7[52]},
      {stage1_7[23]}
   );
   gpc1_1 gpc307 (
      {stage0_7[53]},
      {stage1_7[24]}
   );
   gpc1_1 gpc308 (
      {stage0_8[44]},
      {stage1_8[21]}
   );
   gpc1_1 gpc309 (
      {stage0_8[45]},
      {stage1_8[22]}
   );
   gpc1_1 gpc310 (
      {stage0_8[46]},
      {stage1_8[23]}
   );
   gpc1_1 gpc311 (
      {stage0_8[47]},
      {stage1_8[24]}
   );
   gpc1_1 gpc312 (
      {stage0_8[48]},
      {stage1_8[25]}
   );
   gpc1_1 gpc313 (
      {stage0_8[49]},
      {stage1_8[26]}
   );
   gpc1_1 gpc314 (
      {stage0_8[50]},
      {stage1_8[27]}
   );
   gpc1_1 gpc315 (
      {stage0_8[51]},
      {stage1_8[28]}
   );
   gpc1_1 gpc316 (
      {stage0_8[52]},
      {stage1_8[29]}
   );
   gpc1_1 gpc317 (
      {stage0_8[53]},
      {stage1_8[30]}
   );
   gpc1_1 gpc318 (
      {stage0_10[49]},
      {stage1_10[21]}
   );
   gpc1_1 gpc319 (
      {stage0_10[50]},
      {stage1_10[22]}
   );
   gpc1_1 gpc320 (
      {stage0_10[51]},
      {stage1_10[23]}
   );
   gpc1_1 gpc321 (
      {stage0_10[52]},
      {stage1_10[24]}
   );
   gpc1_1 gpc322 (
      {stage0_10[53]},
      {stage1_10[25]}
   );
   gpc1_1 gpc323 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc324 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc325 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc326 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc327 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc328 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc329 (
      {stage0_12[53]},
      {stage1_12[20]}
   );
   gpc1_1 gpc330 (
      {stage0_13[42]},
      {stage1_13[18]}
   );
   gpc1_1 gpc331 (
      {stage0_13[43]},
      {stage1_13[19]}
   );
   gpc1_1 gpc332 (
      {stage0_13[44]},
      {stage1_13[20]}
   );
   gpc1_1 gpc333 (
      {stage0_13[45]},
      {stage1_13[21]}
   );
   gpc1_1 gpc334 (
      {stage0_13[46]},
      {stage1_13[22]}
   );
   gpc1_1 gpc335 (
      {stage0_13[47]},
      {stage1_13[23]}
   );
   gpc1_1 gpc336 (
      {stage0_13[48]},
      {stage1_13[24]}
   );
   gpc1_1 gpc337 (
      {stage0_13[49]},
      {stage1_13[25]}
   );
   gpc1_1 gpc338 (
      {stage0_13[50]},
      {stage1_13[26]}
   );
   gpc1_1 gpc339 (
      {stage0_13[51]},
      {stage1_13[27]}
   );
   gpc1_1 gpc340 (
      {stage0_13[52]},
      {stage1_13[28]}
   );
   gpc1_1 gpc341 (
      {stage0_13[53]},
      {stage1_13[29]}
   );
   gpc1_1 gpc342 (
      {stage0_14[51]},
      {stage1_14[21]}
   );
   gpc1_1 gpc343 (
      {stage0_14[52]},
      {stage1_14[22]}
   );
   gpc1_1 gpc344 (
      {stage0_14[53]},
      {stage1_14[23]}
   );
   gpc1_1 gpc345 (
      {stage0_15[30]},
      {stage1_15[19]}
   );
   gpc1_1 gpc346 (
      {stage0_15[31]},
      {stage1_15[20]}
   );
   gpc1_1 gpc347 (
      {stage0_15[32]},
      {stage1_15[21]}
   );
   gpc1_1 gpc348 (
      {stage0_15[33]},
      {stage1_15[22]}
   );
   gpc1_1 gpc349 (
      {stage0_15[34]},
      {stage1_15[23]}
   );
   gpc1_1 gpc350 (
      {stage0_15[35]},
      {stage1_15[24]}
   );
   gpc1_1 gpc351 (
      {stage0_15[36]},
      {stage1_15[25]}
   );
   gpc1_1 gpc352 (
      {stage0_15[37]},
      {stage1_15[26]}
   );
   gpc1_1 gpc353 (
      {stage0_15[38]},
      {stage1_15[27]}
   );
   gpc1_1 gpc354 (
      {stage0_15[39]},
      {stage1_15[28]}
   );
   gpc1_1 gpc355 (
      {stage0_15[40]},
      {stage1_15[29]}
   );
   gpc1_1 gpc356 (
      {stage0_15[41]},
      {stage1_15[30]}
   );
   gpc1_1 gpc357 (
      {stage0_15[42]},
      {stage1_15[31]}
   );
   gpc1_1 gpc358 (
      {stage0_15[43]},
      {stage1_15[32]}
   );
   gpc1_1 gpc359 (
      {stage0_15[44]},
      {stage1_15[33]}
   );
   gpc1_1 gpc360 (
      {stage0_15[45]},
      {stage1_15[34]}
   );
   gpc1_1 gpc361 (
      {stage0_15[46]},
      {stage1_15[35]}
   );
   gpc1_1 gpc362 (
      {stage0_15[47]},
      {stage1_15[36]}
   );
   gpc1_1 gpc363 (
      {stage0_15[48]},
      {stage1_15[37]}
   );
   gpc1_1 gpc364 (
      {stage0_15[49]},
      {stage1_15[38]}
   );
   gpc1_1 gpc365 (
      {stage0_15[50]},
      {stage1_15[39]}
   );
   gpc1_1 gpc366 (
      {stage0_15[51]},
      {stage1_15[40]}
   );
   gpc1_1 gpc367 (
      {stage0_15[52]},
      {stage1_15[41]}
   );
   gpc1_1 gpc368 (
      {stage0_15[53]},
      {stage1_15[42]}
   );
   gpc1_1 gpc369 (
      {stage0_16[45]},
      {stage1_16[15]}
   );
   gpc1_1 gpc370 (
      {stage0_16[46]},
      {stage1_16[16]}
   );
   gpc1_1 gpc371 (
      {stage0_16[47]},
      {stage1_16[17]}
   );
   gpc1_1 gpc372 (
      {stage0_16[48]},
      {stage1_16[18]}
   );
   gpc1_1 gpc373 (
      {stage0_16[49]},
      {stage1_16[19]}
   );
   gpc1_1 gpc374 (
      {stage0_16[50]},
      {stage1_16[20]}
   );
   gpc1_1 gpc375 (
      {stage0_16[51]},
      {stage1_16[21]}
   );
   gpc1_1 gpc376 (
      {stage0_16[52]},
      {stage1_16[22]}
   );
   gpc1_1 gpc377 (
      {stage0_16[53]},
      {stage1_16[23]}
   );
   gpc1_1 gpc378 (
      {stage0_18[42]},
      {stage1_18[22]}
   );
   gpc1_1 gpc379 (
      {stage0_18[43]},
      {stage1_18[23]}
   );
   gpc1_1 gpc380 (
      {stage0_18[44]},
      {stage1_18[24]}
   );
   gpc1_1 gpc381 (
      {stage0_18[45]},
      {stage1_18[25]}
   );
   gpc1_1 gpc382 (
      {stage0_18[46]},
      {stage1_18[26]}
   );
   gpc1_1 gpc383 (
      {stage0_18[47]},
      {stage1_18[27]}
   );
   gpc1_1 gpc384 (
      {stage0_18[48]},
      {stage1_18[28]}
   );
   gpc1_1 gpc385 (
      {stage0_18[49]},
      {stage1_18[29]}
   );
   gpc1_1 gpc386 (
      {stage0_18[50]},
      {stage1_18[30]}
   );
   gpc1_1 gpc387 (
      {stage0_18[51]},
      {stage1_18[31]}
   );
   gpc1_1 gpc388 (
      {stage0_18[52]},
      {stage1_18[32]}
   );
   gpc1_1 gpc389 (
      {stage0_18[53]},
      {stage1_18[33]}
   );
   gpc1_1 gpc390 (
      {stage0_19[52]},
      {stage1_19[19]}
   );
   gpc1_1 gpc391 (
      {stage0_19[53]},
      {stage1_19[20]}
   );
   gpc1_1 gpc392 (
      {stage0_20[53]},
      {stage1_20[19]}
   );
   gpc1_1 gpc393 (
      {stage0_21[51]},
      {stage1_21[23]}
   );
   gpc1_1 gpc394 (
      {stage0_21[52]},
      {stage1_21[24]}
   );
   gpc1_1 gpc395 (
      {stage0_21[53]},
      {stage1_21[25]}
   );
   gpc1_1 gpc396 (
      {stage0_24[41]},
      {stage1_24[19]}
   );
   gpc1_1 gpc397 (
      {stage0_24[42]},
      {stage1_24[20]}
   );
   gpc1_1 gpc398 (
      {stage0_24[43]},
      {stage1_24[21]}
   );
   gpc1_1 gpc399 (
      {stage0_24[44]},
      {stage1_24[22]}
   );
   gpc1_1 gpc400 (
      {stage0_24[45]},
      {stage1_24[23]}
   );
   gpc1_1 gpc401 (
      {stage0_24[46]},
      {stage1_24[24]}
   );
   gpc1_1 gpc402 (
      {stage0_24[47]},
      {stage1_24[25]}
   );
   gpc1_1 gpc403 (
      {stage0_24[48]},
      {stage1_24[26]}
   );
   gpc1_1 gpc404 (
      {stage0_24[49]},
      {stage1_24[27]}
   );
   gpc1_1 gpc405 (
      {stage0_24[50]},
      {stage1_24[28]}
   );
   gpc1_1 gpc406 (
      {stage0_24[51]},
      {stage1_24[29]}
   );
   gpc1_1 gpc407 (
      {stage0_24[52]},
      {stage1_24[30]}
   );
   gpc1_1 gpc408 (
      {stage0_24[53]},
      {stage1_24[31]}
   );
   gpc1_1 gpc409 (
      {stage0_25[48]},
      {stage1_25[19]}
   );
   gpc1_1 gpc410 (
      {stage0_25[49]},
      {stage1_25[20]}
   );
   gpc1_1 gpc411 (
      {stage0_25[50]},
      {stage1_25[21]}
   );
   gpc1_1 gpc412 (
      {stage0_25[51]},
      {stage1_25[22]}
   );
   gpc1_1 gpc413 (
      {stage0_25[52]},
      {stage1_25[23]}
   );
   gpc1_1 gpc414 (
      {stage0_25[53]},
      {stage1_25[24]}
   );
   gpc1_1 gpc415 (
      {stage0_26[45]},
      {stage1_26[23]}
   );
   gpc1_1 gpc416 (
      {stage0_26[46]},
      {stage1_26[24]}
   );
   gpc1_1 gpc417 (
      {stage0_26[47]},
      {stage1_26[25]}
   );
   gpc1_1 gpc418 (
      {stage0_26[48]},
      {stage1_26[26]}
   );
   gpc1_1 gpc419 (
      {stage0_26[49]},
      {stage1_26[27]}
   );
   gpc1_1 gpc420 (
      {stage0_26[50]},
      {stage1_26[28]}
   );
   gpc1_1 gpc421 (
      {stage0_26[51]},
      {stage1_26[29]}
   );
   gpc1_1 gpc422 (
      {stage0_26[52]},
      {stage1_26[30]}
   );
   gpc1_1 gpc423 (
      {stage0_26[53]},
      {stage1_26[31]}
   );
   gpc1_1 gpc424 (
      {stage0_27[50]},
      {stage1_27[20]}
   );
   gpc1_1 gpc425 (
      {stage0_27[51]},
      {stage1_27[21]}
   );
   gpc1_1 gpc426 (
      {stage0_27[52]},
      {stage1_27[22]}
   );
   gpc1_1 gpc427 (
      {stage0_27[53]},
      {stage1_27[23]}
   );
   gpc1_1 gpc428 (
      {stage0_29[50]},
      {stage1_29[22]}
   );
   gpc1_1 gpc429 (
      {stage0_29[51]},
      {stage1_29[23]}
   );
   gpc1_1 gpc430 (
      {stage0_29[52]},
      {stage1_29[24]}
   );
   gpc1_1 gpc431 (
      {stage0_29[53]},
      {stage1_29[25]}
   );
   gpc1_1 gpc432 (
      {stage0_30[42]},
      {stage1_30[23]}
   );
   gpc1_1 gpc433 (
      {stage0_30[43]},
      {stage1_30[24]}
   );
   gpc1_1 gpc434 (
      {stage0_30[44]},
      {stage1_30[25]}
   );
   gpc1_1 gpc435 (
      {stage0_30[45]},
      {stage1_30[26]}
   );
   gpc1_1 gpc436 (
      {stage0_30[46]},
      {stage1_30[27]}
   );
   gpc1_1 gpc437 (
      {stage0_30[47]},
      {stage1_30[28]}
   );
   gpc1_1 gpc438 (
      {stage0_30[48]},
      {stage1_30[29]}
   );
   gpc1_1 gpc439 (
      {stage0_30[49]},
      {stage1_30[30]}
   );
   gpc1_1 gpc440 (
      {stage0_30[50]},
      {stage1_30[31]}
   );
   gpc1_1 gpc441 (
      {stage0_30[51]},
      {stage1_30[32]}
   );
   gpc1_1 gpc442 (
      {stage0_30[52]},
      {stage1_30[33]}
   );
   gpc1_1 gpc443 (
      {stage0_30[53]},
      {stage1_30[34]}
   );
   gpc1_1 gpc444 (
      {stage0_31[36]},
      {stage1_31[16]}
   );
   gpc1_1 gpc445 (
      {stage0_31[37]},
      {stage1_31[17]}
   );
   gpc1_1 gpc446 (
      {stage0_31[38]},
      {stage1_31[18]}
   );
   gpc1_1 gpc447 (
      {stage0_31[39]},
      {stage1_31[19]}
   );
   gpc1_1 gpc448 (
      {stage0_31[40]},
      {stage1_31[20]}
   );
   gpc1_1 gpc449 (
      {stage0_31[41]},
      {stage1_31[21]}
   );
   gpc1_1 gpc450 (
      {stage0_31[42]},
      {stage1_31[22]}
   );
   gpc1_1 gpc451 (
      {stage0_31[43]},
      {stage1_31[23]}
   );
   gpc1_1 gpc452 (
      {stage0_31[44]},
      {stage1_31[24]}
   );
   gpc1_1 gpc453 (
      {stage0_31[45]},
      {stage1_31[25]}
   );
   gpc1_1 gpc454 (
      {stage0_31[46]},
      {stage1_31[26]}
   );
   gpc1_1 gpc455 (
      {stage0_31[47]},
      {stage1_31[27]}
   );
   gpc1_1 gpc456 (
      {stage0_31[48]},
      {stage1_31[28]}
   );
   gpc1_1 gpc457 (
      {stage0_31[49]},
      {stage1_31[29]}
   );
   gpc1_1 gpc458 (
      {stage0_31[50]},
      {stage1_31[30]}
   );
   gpc1_1 gpc459 (
      {stage0_31[51]},
      {stage1_31[31]}
   );
   gpc1_1 gpc460 (
      {stage0_31[52]},
      {stage1_31[32]}
   );
   gpc1_1 gpc461 (
      {stage0_31[53]},
      {stage1_31[33]}
   );
   gpc1_1 gpc462 (
      {stage0_32[53]},
      {stage1_32[18]}
   );
   gpc1_1 gpc463 (
      {stage0_33[25]},
      {stage1_33[17]}
   );
   gpc1_1 gpc464 (
      {stage0_33[26]},
      {stage1_33[18]}
   );
   gpc1_1 gpc465 (
      {stage0_33[27]},
      {stage1_33[19]}
   );
   gpc1_1 gpc466 (
      {stage0_33[28]},
      {stage1_33[20]}
   );
   gpc1_1 gpc467 (
      {stage0_33[29]},
      {stage1_33[21]}
   );
   gpc1_1 gpc468 (
      {stage0_33[30]},
      {stage1_33[22]}
   );
   gpc1_1 gpc469 (
      {stage0_33[31]},
      {stage1_33[23]}
   );
   gpc1_1 gpc470 (
      {stage0_33[32]},
      {stage1_33[24]}
   );
   gpc1_1 gpc471 (
      {stage0_33[33]},
      {stage1_33[25]}
   );
   gpc1_1 gpc472 (
      {stage0_33[34]},
      {stage1_33[26]}
   );
   gpc1_1 gpc473 (
      {stage0_33[35]},
      {stage1_33[27]}
   );
   gpc1_1 gpc474 (
      {stage0_33[36]},
      {stage1_33[28]}
   );
   gpc1_1 gpc475 (
      {stage0_33[37]},
      {stage1_33[29]}
   );
   gpc1_1 gpc476 (
      {stage0_33[38]},
      {stage1_33[30]}
   );
   gpc1_1 gpc477 (
      {stage0_33[39]},
      {stage1_33[31]}
   );
   gpc1_1 gpc478 (
      {stage0_33[40]},
      {stage1_33[32]}
   );
   gpc1_1 gpc479 (
      {stage0_33[41]},
      {stage1_33[33]}
   );
   gpc1_1 gpc480 (
      {stage0_33[42]},
      {stage1_33[34]}
   );
   gpc1_1 gpc481 (
      {stage0_33[43]},
      {stage1_33[35]}
   );
   gpc1_1 gpc482 (
      {stage0_33[44]},
      {stage1_33[36]}
   );
   gpc1_1 gpc483 (
      {stage0_33[45]},
      {stage1_33[37]}
   );
   gpc1_1 gpc484 (
      {stage0_33[46]},
      {stage1_33[38]}
   );
   gpc1_1 gpc485 (
      {stage0_33[47]},
      {stage1_33[39]}
   );
   gpc1_1 gpc486 (
      {stage0_33[48]},
      {stage1_33[40]}
   );
   gpc1_1 gpc487 (
      {stage0_33[49]},
      {stage1_33[41]}
   );
   gpc1_1 gpc488 (
      {stage0_33[50]},
      {stage1_33[42]}
   );
   gpc1_1 gpc489 (
      {stage0_33[51]},
      {stage1_33[43]}
   );
   gpc1_1 gpc490 (
      {stage0_33[52]},
      {stage1_33[44]}
   );
   gpc1_1 gpc491 (
      {stage0_33[53]},
      {stage1_33[45]}
   );
   gpc1_1 gpc492 (
      {stage0_34[51]},
      {stage1_34[16]}
   );
   gpc1_1 gpc493 (
      {stage0_34[52]},
      {stage1_34[17]}
   );
   gpc1_1 gpc494 (
      {stage0_34[53]},
      {stage1_34[18]}
   );
   gpc1_1 gpc495 (
      {stage0_35[43]},
      {stage1_35[17]}
   );
   gpc1_1 gpc496 (
      {stage0_35[44]},
      {stage1_35[18]}
   );
   gpc1_1 gpc497 (
      {stage0_35[45]},
      {stage1_35[19]}
   );
   gpc1_1 gpc498 (
      {stage0_35[46]},
      {stage1_35[20]}
   );
   gpc1_1 gpc499 (
      {stage0_35[47]},
      {stage1_35[21]}
   );
   gpc1_1 gpc500 (
      {stage0_35[48]},
      {stage1_35[22]}
   );
   gpc1_1 gpc501 (
      {stage0_35[49]},
      {stage1_35[23]}
   );
   gpc1_1 gpc502 (
      {stage0_35[50]},
      {stage1_35[24]}
   );
   gpc1_1 gpc503 (
      {stage0_35[51]},
      {stage1_35[25]}
   );
   gpc1_1 gpc504 (
      {stage0_35[52]},
      {stage1_35[26]}
   );
   gpc1_1 gpc505 (
      {stage0_35[53]},
      {stage1_35[27]}
   );
   gpc1_1 gpc506 (
      {stage0_36[41]},
      {stage1_36[21]}
   );
   gpc1_1 gpc507 (
      {stage0_36[42]},
      {stage1_36[22]}
   );
   gpc1_1 gpc508 (
      {stage0_36[43]},
      {stage1_36[23]}
   );
   gpc1_1 gpc509 (
      {stage0_36[44]},
      {stage1_36[24]}
   );
   gpc1_1 gpc510 (
      {stage0_36[45]},
      {stage1_36[25]}
   );
   gpc1_1 gpc511 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc512 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc513 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc514 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc515 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc516 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc517 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc518 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc519 (
      {stage0_37[48]},
      {stage1_37[19]}
   );
   gpc1_1 gpc520 (
      {stage0_37[49]},
      {stage1_37[20]}
   );
   gpc1_1 gpc521 (
      {stage0_37[50]},
      {stage1_37[21]}
   );
   gpc1_1 gpc522 (
      {stage0_37[51]},
      {stage1_37[22]}
   );
   gpc1_1 gpc523 (
      {stage0_37[52]},
      {stage1_37[23]}
   );
   gpc1_1 gpc524 (
      {stage0_37[53]},
      {stage1_37[24]}
   );
   gpc1_1 gpc525 (
      {stage0_38[46]},
      {stage1_38[16]}
   );
   gpc1_1 gpc526 (
      {stage0_38[47]},
      {stage1_38[17]}
   );
   gpc1_1 gpc527 (
      {stage0_38[48]},
      {stage1_38[18]}
   );
   gpc1_1 gpc528 (
      {stage0_38[49]},
      {stage1_38[19]}
   );
   gpc1_1 gpc529 (
      {stage0_38[50]},
      {stage1_38[20]}
   );
   gpc1_1 gpc530 (
      {stage0_38[51]},
      {stage1_38[21]}
   );
   gpc1_1 gpc531 (
      {stage0_38[52]},
      {stage1_38[22]}
   );
   gpc1_1 gpc532 (
      {stage0_38[53]},
      {stage1_38[23]}
   );
   gpc1_1 gpc533 (
      {stage0_39[43]},
      {stage1_39[20]}
   );
   gpc1_1 gpc534 (
      {stage0_39[44]},
      {stage1_39[21]}
   );
   gpc1_1 gpc535 (
      {stage0_39[45]},
      {stage1_39[22]}
   );
   gpc1_1 gpc536 (
      {stage0_39[46]},
      {stage1_39[23]}
   );
   gpc1_1 gpc537 (
      {stage0_39[47]},
      {stage1_39[24]}
   );
   gpc1_1 gpc538 (
      {stage0_39[48]},
      {stage1_39[25]}
   );
   gpc1_1 gpc539 (
      {stage0_39[49]},
      {stage1_39[26]}
   );
   gpc1_1 gpc540 (
      {stage0_39[50]},
      {stage1_39[27]}
   );
   gpc1_1 gpc541 (
      {stage0_39[51]},
      {stage1_39[28]}
   );
   gpc1_1 gpc542 (
      {stage0_39[52]},
      {stage1_39[29]}
   );
   gpc1_1 gpc543 (
      {stage0_39[53]},
      {stage1_39[30]}
   );
   gpc1_1 gpc544 (
      {stage0_40[34]},
      {stage1_40[19]}
   );
   gpc1_1 gpc545 (
      {stage0_40[35]},
      {stage1_40[20]}
   );
   gpc1_1 gpc546 (
      {stage0_40[36]},
      {stage1_40[21]}
   );
   gpc1_1 gpc547 (
      {stage0_40[37]},
      {stage1_40[22]}
   );
   gpc1_1 gpc548 (
      {stage0_40[38]},
      {stage1_40[23]}
   );
   gpc1_1 gpc549 (
      {stage0_40[39]},
      {stage1_40[24]}
   );
   gpc1_1 gpc550 (
      {stage0_40[40]},
      {stage1_40[25]}
   );
   gpc1_1 gpc551 (
      {stage0_40[41]},
      {stage1_40[26]}
   );
   gpc1_1 gpc552 (
      {stage0_40[42]},
      {stage1_40[27]}
   );
   gpc1_1 gpc553 (
      {stage0_40[43]},
      {stage1_40[28]}
   );
   gpc1_1 gpc554 (
      {stage0_40[44]},
      {stage1_40[29]}
   );
   gpc1_1 gpc555 (
      {stage0_40[45]},
      {stage1_40[30]}
   );
   gpc1_1 gpc556 (
      {stage0_40[46]},
      {stage1_40[31]}
   );
   gpc1_1 gpc557 (
      {stage0_40[47]},
      {stage1_40[32]}
   );
   gpc1_1 gpc558 (
      {stage0_40[48]},
      {stage1_40[33]}
   );
   gpc1_1 gpc559 (
      {stage0_40[49]},
      {stage1_40[34]}
   );
   gpc1_1 gpc560 (
      {stage0_40[50]},
      {stage1_40[35]}
   );
   gpc1_1 gpc561 (
      {stage0_40[51]},
      {stage1_40[36]}
   );
   gpc1_1 gpc562 (
      {stage0_40[52]},
      {stage1_40[37]}
   );
   gpc1_1 gpc563 (
      {stage0_40[53]},
      {stage1_40[38]}
   );
   gpc1_1 gpc564 (
      {stage0_41[51]},
      {stage1_41[17]}
   );
   gpc1_1 gpc565 (
      {stage0_41[52]},
      {stage1_41[18]}
   );
   gpc1_1 gpc566 (
      {stage0_41[53]},
      {stage1_41[19]}
   );
   gpc1_1 gpc567 (
      {stage0_42[52]},
      {stage1_42[19]}
   );
   gpc1_1 gpc568 (
      {stage0_42[53]},
      {stage1_42[20]}
   );
   gpc1_1 gpc569 (
      {stage0_45[41]},
      {stage1_45[19]}
   );
   gpc1_1 gpc570 (
      {stage0_45[42]},
      {stage1_45[20]}
   );
   gpc1_1 gpc571 (
      {stage0_45[43]},
      {stage1_45[21]}
   );
   gpc1_1 gpc572 (
      {stage0_45[44]},
      {stage1_45[22]}
   );
   gpc1_1 gpc573 (
      {stage0_45[45]},
      {stage1_45[23]}
   );
   gpc1_1 gpc574 (
      {stage0_45[46]},
      {stage1_45[24]}
   );
   gpc1_1 gpc575 (
      {stage0_45[47]},
      {stage1_45[25]}
   );
   gpc1_1 gpc576 (
      {stage0_45[48]},
      {stage1_45[26]}
   );
   gpc1_1 gpc577 (
      {stage0_45[49]},
      {stage1_45[27]}
   );
   gpc1_1 gpc578 (
      {stage0_45[50]},
      {stage1_45[28]}
   );
   gpc1_1 gpc579 (
      {stage0_45[51]},
      {stage1_45[29]}
   );
   gpc1_1 gpc580 (
      {stage0_45[52]},
      {stage1_45[30]}
   );
   gpc1_1 gpc581 (
      {stage0_45[53]},
      {stage1_45[31]}
   );
   gpc1_1 gpc582 (
      {stage0_46[44]},
      {stage1_46[20]}
   );
   gpc1_1 gpc583 (
      {stage0_46[45]},
      {stage1_46[21]}
   );
   gpc1_1 gpc584 (
      {stage0_46[46]},
      {stage1_46[22]}
   );
   gpc1_1 gpc585 (
      {stage0_46[47]},
      {stage1_46[23]}
   );
   gpc1_1 gpc586 (
      {stage0_46[48]},
      {stage1_46[24]}
   );
   gpc1_1 gpc587 (
      {stage0_46[49]},
      {stage1_46[25]}
   );
   gpc1_1 gpc588 (
      {stage0_46[50]},
      {stage1_46[26]}
   );
   gpc1_1 gpc589 (
      {stage0_46[51]},
      {stage1_46[27]}
   );
   gpc1_1 gpc590 (
      {stage0_46[52]},
      {stage1_46[28]}
   );
   gpc1_1 gpc591 (
      {stage0_46[53]},
      {stage1_46[29]}
   );
   gpc1_1 gpc592 (
      {stage0_47[41]},
      {stage1_47[21]}
   );
   gpc1_1 gpc593 (
      {stage0_47[42]},
      {stage1_47[22]}
   );
   gpc1_1 gpc594 (
      {stage0_47[43]},
      {stage1_47[23]}
   );
   gpc1_1 gpc595 (
      {stage0_47[44]},
      {stage1_47[24]}
   );
   gpc1_1 gpc596 (
      {stage0_47[45]},
      {stage1_47[25]}
   );
   gpc1_1 gpc597 (
      {stage0_47[46]},
      {stage1_47[26]}
   );
   gpc1_1 gpc598 (
      {stage0_47[47]},
      {stage1_47[27]}
   );
   gpc1_1 gpc599 (
      {stage0_47[48]},
      {stage1_47[28]}
   );
   gpc1_1 gpc600 (
      {stage0_47[49]},
      {stage1_47[29]}
   );
   gpc1_1 gpc601 (
      {stage0_47[50]},
      {stage1_47[30]}
   );
   gpc1_1 gpc602 (
      {stage0_47[51]},
      {stage1_47[31]}
   );
   gpc1_1 gpc603 (
      {stage0_47[52]},
      {stage1_47[32]}
   );
   gpc1_1 gpc604 (
      {stage0_47[53]},
      {stage1_47[33]}
   );
   gpc1_1 gpc605 (
      {stage0_49[47]},
      {stage1_49[17]}
   );
   gpc1_1 gpc606 (
      {stage0_49[48]},
      {stage1_49[18]}
   );
   gpc1_1 gpc607 (
      {stage0_49[49]},
      {stage1_49[19]}
   );
   gpc1_1 gpc608 (
      {stage0_49[50]},
      {stage1_49[20]}
   );
   gpc1_1 gpc609 (
      {stage0_49[51]},
      {stage1_49[21]}
   );
   gpc1_1 gpc610 (
      {stage0_49[52]},
      {stage1_49[22]}
   );
   gpc1_1 gpc611 (
      {stage0_49[53]},
      {stage1_49[23]}
   );
   gpc1_1 gpc612 (
      {stage0_50[29]},
      {stage1_50[18]}
   );
   gpc1_1 gpc613 (
      {stage0_50[30]},
      {stage1_50[19]}
   );
   gpc1_1 gpc614 (
      {stage0_50[31]},
      {stage1_50[20]}
   );
   gpc1_1 gpc615 (
      {stage0_50[32]},
      {stage1_50[21]}
   );
   gpc1_1 gpc616 (
      {stage0_50[33]},
      {stage1_50[22]}
   );
   gpc1_1 gpc617 (
      {stage0_50[34]},
      {stage1_50[23]}
   );
   gpc1_1 gpc618 (
      {stage0_50[35]},
      {stage1_50[24]}
   );
   gpc1_1 gpc619 (
      {stage0_50[36]},
      {stage1_50[25]}
   );
   gpc1_1 gpc620 (
      {stage0_50[37]},
      {stage1_50[26]}
   );
   gpc1_1 gpc621 (
      {stage0_50[38]},
      {stage1_50[27]}
   );
   gpc1_1 gpc622 (
      {stage0_50[39]},
      {stage1_50[28]}
   );
   gpc1_1 gpc623 (
      {stage0_50[40]},
      {stage1_50[29]}
   );
   gpc1_1 gpc624 (
      {stage0_50[41]},
      {stage1_50[30]}
   );
   gpc1_1 gpc625 (
      {stage0_50[42]},
      {stage1_50[31]}
   );
   gpc1_1 gpc626 (
      {stage0_50[43]},
      {stage1_50[32]}
   );
   gpc1_1 gpc627 (
      {stage0_50[44]},
      {stage1_50[33]}
   );
   gpc1_1 gpc628 (
      {stage0_50[45]},
      {stage1_50[34]}
   );
   gpc1_1 gpc629 (
      {stage0_50[46]},
      {stage1_50[35]}
   );
   gpc1_1 gpc630 (
      {stage0_50[47]},
      {stage1_50[36]}
   );
   gpc1_1 gpc631 (
      {stage0_50[48]},
      {stage1_50[37]}
   );
   gpc1_1 gpc632 (
      {stage0_50[49]},
      {stage1_50[38]}
   );
   gpc1_1 gpc633 (
      {stage0_50[50]},
      {stage1_50[39]}
   );
   gpc1_1 gpc634 (
      {stage0_50[51]},
      {stage1_50[40]}
   );
   gpc1_1 gpc635 (
      {stage0_50[52]},
      {stage1_50[41]}
   );
   gpc1_1 gpc636 (
      {stage0_50[53]},
      {stage1_50[42]}
   );
   gpc1_1 gpc637 (
      {stage0_51[20]},
      {stage1_51[14]}
   );
   gpc1_1 gpc638 (
      {stage0_51[21]},
      {stage1_51[15]}
   );
   gpc1_1 gpc639 (
      {stage0_51[22]},
      {stage1_51[16]}
   );
   gpc1_1 gpc640 (
      {stage0_51[23]},
      {stage1_51[17]}
   );
   gpc1_1 gpc641 (
      {stage0_51[24]},
      {stage1_51[18]}
   );
   gpc1_1 gpc642 (
      {stage0_51[25]},
      {stage1_51[19]}
   );
   gpc1_1 gpc643 (
      {stage0_51[26]},
      {stage1_51[20]}
   );
   gpc1_1 gpc644 (
      {stage0_51[27]},
      {stage1_51[21]}
   );
   gpc1_1 gpc645 (
      {stage0_51[28]},
      {stage1_51[22]}
   );
   gpc1_1 gpc646 (
      {stage0_51[29]},
      {stage1_51[23]}
   );
   gpc1_1 gpc647 (
      {stage0_51[30]},
      {stage1_51[24]}
   );
   gpc1_1 gpc648 (
      {stage0_51[31]},
      {stage1_51[25]}
   );
   gpc1_1 gpc649 (
      {stage0_51[32]},
      {stage1_51[26]}
   );
   gpc1_1 gpc650 (
      {stage0_51[33]},
      {stage1_51[27]}
   );
   gpc1_1 gpc651 (
      {stage0_51[34]},
      {stage1_51[28]}
   );
   gpc1_1 gpc652 (
      {stage0_51[35]},
      {stage1_51[29]}
   );
   gpc1_1 gpc653 (
      {stage0_51[36]},
      {stage1_51[30]}
   );
   gpc1_1 gpc654 (
      {stage0_51[37]},
      {stage1_51[31]}
   );
   gpc1_1 gpc655 (
      {stage0_51[38]},
      {stage1_51[32]}
   );
   gpc1_1 gpc656 (
      {stage0_51[39]},
      {stage1_51[33]}
   );
   gpc1_1 gpc657 (
      {stage0_51[40]},
      {stage1_51[34]}
   );
   gpc1_1 gpc658 (
      {stage0_51[41]},
      {stage1_51[35]}
   );
   gpc1_1 gpc659 (
      {stage0_51[42]},
      {stage1_51[36]}
   );
   gpc1_1 gpc660 (
      {stage0_51[43]},
      {stage1_51[37]}
   );
   gpc1_1 gpc661 (
      {stage0_51[44]},
      {stage1_51[38]}
   );
   gpc1_1 gpc662 (
      {stage0_51[45]},
      {stage1_51[39]}
   );
   gpc1_1 gpc663 (
      {stage0_51[46]},
      {stage1_51[40]}
   );
   gpc1_1 gpc664 (
      {stage0_51[47]},
      {stage1_51[41]}
   );
   gpc1_1 gpc665 (
      {stage0_51[48]},
      {stage1_51[42]}
   );
   gpc1_1 gpc666 (
      {stage0_51[49]},
      {stage1_51[43]}
   );
   gpc1_1 gpc667 (
      {stage0_51[50]},
      {stage1_51[44]}
   );
   gpc1_1 gpc668 (
      {stage0_51[51]},
      {stage1_51[45]}
   );
   gpc1_1 gpc669 (
      {stage0_51[52]},
      {stage1_51[46]}
   );
   gpc1_1 gpc670 (
      {stage0_51[53]},
      {stage1_51[47]}
   );
   gpc1_1 gpc671 (
      {stage0_52[47]},
      {stage1_52[15]}
   );
   gpc1_1 gpc672 (
      {stage0_52[48]},
      {stage1_52[16]}
   );
   gpc1_1 gpc673 (
      {stage0_52[49]},
      {stage1_52[17]}
   );
   gpc1_1 gpc674 (
      {stage0_52[50]},
      {stage1_52[18]}
   );
   gpc1_1 gpc675 (
      {stage0_52[51]},
      {stage1_52[19]}
   );
   gpc1_1 gpc676 (
      {stage0_52[52]},
      {stage1_52[20]}
   );
   gpc1_1 gpc677 (
      {stage0_52[53]},
      {stage1_52[21]}
   );
   gpc1_1 gpc678 (
      {stage0_53[28]},
      {stage1_53[15]}
   );
   gpc1_1 gpc679 (
      {stage0_53[29]},
      {stage1_53[16]}
   );
   gpc1_1 gpc680 (
      {stage0_53[30]},
      {stage1_53[17]}
   );
   gpc1_1 gpc681 (
      {stage0_53[31]},
      {stage1_53[18]}
   );
   gpc1_1 gpc682 (
      {stage0_53[32]},
      {stage1_53[19]}
   );
   gpc1_1 gpc683 (
      {stage0_53[33]},
      {stage1_53[20]}
   );
   gpc1_1 gpc684 (
      {stage0_53[34]},
      {stage1_53[21]}
   );
   gpc1_1 gpc685 (
      {stage0_53[35]},
      {stage1_53[22]}
   );
   gpc1_1 gpc686 (
      {stage0_53[36]},
      {stage1_53[23]}
   );
   gpc1_1 gpc687 (
      {stage0_53[37]},
      {stage1_53[24]}
   );
   gpc1_1 gpc688 (
      {stage0_53[38]},
      {stage1_53[25]}
   );
   gpc1_1 gpc689 (
      {stage0_53[39]},
      {stage1_53[26]}
   );
   gpc1_1 gpc690 (
      {stage0_53[40]},
      {stage1_53[27]}
   );
   gpc1_1 gpc691 (
      {stage0_53[41]},
      {stage1_53[28]}
   );
   gpc1_1 gpc692 (
      {stage0_53[42]},
      {stage1_53[29]}
   );
   gpc1_1 gpc693 (
      {stage0_53[43]},
      {stage1_53[30]}
   );
   gpc1_1 gpc694 (
      {stage0_53[44]},
      {stage1_53[31]}
   );
   gpc1_1 gpc695 (
      {stage0_53[45]},
      {stage1_53[32]}
   );
   gpc1_1 gpc696 (
      {stage0_53[46]},
      {stage1_53[33]}
   );
   gpc1_1 gpc697 (
      {stage0_53[47]},
      {stage1_53[34]}
   );
   gpc1_1 gpc698 (
      {stage0_53[48]},
      {stage1_53[35]}
   );
   gpc1_1 gpc699 (
      {stage0_53[49]},
      {stage1_53[36]}
   );
   gpc1_1 gpc700 (
      {stage0_53[50]},
      {stage1_53[37]}
   );
   gpc1_1 gpc701 (
      {stage0_53[51]},
      {stage1_53[38]}
   );
   gpc1_1 gpc702 (
      {stage0_53[52]},
      {stage1_53[39]}
   );
   gpc1_1 gpc703 (
      {stage0_53[53]},
      {stage1_53[40]}
   );
   gpc1_1 gpc704 (
      {stage0_54[51]},
      {stage1_54[14]}
   );
   gpc1_1 gpc705 (
      {stage0_54[52]},
      {stage1_54[15]}
   );
   gpc1_1 gpc706 (
      {stage0_54[53]},
      {stage1_54[16]}
   );
   gpc1_1 gpc707 (
      {stage0_55[30]},
      {stage1_55[14]}
   );
   gpc1_1 gpc708 (
      {stage0_55[31]},
      {stage1_55[15]}
   );
   gpc1_1 gpc709 (
      {stage0_55[32]},
      {stage1_55[16]}
   );
   gpc1_1 gpc710 (
      {stage0_55[33]},
      {stage1_55[17]}
   );
   gpc1_1 gpc711 (
      {stage0_55[34]},
      {stage1_55[18]}
   );
   gpc1_1 gpc712 (
      {stage0_55[35]},
      {stage1_55[19]}
   );
   gpc1_1 gpc713 (
      {stage0_55[36]},
      {stage1_55[20]}
   );
   gpc1_1 gpc714 (
      {stage0_55[37]},
      {stage1_55[21]}
   );
   gpc1_1 gpc715 (
      {stage0_55[38]},
      {stage1_55[22]}
   );
   gpc1_1 gpc716 (
      {stage0_55[39]},
      {stage1_55[23]}
   );
   gpc1_1 gpc717 (
      {stage0_55[40]},
      {stage1_55[24]}
   );
   gpc1_1 gpc718 (
      {stage0_55[41]},
      {stage1_55[25]}
   );
   gpc1_1 gpc719 (
      {stage0_55[42]},
      {stage1_55[26]}
   );
   gpc1_1 gpc720 (
      {stage0_55[43]},
      {stage1_55[27]}
   );
   gpc1_1 gpc721 (
      {stage0_55[44]},
      {stage1_55[28]}
   );
   gpc1_1 gpc722 (
      {stage0_55[45]},
      {stage1_55[29]}
   );
   gpc1_1 gpc723 (
      {stage0_55[46]},
      {stage1_55[30]}
   );
   gpc1_1 gpc724 (
      {stage0_55[47]},
      {stage1_55[31]}
   );
   gpc1_1 gpc725 (
      {stage0_55[48]},
      {stage1_55[32]}
   );
   gpc1_1 gpc726 (
      {stage0_55[49]},
      {stage1_55[33]}
   );
   gpc1_1 gpc727 (
      {stage0_55[50]},
      {stage1_55[34]}
   );
   gpc1_1 gpc728 (
      {stage0_55[51]},
      {stage1_55[35]}
   );
   gpc1_1 gpc729 (
      {stage0_55[52]},
      {stage1_55[36]}
   );
   gpc1_1 gpc730 (
      {stage0_55[53]},
      {stage1_55[37]}
   );
   gpc1_1 gpc731 (
      {stage0_57[30]},
      {stage1_57[17]}
   );
   gpc1_1 gpc732 (
      {stage0_57[31]},
      {stage1_57[18]}
   );
   gpc1_1 gpc733 (
      {stage0_57[32]},
      {stage1_57[19]}
   );
   gpc1_1 gpc734 (
      {stage0_57[33]},
      {stage1_57[20]}
   );
   gpc1_1 gpc735 (
      {stage0_57[34]},
      {stage1_57[21]}
   );
   gpc1_1 gpc736 (
      {stage0_57[35]},
      {stage1_57[22]}
   );
   gpc1_1 gpc737 (
      {stage0_57[36]},
      {stage1_57[23]}
   );
   gpc1_1 gpc738 (
      {stage0_57[37]},
      {stage1_57[24]}
   );
   gpc1_1 gpc739 (
      {stage0_57[38]},
      {stage1_57[25]}
   );
   gpc1_1 gpc740 (
      {stage0_57[39]},
      {stage1_57[26]}
   );
   gpc1_1 gpc741 (
      {stage0_57[40]},
      {stage1_57[27]}
   );
   gpc1_1 gpc742 (
      {stage0_57[41]},
      {stage1_57[28]}
   );
   gpc1_1 gpc743 (
      {stage0_57[42]},
      {stage1_57[29]}
   );
   gpc1_1 gpc744 (
      {stage0_57[43]},
      {stage1_57[30]}
   );
   gpc1_1 gpc745 (
      {stage0_57[44]},
      {stage1_57[31]}
   );
   gpc1_1 gpc746 (
      {stage0_57[45]},
      {stage1_57[32]}
   );
   gpc1_1 gpc747 (
      {stage0_57[46]},
      {stage1_57[33]}
   );
   gpc1_1 gpc748 (
      {stage0_57[47]},
      {stage1_57[34]}
   );
   gpc1_1 gpc749 (
      {stage0_57[48]},
      {stage1_57[35]}
   );
   gpc1_1 gpc750 (
      {stage0_57[49]},
      {stage1_57[36]}
   );
   gpc1_1 gpc751 (
      {stage0_57[50]},
      {stage1_57[37]}
   );
   gpc1_1 gpc752 (
      {stage0_57[51]},
      {stage1_57[38]}
   );
   gpc1_1 gpc753 (
      {stage0_57[52]},
      {stage1_57[39]}
   );
   gpc1_1 gpc754 (
      {stage0_57[53]},
      {stage1_57[40]}
   );
   gpc1_1 gpc755 (
      {stage0_59[36]},
      {stage1_59[17]}
   );
   gpc1_1 gpc756 (
      {stage0_59[37]},
      {stage1_59[18]}
   );
   gpc1_1 gpc757 (
      {stage0_59[38]},
      {stage1_59[19]}
   );
   gpc1_1 gpc758 (
      {stage0_59[39]},
      {stage1_59[20]}
   );
   gpc1_1 gpc759 (
      {stage0_59[40]},
      {stage1_59[21]}
   );
   gpc1_1 gpc760 (
      {stage0_59[41]},
      {stage1_59[22]}
   );
   gpc1_1 gpc761 (
      {stage0_59[42]},
      {stage1_59[23]}
   );
   gpc1_1 gpc762 (
      {stage0_59[43]},
      {stage1_59[24]}
   );
   gpc1_1 gpc763 (
      {stage0_59[44]},
      {stage1_59[25]}
   );
   gpc1_1 gpc764 (
      {stage0_59[45]},
      {stage1_59[26]}
   );
   gpc1_1 gpc765 (
      {stage0_59[46]},
      {stage1_59[27]}
   );
   gpc1_1 gpc766 (
      {stage0_59[47]},
      {stage1_59[28]}
   );
   gpc1_1 gpc767 (
      {stage0_59[48]},
      {stage1_59[29]}
   );
   gpc1_1 gpc768 (
      {stage0_59[49]},
      {stage1_59[30]}
   );
   gpc1_1 gpc769 (
      {stage0_59[50]},
      {stage1_59[31]}
   );
   gpc1_1 gpc770 (
      {stage0_59[51]},
      {stage1_59[32]}
   );
   gpc1_1 gpc771 (
      {stage0_59[52]},
      {stage1_59[33]}
   );
   gpc1_1 gpc772 (
      {stage0_59[53]},
      {stage1_59[34]}
   );
   gpc1_1 gpc773 (
      {stage0_62[48]},
      {stage1_62[18]}
   );
   gpc1_1 gpc774 (
      {stage0_62[49]},
      {stage1_62[19]}
   );
   gpc1_1 gpc775 (
      {stage0_62[50]},
      {stage1_62[20]}
   );
   gpc1_1 gpc776 (
      {stage0_62[51]},
      {stage1_62[21]}
   );
   gpc1_1 gpc777 (
      {stage0_62[52]},
      {stage1_62[22]}
   );
   gpc1_1 gpc778 (
      {stage0_62[53]},
      {stage1_62[23]}
   );
   gpc1_1 gpc779 (
      {stage0_63[36]},
      {stage1_63[17]}
   );
   gpc1_1 gpc780 (
      {stage0_63[37]},
      {stage1_63[18]}
   );
   gpc1_1 gpc781 (
      {stage0_63[38]},
      {stage1_63[19]}
   );
   gpc1_1 gpc782 (
      {stage0_63[39]},
      {stage1_63[20]}
   );
   gpc1_1 gpc783 (
      {stage0_63[40]},
      {stage1_63[21]}
   );
   gpc1_1 gpc784 (
      {stage0_63[41]},
      {stage1_63[22]}
   );
   gpc1_1 gpc785 (
      {stage0_63[42]},
      {stage1_63[23]}
   );
   gpc1_1 gpc786 (
      {stage0_63[43]},
      {stage1_63[24]}
   );
   gpc1_1 gpc787 (
      {stage0_63[44]},
      {stage1_63[25]}
   );
   gpc1_1 gpc788 (
      {stage0_63[45]},
      {stage1_63[26]}
   );
   gpc1_1 gpc789 (
      {stage0_63[46]},
      {stage1_63[27]}
   );
   gpc1_1 gpc790 (
      {stage0_63[47]},
      {stage1_63[28]}
   );
   gpc1_1 gpc791 (
      {stage0_63[48]},
      {stage1_63[29]}
   );
   gpc1_1 gpc792 (
      {stage0_63[49]},
      {stage1_63[30]}
   );
   gpc1_1 gpc793 (
      {stage0_63[50]},
      {stage1_63[31]}
   );
   gpc1_1 gpc794 (
      {stage0_63[51]},
      {stage1_63[32]}
   );
   gpc1_1 gpc795 (
      {stage0_63[52]},
      {stage1_63[33]}
   );
   gpc1_1 gpc796 (
      {stage0_63[53]},
      {stage1_63[34]}
   );
   gpc1163_5 gpc797 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc798 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc799 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[6]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc800 (
      {stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage1_3[1]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc801 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc802 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[5],stage2_3[5]}
   );
   gpc615_5 gpc803 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[3]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc804 (
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage1_4[4]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc2135_5 gpc805 (
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[5],stage2_4[8]}
   );
   gpc2135_5 gpc806 (
      {stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_6[1]},
      {stage1_7[2], stage1_7[3]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc807 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc808 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage2_9[0],stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[8]}
   );
   gpc606_5 gpc809 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage2_9[1],stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[9]}
   );
   gpc615_5 gpc810 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[16]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[5],stage2_7[8],stage2_6[8]}
   );
   gpc615_5 gpc811 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[17]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[6],stage2_7[9],stage2_6[9]}
   );
   gpc615_5 gpc812 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[4],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc813 (
      {stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[3],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc814 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[4],stage2_9[6],stage2_8[9]}
   );
   gpc606_5 gpc815 (
      {stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[5],stage2_9[7],stage2_8[10]}
   );
   gpc615_5 gpc816 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[0]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[3],stage2_11[4],stage2_10[6]}
   );
   gpc1415_5 gpc817 (
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[4],stage2_11[5]}
   );
   gpc1415_5 gpc818 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[7]},
      {stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[5],stage2_11[6]}
   );
   gpc1163_5 gpc819 (
      {stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_13[8]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[6],stage2_11[7]}
   );
   gpc1163_5 gpc820 (
      {stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_13[9]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[7],stage2_11[8]}
   );
   gpc615_5 gpc821 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[20]},
      {stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[8],stage2_11[9]}
   );
   gpc615_5 gpc822 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {1'b0},
      {stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[9],stage2_11[10]}
   );
   gpc606_5 gpc823 (
      {stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[6],stage2_14[7],stage2_13[7]}
   );
   gpc1343_5 gpc824 (
      {stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage1_16[0], stage1_16[1], stage1_16[2]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[7],stage2_14[8]}
   );
   gpc1343_5 gpc825 (
      {stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[8],stage2_14[9]}
   );
   gpc1163_5 gpc826 (
      {stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_16[6]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[9],stage2_14[10]}
   );
   gpc1163_5 gpc827 (
      {stage1_14[13], stage1_14[14], stage1_14[15]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_16[7]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[4],stage2_16[4],stage2_15[10],stage2_14[11]}
   );
   gpc1163_5 gpc828 (
      {stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_16[8]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[5],stage2_16[5],stage2_15[11],stage2_14[12]}
   );
   gpc1163_5 gpc829 (
      {stage1_14[19], stage1_14[20], stage1_14[21]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[9]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[6],stage2_16[6],stage2_15[12],stage2_14[13]}
   );
   gpc1163_5 gpc830 (
      {stage1_14[22], stage1_14[23], 1'b0},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], 1'b0},
      {stage1_16[10]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[7],stage2_16[7],stage2_15[13],stage2_14[14]}
   );
   gpc606_5 gpc831 (
      {stage1_16[11], stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[7],stage2_17[8],stage2_16[8]}
   );
   gpc606_5 gpc832 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[8],stage2_17[9],stage2_16[9]}
   );
   gpc606_5 gpc833 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[9],stage2_17[10]}
   );
   gpc615_5 gpc834 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_18[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[10],stage2_17[11]}
   );
   gpc615_5 gpc835 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_19[12]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[11]}
   );
   gpc615_5 gpc836 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage1_19[13]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[12]}
   );
   gpc615_5 gpc837 (
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27]},
      {stage1_19[14]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[13]}
   );
   gpc615_5 gpc838 (
      {stage1_19[15], stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[5],stage2_20[7],stage2_19[7]}
   );
   gpc1343_5 gpc839 (
      {stage1_21[6], stage1_21[7], stage1_21[8]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3]},
      {stage1_23[0], stage1_23[1], stage1_23[2]},
      {stage1_24[0]},
      {stage2_25[0],stage2_24[0],stage2_23[1],stage2_22[4],stage2_21[6]}
   );
   gpc1343_5 gpc840 (
      {stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage1_22[4], stage1_22[5], stage1_22[6], stage1_22[7]},
      {stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage1_24[1]},
      {stage2_25[1],stage2_24[1],stage2_23[2],stage2_22[5],stage2_21[7]}
   );
   gpc606_5 gpc841 (
      {stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11], stage1_22[12], stage1_22[13]},
      {stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7]},
      {stage2_26[0],stage2_25[2],stage2_24[2],stage2_23[3],stage2_22[6]}
   );
   gpc606_5 gpc842 (
      {stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17], stage1_22[18], stage1_22[19]},
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage2_26[1],stage2_25[3],stage2_24[3],stage2_23[4],stage2_22[7]}
   );
   gpc615_5 gpc843 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage1_25[0]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[4],stage2_24[4]}
   );
   gpc615_5 gpc844 (
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage1_25[1]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[5],stage2_24[5]}
   );
   gpc615_5 gpc845 (
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28]},
      {stage1_25[2]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[6],stage2_24[6]}
   );
   gpc615_5 gpc846 (
      {stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage1_26[18]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[7]}
   );
   gpc615_5 gpc847 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage1_26[19]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[4],stage2_27[4],stage2_26[6],stage2_25[8]}
   );
   gpc615_5 gpc848 (
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage1_26[20]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[5],stage2_27[5],stage2_26[7],stage2_25[9]}
   );
   gpc615_5 gpc849 (
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22]},
      {stage1_26[21]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[6],stage2_27[6],stage2_26[8],stage2_25[10]}
   );
   gpc1343_5 gpc850 (
      {stage1_28[0], stage1_28[1], stage1_28[2]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage2_32[0],stage2_31[0],stage2_30[0],stage2_29[4],stage2_28[7]}
   );
   gpc1343_5 gpc851 (
      {stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_29[4], stage1_29[5], stage1_29[6], stage1_29[7]},
      {stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_31[1]},
      {stage2_32[1],stage2_31[1],stage2_30[1],stage2_29[5],stage2_28[8]}
   );
   gpc1343_5 gpc852 (
      {stage1_28[6], stage1_28[7], stage1_28[8]},
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_31[2]},
      {stage2_32[2],stage2_31[2],stage2_30[2],stage2_29[6],stage2_28[9]}
   );
   gpc606_5 gpc853 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage2_32[3],stage2_31[3],stage2_30[3],stage2_29[7],stage2_28[10]}
   );
   gpc615_5 gpc854 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_30[15]},
      {stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8]},
      {stage2_33[0],stage2_32[4],stage2_31[4],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc855 (
      {stage1_30[16], stage1_30[17], stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[5],stage2_31[5],stage2_30[5]}
   );
   gpc606_5 gpc856 (
      {stage1_30[22], stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[2],stage2_32[6],stage2_31[6],stage2_30[6]}
   );
   gpc615_5 gpc857 (
      {stage1_30[28], stage1_30[29], stage1_30[30], stage1_30[31], stage1_30[32]},
      {stage1_31[9]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[3],stage2_32[7],stage2_31[7],stage2_30[7]}
   );
   gpc606_5 gpc858 (
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[3],stage2_33[4],stage2_32[8],stage2_31[8]}
   );
   gpc606_5 gpc859 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[4],stage2_33[5],stage2_32[9],stage2_31[9]}
   );
   gpc606_5 gpc860 (
      {stage1_31[22], stage1_31[23], stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[5],stage2_33[6],stage2_32[10],stage2_31[10]}
   );
   gpc606_5 gpc861 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[0],stage2_35[3],stage2_34[6],stage2_33[7]}
   );
   gpc606_5 gpc862 (
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[1],stage2_35[4],stage2_34[7],stage2_33[8]}
   );
   gpc606_5 gpc863 (
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[2],stage2_35[5],stage2_34[8],stage2_33[9]}
   );
   gpc615_5 gpc864 (
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40]},
      {stage1_34[0]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[3],stage2_35[6],stage2_34[9],stage2_33[10]}
   );
   gpc615_5 gpc865 (
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage1_35[24]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[4],stage2_36[4],stage2_35[7],stage2_34[10]}
   );
   gpc615_5 gpc866 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[25]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[5],stage2_36[5],stage2_35[8],stage2_34[11]}
   );
   gpc615_5 gpc867 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[26]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[6],stage2_36[6],stage2_35[9],stage2_34[12]}
   );
   gpc615_5 gpc868 (
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22]},
      {stage1_37[0]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[0],stage2_38[3],stage2_37[7],stage2_36[7]}
   );
   gpc606_5 gpc869 (
      {stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5], stage1_37[6]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[4],stage2_37[8]}
   );
   gpc606_5 gpc870 (
      {stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11], stage1_37[12]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[5],stage2_37[9]}
   );
   gpc606_5 gpc871 (
      {stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17], stage1_37[18]},
      {stage1_39[12], stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17]},
      {stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[6],stage2_37[10]}
   );
   gpc615_5 gpc872 (
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10]},
      {stage1_39[18]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[3],stage2_40[4],stage2_39[4],stage2_38[7]}
   );
   gpc615_5 gpc873 (
      {stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage1_39[19]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[4],stage2_40[5],stage2_39[5],stage2_38[8]}
   );
   gpc615_5 gpc874 (
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage1_39[20]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[5],stage2_40[6],stage2_39[6],stage2_38[9]}
   );
   gpc1163_5 gpc875 (
      {stage1_40[18], stage1_40[19], stage1_40[20]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_42[0]},
      {stage1_43[0]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[6],stage2_40[7]}
   );
   gpc1163_5 gpc876 (
      {stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_42[1]},
      {stage1_43[1]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[7],stage2_40[8]}
   );
   gpc1163_5 gpc877 (
      {stage1_40[24], stage1_40[25], stage1_40[26]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_42[2]},
      {stage1_43[2]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[8],stage2_40[9]}
   );
   gpc606_5 gpc878 (
      {stage1_40[27], stage1_40[28], stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32]},
      {stage1_42[3], stage1_42[4], stage1_42[5], stage1_42[6], stage1_42[7], stage1_42[8]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[9],stage2_40[10]}
   );
   gpc606_5 gpc879 (
      {stage1_40[33], stage1_40[34], stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38]},
      {stage1_42[9], stage1_42[10], stage1_42[11], stage1_42[12], stage1_42[13], stage1_42[14]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[10],stage2_40[11]}
   );
   gpc606_5 gpc880 (
      {stage1_43[3], stage1_43[4], stage1_43[5], stage1_43[6], stage1_43[7], stage1_43[8]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[0],stage2_44[5],stage2_43[5]}
   );
   gpc606_5 gpc881 (
      {stage1_43[9], stage1_43[10], stage1_43[11], stage1_43[12], stage1_43[13], stage1_43[14]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[1],stage2_44[6],stage2_43[6]}
   );
   gpc606_5 gpc882 (
      {stage1_43[15], stage1_43[16], stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[2],stage2_44[7],stage2_43[7]}
   );
   gpc606_5 gpc883 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[3],stage2_46[3],stage2_45[3],stage2_44[8]}
   );
   gpc606_5 gpc884 (
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[4],stage2_46[4],stage2_45[4],stage2_44[9]}
   );
   gpc606_5 gpc885 (
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[5],stage2_46[5],stage2_45[5],stage2_44[10]}
   );
   gpc615_5 gpc886 (
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22]},
      {stage1_46[18]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[6],stage2_46[6],stage2_45[6]}
   );
   gpc615_5 gpc887 (
      {stage1_45[23], stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27]},
      {stage1_46[19]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[7],stage2_46[7],stage2_45[7]}
   );
   gpc615_5 gpc888 (
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16]},
      {stage1_48[0]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[2],stage2_48[5],stage2_47[8]}
   );
   gpc615_5 gpc889 (
      {stage1_47[17], stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21]},
      {stage1_48[1]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[3],stage2_48[6],stage2_47[9]}
   );
   gpc606_5 gpc890 (
      {stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6], stage1_48[7]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[2],stage2_50[2],stage2_49[4],stage2_48[7]}
   );
   gpc606_5 gpc891 (
      {stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[3],stage2_50[3],stage2_49[5],stage2_48[8]}
   );
   gpc2135_5 gpc892 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16]},
      {stage1_51[0], stage1_51[1], stage1_51[2]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[0],stage2_52[2],stage2_51[4],stage2_50[4]}
   );
   gpc2135_5 gpc893 (
      {stage1_50[17], stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21]},
      {stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[1]},
      {stage1_53[2], stage1_53[3]},
      {stage2_54[1],stage2_53[1],stage2_52[3],stage2_51[5],stage2_50[5]}
   );
   gpc2135_5 gpc894 (
      {stage1_50[22], stage1_50[23], stage1_50[24], stage1_50[25], stage1_50[26]},
      {stage1_51[6], stage1_51[7], stage1_51[8]},
      {stage1_52[2]},
      {stage1_53[4], stage1_53[5]},
      {stage2_54[2],stage2_53[2],stage2_52[4],stage2_51[6],stage2_50[6]}
   );
   gpc2135_5 gpc895 (
      {stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30], stage1_50[31]},
      {stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage1_52[3]},
      {stage1_53[6], stage1_53[7]},
      {stage2_54[3],stage2_53[3],stage2_52[5],stage2_51[7],stage2_50[7]}
   );
   gpc2135_5 gpc896 (
      {stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_51[12], stage1_51[13], stage1_51[14]},
      {stage1_52[4]},
      {stage1_53[8], stage1_53[9]},
      {stage2_54[4],stage2_53[4],stage2_52[6],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc897 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[15]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[5],stage2_52[7],stage2_51[9],stage2_50[9]}
   );
   gpc606_5 gpc898 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15]},
      {stage2_55[0],stage2_54[6],stage2_53[6],stage2_52[8],stage2_51[10]}
   );
   gpc606_5 gpc899 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27]},
      {stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage2_55[1],stage2_54[7],stage2_53[7],stage2_52[9],stage2_51[11]}
   );
   gpc606_5 gpc900 (
      {stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33]},
      {stage1_53[22], stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27]},
      {stage2_55[2],stage2_54[8],stage2_53[8],stage2_52[10],stage2_51[12]}
   );
   gpc606_5 gpc901 (
      {stage1_51[34], stage1_51[35], stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39]},
      {stage1_53[28], stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33]},
      {stage2_55[3],stage2_54[9],stage2_53[9],stage2_52[11],stage2_51[13]}
   );
   gpc606_5 gpc902 (
      {stage1_51[40], stage1_51[41], stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45]},
      {stage1_53[34], stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage2_55[4],stage2_54[10],stage2_53[10],stage2_52[12],stage2_51[14]}
   );
   gpc606_5 gpc903 (
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[5],stage2_54[11],stage2_53[11],stage2_52[13]}
   );
   gpc615_5 gpc904 (
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10]},
      {stage1_55[0]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[0],stage2_56[1],stage2_55[6],stage2_54[12]}
   );
   gpc615_5 gpc905 (
      {stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage1_55[1]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[1],stage2_56[2],stage2_55[7],stage2_54[13]}
   );
   gpc606_5 gpc906 (
      {stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5], stage1_55[6], stage1_55[7]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[2],stage2_56[3],stage2_55[8]}
   );
   gpc606_5 gpc907 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12], stage1_55[13]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[3],stage2_56[4],stage2_55[9]}
   );
   gpc606_5 gpc908 (
      {stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17], stage1_55[18], stage1_55[19]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[4],stage2_56[5],stage2_55[10]}
   );
   gpc606_5 gpc909 (
      {stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23], stage1_55[24], stage1_55[25]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[5],stage2_56[6],stage2_55[11]}
   );
   gpc606_5 gpc910 (
      {stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[6],stage2_56[7],stage2_55[12]}
   );
   gpc615_5 gpc911 (
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16]},
      {stage1_57[30]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[5],stage2_58[7],stage2_57[7],stage2_56[8]}
   );
   gpc606_5 gpc912 (
      {stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35], stage1_57[36]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[1],stage2_59[6],stage2_58[8],stage2_57[8]}
   );
   gpc135_4 gpc913 (
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10]},
      {stage1_60[0], stage1_60[1], stage1_60[2]},
      {stage1_61[0]},
      {stage2_62[0],stage2_61[1],stage2_60[2],stage2_59[7]}
   );
   gpc135_4 gpc914 (
      {stage1_59[11], stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15]},
      {stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage1_61[1]},
      {stage2_62[1],stage2_61[2],stage2_60[3],stage2_59[8]}
   );
   gpc135_4 gpc915 (
      {stage1_59[16], stage1_59[17], stage1_59[18], stage1_59[19], stage1_59[20]},
      {stage1_60[6], stage1_60[7], stage1_60[8]},
      {stage1_61[2]},
      {stage2_62[2],stage2_61[3],stage2_60[4],stage2_59[9]}
   );
   gpc135_4 gpc916 (
      {stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24], stage1_59[25]},
      {stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage1_61[3]},
      {stage2_62[3],stage2_61[4],stage2_60[5],stage2_59[10]}
   );
   gpc135_4 gpc917 (
      {stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30]},
      {stage1_60[12], stage1_60[13], stage1_60[14]},
      {stage1_61[4]},
      {stage2_62[4],stage2_61[5],stage2_60[6],stage2_59[11]}
   );
   gpc135_4 gpc918 (
      {stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], 1'b0},
      {stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage1_61[5]},
      {stage2_62[5],stage2_61[6],stage2_60[7],stage2_59[12]}
   );
   gpc606_5 gpc919 (
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[0],stage2_63[0],stage2_62[6],stage2_61[7]}
   );
   gpc606_5 gpc920 (
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[1],stage2_63[1],stage2_62[7],stage2_61[8]}
   );
   gpc1163_5 gpc921 (
      {stage1_62[0], stage1_62[1], stage1_62[2]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[2],stage2_64[2],stage2_63[2],stage2_62[8]}
   );
   gpc1163_5 gpc922 (
      {stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[3],stage2_64[3],stage2_63[3],stage2_62[9]}
   );
   gpc606_5 gpc923 (
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7]},
      {stage2_66[2],stage2_65[4],stage2_64[4],stage2_63[4],stage2_62[10]}
   );
   gpc606_5 gpc924 (
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13]},
      {stage2_66[3],stage2_65[5],stage2_64[5],stage2_63[5],stage2_62[11]}
   );
   gpc1_1 gpc925 (
      {stage1_0[14]},
      {stage2_0[3]}
   );
   gpc1_1 gpc926 (
      {stage1_0[15]},
      {stage2_0[4]}
   );
   gpc1_1 gpc927 (
      {stage1_0[16]},
      {stage2_0[5]}
   );
   gpc1_1 gpc928 (
      {stage1_1[18]},
      {stage2_1[5]}
   );
   gpc1_1 gpc929 (
      {stage1_1[19]},
      {stage2_1[6]}
   );
   gpc1_1 gpc930 (
      {stage1_2[16]},
      {stage2_2[5]}
   );
   gpc1_1 gpc931 (
      {stage1_2[17]},
      {stage2_2[6]}
   );
   gpc1_1 gpc932 (
      {stage1_2[18]},
      {stage2_2[7]}
   );
   gpc1_1 gpc933 (
      {stage1_2[19]},
      {stage2_2[8]}
   );
   gpc1_1 gpc934 (
      {stage1_2[20]},
      {stage2_2[9]}
   );
   gpc1_1 gpc935 (
      {stage1_2[21]},
      {stage2_2[10]}
   );
   gpc1_1 gpc936 (
      {stage1_2[22]},
      {stage2_2[11]}
   );
   gpc1_1 gpc937 (
      {stage1_2[23]},
      {stage2_2[12]}
   );
   gpc1_1 gpc938 (
      {stage1_2[24]},
      {stage2_2[13]}
   );
   gpc1_1 gpc939 (
      {stage1_3[23]},
      {stage2_3[8]}
   );
   gpc1_1 gpc940 (
      {stage1_4[21]},
      {stage2_4[11]}
   );
   gpc1_1 gpc941 (
      {stage1_4[22]},
      {stage2_4[12]}
   );
   gpc1_1 gpc942 (
      {stage1_4[23]},
      {stage2_4[13]}
   );
   gpc1_1 gpc943 (
      {stage1_4[24]},
      {stage2_4[14]}
   );
   gpc1_1 gpc944 (
      {stage1_4[25]},
      {stage2_4[15]}
   );
   gpc1_1 gpc945 (
      {stage1_4[26]},
      {stage2_4[16]}
   );
   gpc1_1 gpc946 (
      {stage1_4[27]},
      {stage2_4[17]}
   );
   gpc1_1 gpc947 (
      {stage1_4[28]},
      {stage2_4[18]}
   );
   gpc1_1 gpc948 (
      {stage1_4[29]},
      {stage2_4[19]}
   );
   gpc1_1 gpc949 (
      {stage1_4[30]},
      {stage2_4[20]}
   );
   gpc1_1 gpc950 (
      {stage1_4[31]},
      {stage2_4[21]}
   );
   gpc1_1 gpc951 (
      {stage1_4[32]},
      {stage2_4[22]}
   );
   gpc1_1 gpc952 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc953 (
      {stage1_7[23]},
      {stage2_7[11]}
   );
   gpc1_1 gpc954 (
      {stage1_7[24]},
      {stage2_7[12]}
   );
   gpc1_1 gpc955 (
      {stage1_9[6]},
      {stage2_9[8]}
   );
   gpc1_1 gpc956 (
      {stage1_9[7]},
      {stage2_9[9]}
   );
   gpc1_1 gpc957 (
      {stage1_9[8]},
      {stage2_9[10]}
   );
   gpc1_1 gpc958 (
      {stage1_9[9]},
      {stage2_9[11]}
   );
   gpc1_1 gpc959 (
      {stage1_9[10]},
      {stage2_9[12]}
   );
   gpc1_1 gpc960 (
      {stage1_9[11]},
      {stage2_9[13]}
   );
   gpc1_1 gpc961 (
      {stage1_9[12]},
      {stage2_9[14]}
   );
   gpc1_1 gpc962 (
      {stage1_9[13]},
      {stage2_9[15]}
   );
   gpc1_1 gpc963 (
      {stage1_9[14]},
      {stage2_9[16]}
   );
   gpc1_1 gpc964 (
      {stage1_9[15]},
      {stage2_9[17]}
   );
   gpc1_1 gpc965 (
      {stage1_9[16]},
      {stage2_9[18]}
   );
   gpc1_1 gpc966 (
      {stage1_9[17]},
      {stage2_9[19]}
   );
   gpc1_1 gpc967 (
      {stage1_10[23]},
      {stage2_10[7]}
   );
   gpc1_1 gpc968 (
      {stage1_10[24]},
      {stage2_10[8]}
   );
   gpc1_1 gpc969 (
      {stage1_10[25]},
      {stage2_10[9]}
   );
   gpc1_1 gpc970 (
      {stage1_11[27]},
      {stage2_11[11]}
   );
   gpc1_1 gpc971 (
      {stage1_11[28]},
      {stage2_11[12]}
   );
   gpc1_1 gpc972 (
      {stage1_13[28]},
      {stage2_13[8]}
   );
   gpc1_1 gpc973 (
      {stage1_13[29]},
      {stage2_13[9]}
   );
   gpc1_1 gpc974 (
      {stage1_16[23]},
      {stage2_16[10]}
   );
   gpc1_1 gpc975 (
      {stage1_18[28]},
      {stage2_18[14]}
   );
   gpc1_1 gpc976 (
      {stage1_18[29]},
      {stage2_18[15]}
   );
   gpc1_1 gpc977 (
      {stage1_18[30]},
      {stage2_18[16]}
   );
   gpc1_1 gpc978 (
      {stage1_18[31]},
      {stage2_18[17]}
   );
   gpc1_1 gpc979 (
      {stage1_18[32]},
      {stage2_18[18]}
   );
   gpc1_1 gpc980 (
      {stage1_18[33]},
      {stage2_18[19]}
   );
   gpc1_1 gpc981 (
      {stage1_19[20]},
      {stage2_19[8]}
   );
   gpc1_1 gpc982 (
      {stage1_20[19]},
      {stage2_20[8]}
   );
   gpc1_1 gpc983 (
      {stage1_21[12]},
      {stage2_21[8]}
   );
   gpc1_1 gpc984 (
      {stage1_21[13]},
      {stage2_21[9]}
   );
   gpc1_1 gpc985 (
      {stage1_21[14]},
      {stage2_21[10]}
   );
   gpc1_1 gpc986 (
      {stage1_21[15]},
      {stage2_21[11]}
   );
   gpc1_1 gpc987 (
      {stage1_21[16]},
      {stage2_21[12]}
   );
   gpc1_1 gpc988 (
      {stage1_21[17]},
      {stage2_21[13]}
   );
   gpc1_1 gpc989 (
      {stage1_21[18]},
      {stage2_21[14]}
   );
   gpc1_1 gpc990 (
      {stage1_21[19]},
      {stage2_21[15]}
   );
   gpc1_1 gpc991 (
      {stage1_21[20]},
      {stage2_21[16]}
   );
   gpc1_1 gpc992 (
      {stage1_21[21]},
      {stage2_21[17]}
   );
   gpc1_1 gpc993 (
      {stage1_21[22]},
      {stage2_21[18]}
   );
   gpc1_1 gpc994 (
      {stage1_21[23]},
      {stage2_21[19]}
   );
   gpc1_1 gpc995 (
      {stage1_21[24]},
      {stage2_21[20]}
   );
   gpc1_1 gpc996 (
      {stage1_21[25]},
      {stage2_21[21]}
   );
   gpc1_1 gpc997 (
      {stage1_22[20]},
      {stage2_22[8]}
   );
   gpc1_1 gpc998 (
      {stage1_22[21]},
      {stage2_22[9]}
   );
   gpc1_1 gpc999 (
      {stage1_22[22]},
      {stage2_22[10]}
   );
   gpc1_1 gpc1000 (
      {stage1_23[6]},
      {stage2_23[5]}
   );
   gpc1_1 gpc1001 (
      {stage1_23[7]},
      {stage2_23[6]}
   );
   gpc1_1 gpc1002 (
      {stage1_23[8]},
      {stage2_23[7]}
   );
   gpc1_1 gpc1003 (
      {stage1_23[9]},
      {stage2_23[8]}
   );
   gpc1_1 gpc1004 (
      {stage1_23[10]},
      {stage2_23[9]}
   );
   gpc1_1 gpc1005 (
      {stage1_23[11]},
      {stage2_23[10]}
   );
   gpc1_1 gpc1006 (
      {stage1_23[12]},
      {stage2_23[11]}
   );
   gpc1_1 gpc1007 (
      {stage1_23[13]},
      {stage2_23[12]}
   );
   gpc1_1 gpc1008 (
      {stage1_23[14]},
      {stage2_23[13]}
   );
   gpc1_1 gpc1009 (
      {stage1_23[15]},
      {stage2_23[14]}
   );
   gpc1_1 gpc1010 (
      {stage1_23[16]},
      {stage2_23[15]}
   );
   gpc1_1 gpc1011 (
      {stage1_23[17]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1012 (
      {stage1_23[18]},
      {stage2_23[17]}
   );
   gpc1_1 gpc1013 (
      {stage1_23[19]},
      {stage2_23[18]}
   );
   gpc1_1 gpc1014 (
      {stage1_23[20]},
      {stage2_23[19]}
   );
   gpc1_1 gpc1015 (
      {stage1_23[21]},
      {stage2_23[20]}
   );
   gpc1_1 gpc1016 (
      {stage1_24[29]},
      {stage2_24[7]}
   );
   gpc1_1 gpc1017 (
      {stage1_24[30]},
      {stage2_24[8]}
   );
   gpc1_1 gpc1018 (
      {stage1_24[31]},
      {stage2_24[9]}
   );
   gpc1_1 gpc1019 (
      {stage1_25[23]},
      {stage2_25[11]}
   );
   gpc1_1 gpc1020 (
      {stage1_25[24]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1021 (
      {stage1_26[22]},
      {stage2_26[9]}
   );
   gpc1_1 gpc1022 (
      {stage1_26[23]},
      {stage2_26[10]}
   );
   gpc1_1 gpc1023 (
      {stage1_26[24]},
      {stage2_26[11]}
   );
   gpc1_1 gpc1024 (
      {stage1_26[25]},
      {stage2_26[12]}
   );
   gpc1_1 gpc1025 (
      {stage1_26[26]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1026 (
      {stage1_26[27]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1027 (
      {stage1_26[28]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1028 (
      {stage1_26[29]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1029 (
      {stage1_26[30]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1030 (
      {stage1_26[31]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1031 (
      {stage1_28[15]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1032 (
      {stage1_28[16]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1033 (
      {stage1_28[17]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1034 (
      {stage1_29[17]},
      {stage2_29[9]}
   );
   gpc1_1 gpc1035 (
      {stage1_29[18]},
      {stage2_29[10]}
   );
   gpc1_1 gpc1036 (
      {stage1_29[19]},
      {stage2_29[11]}
   );
   gpc1_1 gpc1037 (
      {stage1_29[20]},
      {stage2_29[12]}
   );
   gpc1_1 gpc1038 (
      {stage1_29[21]},
      {stage2_29[13]}
   );
   gpc1_1 gpc1039 (
      {stage1_29[22]},
      {stage2_29[14]}
   );
   gpc1_1 gpc1040 (
      {stage1_29[23]},
      {stage2_29[15]}
   );
   gpc1_1 gpc1041 (
      {stage1_29[24]},
      {stage2_29[16]}
   );
   gpc1_1 gpc1042 (
      {stage1_29[25]},
      {stage2_29[17]}
   );
   gpc1_1 gpc1043 (
      {stage1_30[33]},
      {stage2_30[8]}
   );
   gpc1_1 gpc1044 (
      {stage1_30[34]},
      {stage2_30[9]}
   );
   gpc1_1 gpc1045 (
      {stage1_31[28]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1046 (
      {stage1_31[29]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1047 (
      {stage1_31[30]},
      {stage2_31[13]}
   );
   gpc1_1 gpc1048 (
      {stage1_31[31]},
      {stage2_31[14]}
   );
   gpc1_1 gpc1049 (
      {stage1_31[32]},
      {stage2_31[15]}
   );
   gpc1_1 gpc1050 (
      {stage1_31[33]},
      {stage2_31[16]}
   );
   gpc1_1 gpc1051 (
      {stage1_32[18]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1052 (
      {stage1_33[41]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1053 (
      {stage1_33[42]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1054 (
      {stage1_33[43]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1055 (
      {stage1_33[44]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1056 (
      {stage1_33[45]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1057 (
      {stage1_34[16]},
      {stage2_34[13]}
   );
   gpc1_1 gpc1058 (
      {stage1_34[17]},
      {stage2_34[14]}
   );
   gpc1_1 gpc1059 (
      {stage1_34[18]},
      {stage2_34[15]}
   );
   gpc1_1 gpc1060 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1061 (
      {stage1_36[23]},
      {stage2_36[8]}
   );
   gpc1_1 gpc1062 (
      {stage1_36[24]},
      {stage2_36[9]}
   );
   gpc1_1 gpc1063 (
      {stage1_36[25]},
      {stage2_36[10]}
   );
   gpc1_1 gpc1064 (
      {stage1_36[26]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1065 (
      {stage1_36[27]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1066 (
      {stage1_36[28]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1067 (
      {stage1_36[29]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1068 (
      {stage1_36[30]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1069 (
      {stage1_36[31]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1070 (
      {stage1_36[32]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1071 (
      {stage1_36[33]},
      {stage2_36[18]}
   );
   gpc1_1 gpc1072 (
      {stage1_37[19]},
      {stage2_37[11]}
   );
   gpc1_1 gpc1073 (
      {stage1_37[20]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1074 (
      {stage1_37[21]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1075 (
      {stage1_37[22]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1076 (
      {stage1_37[23]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1077 (
      {stage1_37[24]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1078 (
      {stage1_38[21]},
      {stage2_38[10]}
   );
   gpc1_1 gpc1079 (
      {stage1_38[22]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1080 (
      {stage1_38[23]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1081 (
      {stage1_39[21]},
      {stage2_39[7]}
   );
   gpc1_1 gpc1082 (
      {stage1_39[22]},
      {stage2_39[8]}
   );
   gpc1_1 gpc1083 (
      {stage1_39[23]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_39[24]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_39[25]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_39[26]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_39[27]},
      {stage2_39[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_39[28]},
      {stage2_39[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_39[29]},
      {stage2_39[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_39[30]},
      {stage2_39[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_41[18]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1092 (
      {stage1_41[19]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1093 (
      {stage1_42[15]},
      {stage2_42[8]}
   );
   gpc1_1 gpc1094 (
      {stage1_42[16]},
      {stage2_42[9]}
   );
   gpc1_1 gpc1095 (
      {stage1_42[17]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1096 (
      {stage1_42[18]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1097 (
      {stage1_42[19]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1098 (
      {stage1_42[20]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1099 (
      {stage1_43[21]},
      {stage2_43[8]}
   );
   gpc1_1 gpc1100 (
      {stage1_43[22]},
      {stage2_43[9]}
   );
   gpc1_1 gpc1101 (
      {stage1_44[18]},
      {stage2_44[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_44[19]},
      {stage2_44[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_44[20]},
      {stage2_44[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_44[21]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_45[28]},
      {stage2_45[8]}
   );
   gpc1_1 gpc1106 (
      {stage1_45[29]},
      {stage2_45[9]}
   );
   gpc1_1 gpc1107 (
      {stage1_45[30]},
      {stage2_45[10]}
   );
   gpc1_1 gpc1108 (
      {stage1_45[31]},
      {stage2_45[11]}
   );
   gpc1_1 gpc1109 (
      {stage1_46[20]},
      {stage2_46[8]}
   );
   gpc1_1 gpc1110 (
      {stage1_46[21]},
      {stage2_46[9]}
   );
   gpc1_1 gpc1111 (
      {stage1_46[22]},
      {stage2_46[10]}
   );
   gpc1_1 gpc1112 (
      {stage1_46[23]},
      {stage2_46[11]}
   );
   gpc1_1 gpc1113 (
      {stage1_46[24]},
      {stage2_46[12]}
   );
   gpc1_1 gpc1114 (
      {stage1_46[25]},
      {stage2_46[13]}
   );
   gpc1_1 gpc1115 (
      {stage1_46[26]},
      {stage2_46[14]}
   );
   gpc1_1 gpc1116 (
      {stage1_46[27]},
      {stage2_46[15]}
   );
   gpc1_1 gpc1117 (
      {stage1_46[28]},
      {stage2_46[16]}
   );
   gpc1_1 gpc1118 (
      {stage1_46[29]},
      {stage2_46[17]}
   );
   gpc1_1 gpc1119 (
      {stage1_47[22]},
      {stage2_47[10]}
   );
   gpc1_1 gpc1120 (
      {stage1_47[23]},
      {stage2_47[11]}
   );
   gpc1_1 gpc1121 (
      {stage1_47[24]},
      {stage2_47[12]}
   );
   gpc1_1 gpc1122 (
      {stage1_47[25]},
      {stage2_47[13]}
   );
   gpc1_1 gpc1123 (
      {stage1_47[26]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1124 (
      {stage1_47[27]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1125 (
      {stage1_47[28]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1126 (
      {stage1_47[29]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1127 (
      {stage1_47[30]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1128 (
      {stage1_47[31]},
      {stage2_47[19]}
   );
   gpc1_1 gpc1129 (
      {stage1_47[32]},
      {stage2_47[20]}
   );
   gpc1_1 gpc1130 (
      {stage1_47[33]},
      {stage2_47[21]}
   );
   gpc1_1 gpc1131 (
      {stage1_48[14]},
      {stage2_48[9]}
   );
   gpc1_1 gpc1132 (
      {stage1_48[15]},
      {stage2_48[10]}
   );
   gpc1_1 gpc1133 (
      {stage1_48[16]},
      {stage2_48[11]}
   );
   gpc1_1 gpc1134 (
      {stage1_48[17]},
      {stage2_48[12]}
   );
   gpc1_1 gpc1135 (
      {stage1_49[12]},
      {stage2_49[6]}
   );
   gpc1_1 gpc1136 (
      {stage1_49[13]},
      {stage2_49[7]}
   );
   gpc1_1 gpc1137 (
      {stage1_49[14]},
      {stage2_49[8]}
   );
   gpc1_1 gpc1138 (
      {stage1_49[15]},
      {stage2_49[9]}
   );
   gpc1_1 gpc1139 (
      {stage1_49[16]},
      {stage2_49[10]}
   );
   gpc1_1 gpc1140 (
      {stage1_49[17]},
      {stage2_49[11]}
   );
   gpc1_1 gpc1141 (
      {stage1_49[18]},
      {stage2_49[12]}
   );
   gpc1_1 gpc1142 (
      {stage1_49[19]},
      {stage2_49[13]}
   );
   gpc1_1 gpc1143 (
      {stage1_49[20]},
      {stage2_49[14]}
   );
   gpc1_1 gpc1144 (
      {stage1_49[21]},
      {stage2_49[15]}
   );
   gpc1_1 gpc1145 (
      {stage1_49[22]},
      {stage2_49[16]}
   );
   gpc1_1 gpc1146 (
      {stage1_49[23]},
      {stage2_49[17]}
   );
   gpc1_1 gpc1147 (
      {stage1_50[42]},
      {stage2_50[10]}
   );
   gpc1_1 gpc1148 (
      {stage1_51[46]},
      {stage2_51[15]}
   );
   gpc1_1 gpc1149 (
      {stage1_51[47]},
      {stage2_51[16]}
   );
   gpc1_1 gpc1150 (
      {stage1_52[17]},
      {stage2_52[14]}
   );
   gpc1_1 gpc1151 (
      {stage1_52[18]},
      {stage2_52[15]}
   );
   gpc1_1 gpc1152 (
      {stage1_52[19]},
      {stage2_52[16]}
   );
   gpc1_1 gpc1153 (
      {stage1_52[20]},
      {stage2_52[17]}
   );
   gpc1_1 gpc1154 (
      {stage1_52[21]},
      {stage2_52[18]}
   );
   gpc1_1 gpc1155 (
      {stage1_53[40]},
      {stage2_53[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_54[16]},
      {stage2_54[14]}
   );
   gpc1_1 gpc1157 (
      {stage1_55[32]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1158 (
      {stage1_55[33]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1159 (
      {stage1_55[34]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1160 (
      {stage1_55[35]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1161 (
      {stage1_55[36]},
      {stage2_55[17]}
   );
   gpc1_1 gpc1162 (
      {stage1_55[37]},
      {stage2_55[18]}
   );
   gpc1_1 gpc1163 (
      {stage1_56[17]},
      {stage2_56[9]}
   );
   gpc1_1 gpc1164 (
      {stage1_56[18]},
      {stage2_56[10]}
   );
   gpc1_1 gpc1165 (
      {stage1_56[19]},
      {stage2_56[11]}
   );
   gpc1_1 gpc1166 (
      {stage1_56[20]},
      {stage2_56[12]}
   );
   gpc1_1 gpc1167 (
      {stage1_57[37]},
      {stage2_57[9]}
   );
   gpc1_1 gpc1168 (
      {stage1_57[38]},
      {stage2_57[10]}
   );
   gpc1_1 gpc1169 (
      {stage1_57[39]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1170 (
      {stage1_57[40]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1171 (
      {stage1_58[6]},
      {stage2_58[9]}
   );
   gpc1_1 gpc1172 (
      {stage1_58[7]},
      {stage2_58[10]}
   );
   gpc1_1 gpc1173 (
      {stage1_58[8]},
      {stage2_58[11]}
   );
   gpc1_1 gpc1174 (
      {stage1_58[9]},
      {stage2_58[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_58[10]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_58[11]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_58[12]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1178 (
      {stage1_58[13]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1179 (
      {stage1_58[14]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1180 (
      {stage1_60[18]},
      {stage2_60[8]}
   );
   gpc1_1 gpc1181 (
      {stage1_60[19]},
      {stage2_60[9]}
   );
   gpc1_1 gpc1182 (
      {stage1_60[20]},
      {stage2_60[10]}
   );
   gpc1_1 gpc1183 (
      {stage1_60[21]},
      {stage2_60[11]}
   );
   gpc1_1 gpc1184 (
      {stage1_60[22]},
      {stage2_60[12]}
   );
   gpc1_1 gpc1185 (
      {stage1_61[18]},
      {stage2_61[9]}
   );
   gpc1_1 gpc1186 (
      {stage1_61[19]},
      {stage2_61[10]}
   );
   gpc1_1 gpc1187 (
      {stage1_61[20]},
      {stage2_61[11]}
   );
   gpc1_1 gpc1188 (
      {stage1_62[18]},
      {stage2_62[12]}
   );
   gpc1_1 gpc1189 (
      {stage1_62[19]},
      {stage2_62[13]}
   );
   gpc1_1 gpc1190 (
      {stage1_62[20]},
      {stage2_62[14]}
   );
   gpc1_1 gpc1191 (
      {stage1_62[21]},
      {stage2_62[15]}
   );
   gpc1_1 gpc1192 (
      {stage1_62[22]},
      {stage2_62[16]}
   );
   gpc1_1 gpc1193 (
      {stage1_62[23]},
      {stage2_62[17]}
   );
   gpc1_1 gpc1194 (
      {stage1_63[24]},
      {stage2_63[6]}
   );
   gpc1_1 gpc1195 (
      {stage1_63[25]},
      {stage2_63[7]}
   );
   gpc1_1 gpc1196 (
      {stage1_63[26]},
      {stage2_63[8]}
   );
   gpc1_1 gpc1197 (
      {stage1_63[27]},
      {stage2_63[9]}
   );
   gpc1_1 gpc1198 (
      {stage1_63[28]},
      {stage2_63[10]}
   );
   gpc1_1 gpc1199 (
      {stage1_63[29]},
      {stage2_63[11]}
   );
   gpc1_1 gpc1200 (
      {stage1_63[30]},
      {stage2_63[12]}
   );
   gpc1_1 gpc1201 (
      {stage1_63[31]},
      {stage2_63[13]}
   );
   gpc1_1 gpc1202 (
      {stage1_63[32]},
      {stage2_63[14]}
   );
   gpc1_1 gpc1203 (
      {stage1_63[33]},
      {stage2_63[15]}
   );
   gpc1_1 gpc1204 (
      {stage1_63[34]},
      {stage2_63[16]}
   );
   gpc1_1 gpc1205 (
      {stage1_65[2]},
      {stage2_65[6]}
   );
   gpc1_1 gpc1206 (
      {stage1_65[3]},
      {stage2_65[7]}
   );
   gpc1_1 gpc1207 (
      {stage1_65[4]},
      {stage2_65[8]}
   );
   gpc1_1 gpc1208 (
      {stage1_65[5]},
      {stage2_65[9]}
   );
   gpc615_5 gpc1209 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1210 (
      {stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc1211 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc1212 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3]}
   );
   gpc2135_5 gpc1213 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4]},
      {stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3]}
   );
   gpc615_5 gpc1214 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc1215 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[2]}
   );
   gpc606_5 gpc1216 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[3]}
   );
   gpc615_5 gpc1217 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2],stage3_12[3]}
   );
   gpc615_5 gpc1218 (
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage2_13[1]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[1],stage3_14[1],stage3_13[3],stage3_12[4]}
   );
   gpc623_5 gpc1219 (
      {stage2_13[2], stage2_13[3], stage2_13[4]},
      {stage2_14[12], stage2_14[13]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[2],stage3_15[2],stage3_14[2],stage3_13[4]}
   );
   gpc623_5 gpc1220 (
      {stage2_13[5], stage2_13[6], stage2_13[7]},
      {stage2_14[14], 1'b0},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[3],stage3_15[3],stage3_14[3],stage3_13[5]}
   );
   gpc135_4 gpc1221 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4]},
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[2],stage3_16[4]}
   );
   gpc606_5 gpc1222 (
      {stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[1],stage3_18[1],stage3_17[3],stage3_16[5]}
   );
   gpc606_5 gpc1223 (
      {stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[2],stage3_18[2],stage3_17[4]}
   );
   gpc1406_5 gpc1224 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[1],stage3_20[2],stage3_19[3],stage3_18[3]}
   );
   gpc1406_5 gpc1225 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[2],stage3_20[3],stage3_19[4],stage3_18[4]}
   );
   gpc615_5 gpc1226 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[3]}
   );
   gpc615_5 gpc1227 (
      {stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3],stage3_21[4]}
   );
   gpc615_5 gpc1228 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4],stage3_21[5]}
   );
   gpc1325_5 gpc1229 (
      {stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[3], stage2_22[4]},
      {stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage2_24[0]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5],stage3_21[6]}
   );
   gpc606_5 gpc1230 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6]},
      {stage3_26[0],stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[6]}
   );
   gpc1343_5 gpc1231 (
      {stage2_24[7], stage2_24[8], stage2_24[9]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3]},
      {stage2_26[0], stage2_26[1], stage2_26[2]},
      {stage2_27[0]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[5],stage3_24[5]}
   );
   gpc1325_5 gpc1232 (
      {stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_26[3], stage2_26[4]},
      {stage2_27[1], stage2_27[2], stage2_27[3]},
      {stage2_28[0]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[6]}
   );
   gpc1325_5 gpc1233 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], 1'b0},
      {stage2_26[5], stage2_26[6]},
      {stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage2_28[1]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[7]}
   );
   gpc606_5 gpc1234 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7]},
      {stage3_30[0],stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc606_5 gpc1235 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18]},
      {stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage3_30[1],stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc606_5 gpc1236 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[2],stage3_29[4]}
   );
   gpc606_5 gpc1237 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[1],stage3_31[1],stage3_30[3],stage3_29[5]}
   );
   gpc615_5 gpc1238 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[2],stage3_31[2],stage3_30[4]}
   );
   gpc615_5 gpc1239 (
      {stage2_30[5], stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[3],stage3_31[3],stage3_30[5]}
   );
   gpc606_5 gpc1240 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[0],stage3_35[0],stage3_34[2],stage3_33[4]}
   );
   gpc606_5 gpc1241 (
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[1],stage3_35[1],stage3_34[3]}
   );
   gpc606_5 gpc1242 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[2],stage3_35[2],stage3_34[4]}
   );
   gpc615_5 gpc1243 (
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[3],stage3_35[3]}
   );
   gpc615_5 gpc1244 (
      {stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage2_37[6]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4],stage3_36[4]}
   );
   gpc615_5 gpc1245 (
      {stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_38[6]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc615_5 gpc1246 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16]},
      {stage2_38[7]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[2],stage3_39[3],stage3_38[5],stage3_37[6]}
   );
   gpc207_4 gpc1247 (
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], 1'b0, 1'b0},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc615_5 gpc1248 (
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16]},
      {stage2_40[2]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[0],stage3_41[3],stage3_40[4],stage3_39[5]}
   );
   gpc606_5 gpc1249 (
      {stage2_40[3], stage2_40[4], stage2_40[5], stage2_40[6], stage2_40[7], stage2_40[8]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[1],stage3_42[1],stage3_41[4],stage3_40[5]}
   );
   gpc623_5 gpc1250 (
      {stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_41[6], stage2_41[7]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[2],stage3_42[2],stage3_41[5],stage3_40[6]}
   );
   gpc606_5 gpc1251 (
      {stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11], stage2_41[12], 1'b0},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[2],stage3_43[3],stage3_42[3],stage3_41[6]}
   );
   gpc606_5 gpc1252 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[0],stage3_46[0],stage3_45[1],stage3_44[3]}
   );
   gpc606_5 gpc1253 (
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[1],stage3_46[1],stage3_45[2],stage3_44[4]}
   );
   gpc606_5 gpc1254 (
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[2],stage3_46[2],stage3_45[3]}
   );
   gpc606_5 gpc1255 (
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[3],stage3_46[3],stage3_45[4]}
   );
   gpc615_5 gpc1256 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16]},
      {stage2_47[12]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[2],stage3_48[4],stage3_47[4],stage3_46[4]}
   );
   gpc606_5 gpc1257 (
      {stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17], stage2_47[18]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[1],stage3_49[3],stage3_48[5],stage3_47[5]}
   );
   gpc606_5 gpc1258 (
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[0],stage3_51[1],stage3_50[2],stage3_49[4]}
   );
   gpc606_5 gpc1259 (
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[1],stage3_51[2],stage3_50[3],stage3_49[5]}
   );
   gpc615_5 gpc1260 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4]},
      {stage2_51[12]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[2],stage3_52[2],stage3_51[3],stage3_50[4]}
   );
   gpc606_5 gpc1261 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[0],stage3_54[1],stage3_53[3],stage3_52[3]}
   );
   gpc606_5 gpc1262 (
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[1],stage3_55[1],stage3_54[2],stage3_53[4]}
   );
   gpc606_5 gpc1263 (
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[2],stage3_55[2],stage3_54[3],stage3_53[5]}
   );
   gpc135_4 gpc1264 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10]},
      {stage2_55[12], stage2_55[13], stage2_55[14]},
      {stage2_56[0]},
      {stage3_57[2],stage3_56[3],stage3_55[3],stage3_54[4]}
   );
   gpc135_4 gpc1265 (
      {stage2_54[11], stage2_54[12], stage2_54[13], stage2_54[14], 1'b0},
      {stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage2_56[1]},
      {stage3_57[3],stage3_56[4],stage3_55[4],stage3_54[5]}
   );
   gpc606_5 gpc1266 (
      {stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5], stage2_56[6], stage2_56[7]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[4],stage3_56[5]}
   );
   gpc135_4 gpc1267 (
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4]},
      {stage2_58[6], stage2_58[7], stage2_58[8]},
      {stage2_59[0]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[5]}
   );
   gpc135_4 gpc1268 (
      {stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9]},
      {stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage2_59[1]},
      {stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[6]}
   );
   gpc1163_5 gpc1269 (
      {stage2_57[10], stage2_57[11], stage2_57[12]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage2_59[2]},
      {stage2_60[0]},
      {stage3_61[0],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[7]}
   );
   gpc606_5 gpc1270 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[0],stage3_62[0],stage3_61[1],stage3_60[4]}
   );
   gpc606_5 gpc1271 (
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[1],stage3_62[1],stage3_61[2],stage3_60[5]}
   );
   gpc606_5 gpc1272 (
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[2],stage3_63[2],stage3_62[2],stage3_61[3]}
   );
   gpc606_5 gpc1273 (
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[3],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1274 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[4],stage3_63[4]}
   );
   gpc1_1 gpc1275 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1276 (
      {stage2_2[12]},
      {stage3_2[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_2[13]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc1279 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1280 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc1281 (
      {stage2_4[12]},
      {stage3_4[4]}
   );
   gpc1_1 gpc1282 (
      {stage2_4[13]},
      {stage3_4[5]}
   );
   gpc1_1 gpc1283 (
      {stage2_4[14]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1284 (
      {stage2_4[15]},
      {stage3_4[7]}
   );
   gpc1_1 gpc1285 (
      {stage2_4[16]},
      {stage3_4[8]}
   );
   gpc1_1 gpc1286 (
      {stage2_4[17]},
      {stage3_4[9]}
   );
   gpc1_1 gpc1287 (
      {stage2_4[18]},
      {stage3_4[10]}
   );
   gpc1_1 gpc1288 (
      {stage2_4[19]},
      {stage3_4[11]}
   );
   gpc1_1 gpc1289 (
      {stage2_4[20]},
      {stage3_4[12]}
   );
   gpc1_1 gpc1290 (
      {stage2_4[21]},
      {stage3_4[13]}
   );
   gpc1_1 gpc1291 (
      {stage2_4[22]},
      {stage3_4[14]}
   );
   gpc1_1 gpc1292 (
      {stage2_5[5]},
      {stage3_5[4]}
   );
   gpc1_1 gpc1293 (
      {stage2_5[6]},
      {stage3_5[5]}
   );
   gpc1_1 gpc1294 (
      {stage2_5[7]},
      {stage3_5[6]}
   );
   gpc1_1 gpc1295 (
      {stage2_5[8]},
      {stage3_5[7]}
   );
   gpc1_1 gpc1296 (
      {stage2_5[9]},
      {stage3_5[8]}
   );
   gpc1_1 gpc1297 (
      {stage2_6[9]},
      {stage3_6[3]}
   );
   gpc1_1 gpc1298 (
      {stage2_6[10]},
      {stage3_6[4]}
   );
   gpc1_1 gpc1299 (
      {stage2_7[1]},
      {stage3_7[2]}
   );
   gpc1_1 gpc1300 (
      {stage2_7[2]},
      {stage3_7[3]}
   );
   gpc1_1 gpc1301 (
      {stage2_7[3]},
      {stage3_7[4]}
   );
   gpc1_1 gpc1302 (
      {stage2_7[4]},
      {stage3_7[5]}
   );
   gpc1_1 gpc1303 (
      {stage2_7[5]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1304 (
      {stage2_7[6]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1305 (
      {stage2_7[7]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1306 (
      {stage2_7[8]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1307 (
      {stage2_7[9]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[10]},
      {stage3_7[11]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[11]},
      {stage3_7[12]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[12]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1311 (
      {stage2_8[7]},
      {stage3_8[3]}
   );
   gpc1_1 gpc1312 (
      {stage2_8[8]},
      {stage3_8[4]}
   );
   gpc1_1 gpc1313 (
      {stage2_8[9]},
      {stage3_8[5]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[10]},
      {stage3_8[6]}
   );
   gpc1_1 gpc1315 (
      {stage2_9[13]},
      {stage3_9[4]}
   );
   gpc1_1 gpc1316 (
      {stage2_9[14]},
      {stage3_9[5]}
   );
   gpc1_1 gpc1317 (
      {stage2_9[15]},
      {stage3_9[6]}
   );
   gpc1_1 gpc1318 (
      {stage2_9[16]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1319 (
      {stage2_9[17]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1320 (
      {stage2_9[18]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[19]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1322 (
      {stage2_10[6]},
      {stage3_10[3]}
   );
   gpc1_1 gpc1323 (
      {stage2_10[7]},
      {stage3_10[4]}
   );
   gpc1_1 gpc1324 (
      {stage2_10[8]},
      {stage3_10[5]}
   );
   gpc1_1 gpc1325 (
      {stage2_10[9]},
      {stage3_10[6]}
   );
   gpc1_1 gpc1326 (
      {stage2_11[12]},
      {stage3_11[3]}
   );
   gpc1_1 gpc1327 (
      {stage2_13[8]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1328 (
      {stage2_13[9]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1329 (
      {stage2_15[12]},
      {stage3_15[4]}
   );
   gpc1_1 gpc1330 (
      {stage2_15[13]},
      {stage3_15[5]}
   );
   gpc1_1 gpc1331 (
      {stage2_17[9]},
      {stage3_17[5]}
   );
   gpc1_1 gpc1332 (
      {stage2_17[10]},
      {stage3_17[6]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[11]},
      {stage3_17[7]}
   );
   gpc1_1 gpc1334 (
      {stage2_18[19]},
      {stage3_18[5]}
   );
   gpc1_1 gpc1335 (
      {stage2_19[6]},
      {stage3_19[5]}
   );
   gpc1_1 gpc1336 (
      {stage2_19[7]},
      {stage3_19[6]}
   );
   gpc1_1 gpc1337 (
      {stage2_19[8]},
      {stage3_19[7]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[8]},
      {stage3_20[4]}
   );
   gpc1_1 gpc1339 (
      {stage2_29[12]},
      {stage3_29[6]}
   );
   gpc1_1 gpc1340 (
      {stage2_29[13]},
      {stage3_29[7]}
   );
   gpc1_1 gpc1341 (
      {stage2_29[14]},
      {stage3_29[8]}
   );
   gpc1_1 gpc1342 (
      {stage2_29[15]},
      {stage3_29[9]}
   );
   gpc1_1 gpc1343 (
      {stage2_29[16]},
      {stage3_29[10]}
   );
   gpc1_1 gpc1344 (
      {stage2_29[17]},
      {stage3_29[11]}
   );
   gpc1_1 gpc1345 (
      {stage2_31[14]},
      {stage3_31[4]}
   );
   gpc1_1 gpc1346 (
      {stage2_31[15]},
      {stage3_31[5]}
   );
   gpc1_1 gpc1347 (
      {stage2_31[16]},
      {stage3_31[6]}
   );
   gpc1_1 gpc1348 (
      {stage2_33[6]},
      {stage3_33[5]}
   );
   gpc1_1 gpc1349 (
      {stage2_33[7]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1350 (
      {stage2_33[8]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1351 (
      {stage2_33[9]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1352 (
      {stage2_33[10]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1353 (
      {stage2_33[11]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1354 (
      {stage2_33[12]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1355 (
      {stage2_33[13]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1356 (
      {stage2_33[14]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1357 (
      {stage2_33[15]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1358 (
      {stage2_34[12]},
      {stage3_34[5]}
   );
   gpc1_1 gpc1359 (
      {stage2_34[13]},
      {stage3_34[6]}
   );
   gpc1_1 gpc1360 (
      {stage2_34[14]},
      {stage3_34[7]}
   );
   gpc1_1 gpc1361 (
      {stage2_34[15]},
      {stage3_34[8]}
   );
   gpc1_1 gpc1362 (
      {stage2_36[18]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1363 (
      {stage2_42[12]},
      {stage3_42[4]}
   );
   gpc1_1 gpc1364 (
      {stage2_42[13]},
      {stage3_42[5]}
   );
   gpc1_1 gpc1365 (
      {stage2_43[6]},
      {stage3_43[4]}
   );
   gpc1_1 gpc1366 (
      {stage2_43[7]},
      {stage3_43[5]}
   );
   gpc1_1 gpc1367 (
      {stage2_43[8]},
      {stage3_43[6]}
   );
   gpc1_1 gpc1368 (
      {stage2_43[9]},
      {stage3_43[7]}
   );
   gpc1_1 gpc1369 (
      {stage2_44[12]},
      {stage3_44[5]}
   );
   gpc1_1 gpc1370 (
      {stage2_44[13]},
      {stage3_44[6]}
   );
   gpc1_1 gpc1371 (
      {stage2_44[14]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1372 (
      {stage2_46[17]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1373 (
      {stage2_47[19]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1374 (
      {stage2_47[20]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1375 (
      {stage2_47[21]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1376 (
      {stage2_48[6]},
      {stage3_48[6]}
   );
   gpc1_1 gpc1377 (
      {stage2_48[7]},
      {stage3_48[7]}
   );
   gpc1_1 gpc1378 (
      {stage2_48[8]},
      {stage3_48[8]}
   );
   gpc1_1 gpc1379 (
      {stage2_48[9]},
      {stage3_48[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_48[10]},
      {stage3_48[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_48[11]},
      {stage3_48[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_48[12]},
      {stage3_48[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_50[5]},
      {stage3_50[5]}
   );
   gpc1_1 gpc1384 (
      {stage2_50[6]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1385 (
      {stage2_50[7]},
      {stage3_50[7]}
   );
   gpc1_1 gpc1386 (
      {stage2_50[8]},
      {stage3_50[8]}
   );
   gpc1_1 gpc1387 (
      {stage2_50[9]},
      {stage3_50[9]}
   );
   gpc1_1 gpc1388 (
      {stage2_50[10]},
      {stage3_50[10]}
   );
   gpc1_1 gpc1389 (
      {stage2_51[13]},
      {stage3_51[4]}
   );
   gpc1_1 gpc1390 (
      {stage2_51[14]},
      {stage3_51[5]}
   );
   gpc1_1 gpc1391 (
      {stage2_51[15]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1392 (
      {stage2_51[16]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1393 (
      {stage2_52[12]},
      {stage3_52[4]}
   );
   gpc1_1 gpc1394 (
      {stage2_52[13]},
      {stage3_52[5]}
   );
   gpc1_1 gpc1395 (
      {stage2_52[14]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1396 (
      {stage2_52[15]},
      {stage3_52[7]}
   );
   gpc1_1 gpc1397 (
      {stage2_52[16]},
      {stage3_52[8]}
   );
   gpc1_1 gpc1398 (
      {stage2_52[17]},
      {stage3_52[9]}
   );
   gpc1_1 gpc1399 (
      {stage2_52[18]},
      {stage3_52[10]}
   );
   gpc1_1 gpc1400 (
      {stage2_53[12]},
      {stage3_53[6]}
   );
   gpc1_1 gpc1401 (
      {stage2_55[18]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1402 (
      {stage2_56[8]},
      {stage3_56[6]}
   );
   gpc1_1 gpc1403 (
      {stage2_56[9]},
      {stage3_56[7]}
   );
   gpc1_1 gpc1404 (
      {stage2_56[10]},
      {stage3_56[8]}
   );
   gpc1_1 gpc1405 (
      {stage2_56[11]},
      {stage3_56[9]}
   );
   gpc1_1 gpc1406 (
      {stage2_56[12]},
      {stage3_56[10]}
   );
   gpc1_1 gpc1407 (
      {stage2_59[3]},
      {stage3_59[4]}
   );
   gpc1_1 gpc1408 (
      {stage2_59[4]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1409 (
      {stage2_59[5]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1410 (
      {stage2_59[6]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1411 (
      {stage2_59[7]},
      {stage3_59[8]}
   );
   gpc1_1 gpc1412 (
      {stage2_59[8]},
      {stage3_59[9]}
   );
   gpc1_1 gpc1413 (
      {stage2_59[9]},
      {stage3_59[10]}
   );
   gpc1_1 gpc1414 (
      {stage2_59[10]},
      {stage3_59[11]}
   );
   gpc1_1 gpc1415 (
      {stage2_59[11]},
      {stage3_59[12]}
   );
   gpc1_1 gpc1416 (
      {stage2_59[12]},
      {stage3_59[13]}
   );
   gpc1_1 gpc1417 (
      {stage2_61[6]},
      {stage3_61[4]}
   );
   gpc1_1 gpc1418 (
      {stage2_61[7]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1419 (
      {stage2_61[8]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1420 (
      {stage2_61[9]},
      {stage3_61[7]}
   );
   gpc1_1 gpc1421 (
      {stage2_61[10]},
      {stage3_61[8]}
   );
   gpc1_1 gpc1422 (
      {stage2_61[11]},
      {stage3_61[9]}
   );
   gpc1_1 gpc1423 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1424 (
      {stage2_63[13]},
      {stage3_63[6]}
   );
   gpc1_1 gpc1425 (
      {stage2_63[14]},
      {stage3_63[7]}
   );
   gpc1_1 gpc1426 (
      {stage2_63[15]},
      {stage3_63[8]}
   );
   gpc1_1 gpc1427 (
      {stage2_63[16]},
      {stage3_63[9]}
   );
   gpc1_1 gpc1428 (
      {stage2_65[6]},
      {stage3_65[3]}
   );
   gpc1_1 gpc1429 (
      {stage2_65[7]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1430 (
      {stage2_65[8]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1431 (
      {stage2_65[9]},
      {stage3_65[6]}
   );
   gpc1_1 gpc1432 (
      {stage2_66[0]},
      {stage3_66[2]}
   );
   gpc1_1 gpc1433 (
      {stage2_66[1]},
      {stage3_66[3]}
   );
   gpc1_1 gpc1434 (
      {stage2_66[2]},
      {stage3_66[4]}
   );
   gpc1_1 gpc1435 (
      {stage2_66[3]},
      {stage3_66[5]}
   );
   gpc615_5 gpc1436 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc1437 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1]}
   );
   gpc2135_5 gpc1438 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[2]}
   );
   gpc615_5 gpc1439 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], 1'b0},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[3]}
   );
   gpc615_5 gpc1440 (
      {stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1441 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12]},
      {1'b0},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], 1'b0},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc7_3 gpc1442 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1443 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], 1'b0},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[3]}
   );
   gpc207_4 gpc1444 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1]}
   );
   gpc1415_5 gpc1445 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], 1'b0},
      {stage3_15[2]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[2]}
   );
   gpc117_4 gpc1446 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1]}
   );
   gpc1406_5 gpc1447 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc615_5 gpc1448 (
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[4]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1],stage4_20[2]}
   );
   gpc615_5 gpc1449 (
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[2]}
   );
   gpc15_3 gpc1450 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[6]},
      {stage4_26[1],stage4_25[1],stage4_24[2]}
   );
   gpc615_5 gpc1451 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4]},
      {stage3_27[0]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], 1'b0},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[2]}
   );
   gpc1163_5 gpc1452 (
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[1]}
   );
   gpc606_5 gpc1453 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage4_33[1],stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[2]}
   );
   gpc3_2 gpc1454 (
      {stage3_32[1], stage3_32[2], stage3_32[3]},
      {stage4_33[2],stage4_32[2]}
   );
   gpc2135_5 gpc1455 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[3]}
   );
   gpc2135_5 gpc1456 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[1],stage4_33[4]}
   );
   gpc2135_5 gpc1457 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_34[6], stage3_34[7], stage3_34[8]},
      {stage3_35[2]},
      {stage3_36[4], stage3_36[5]},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[2],stage4_33[5]}
   );
   gpc615_5 gpc1458 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4]},
      {stage3_38[0]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3]}
   );
   gpc2116_5 gpc1459 (
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage3_41[0]},
      {stage3_42[0]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1],stage4_40[1]}
   );
   gpc207_4 gpc1460 (
      {stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], 1'b0},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[1],stage4_41[2]}
   );
   gpc2135_5 gpc1461 (
      {stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage3_43[4], stage3_43[5], stage3_43[6]},
      {stage3_44[0]},
      {stage3_45[0], stage3_45[1]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[2]}
   );
   gpc2135_5 gpc1462 (
      {stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage3_45[2], stage3_45[3], stage3_45[4]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc615_5 gpc1463 (
      {stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[2]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[2]}
   );
   gpc615_5 gpc1464 (
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7]},
      {stage3_48[6]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[2],stage4_47[2]}
   );
   gpc606_5 gpc1465 (
      {stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11], stage3_48[12]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[1],stage4_50[2],stage4_49[2],stage4_48[3]}
   );
   gpc615_5 gpc1466 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[1],stage4_51[2],stage4_50[3]}
   );
   gpc606_5 gpc1467 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5], stage3_51[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[2],stage4_51[3]}
   );
   gpc615_5 gpc1468 (
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[2],stage4_53[2],stage4_52[3]}
   );
   gpc1343_5 gpc1469 (
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3]},
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2]}
   );
   gpc1343_5 gpc1470 (
      {stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_56[4], stage3_56[5], stage3_56[6], stage3_56[7]},
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[1]},
      {stage4_59[1],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc623_5 gpc1471 (
      {stage3_57[6], stage3_57[7], 1'b0},
      {stage3_58[2], stage3_58[3]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[2],stage4_58[2],stage4_57[2]}
   );
   gpc606_5 gpc1472 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[1],stage4_59[3]}
   );
   gpc117_4 gpc1473 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5], 1'b0},
      {stage3_61[6]},
      {stage3_62[0]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc2223_5 gpc1474 (
      {stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0], stage3_63[1]},
      {stage3_64[0], stage3_64[1]},
      {stage3_65[0], stage3_65[1]},
      {stage4_66[0],stage4_65[0],stage4_64[0],stage4_63[2],stage4_62[2]}
   );
   gpc606_5 gpc1475 (
      {stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6], stage3_63[7]},
      {stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5], stage3_65[6], 1'b0},
      {stage4_67[0],stage4_66[1],stage4_65[1],stage4_64[1],stage4_63[3]}
   );
   gpc606_5 gpc1476 (
      {stage3_64[2], stage3_64[3], stage3_64[4], 1'b0, 1'b0, 1'b0},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[2],stage4_65[2],stage4_64[2]}
   );
   gpc1_1 gpc1477 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1478 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1479 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc1480 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1481 (
      {stage3_4[12]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1482 (
      {stage3_4[13]},
      {stage4_4[4]}
   );
   gpc1_1 gpc1483 (
      {stage3_4[14]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1484 (
      {stage3_7[13]},
      {stage4_7[5]}
   );
   gpc1_1 gpc1485 (
      {stage3_12[3]},
      {stage4_12[2]}
   );
   gpc1_1 gpc1486 (
      {stage3_12[4]},
      {stage4_12[3]}
   );
   gpc1_1 gpc1487 (
      {stage3_15[3]},
      {stage4_15[2]}
   );
   gpc1_1 gpc1488 (
      {stage3_15[4]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1489 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc1490 (
      {stage3_16[4]},
      {stage4_16[2]}
   );
   gpc1_1 gpc1491 (
      {stage3_16[5]},
      {stage4_16[3]}
   );
   gpc1_1 gpc1492 (
      {stage3_18[1]},
      {stage4_18[2]}
   );
   gpc1_1 gpc1493 (
      {stage3_18[2]},
      {stage4_18[3]}
   );
   gpc1_1 gpc1494 (
      {stage3_18[3]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1495 (
      {stage3_18[4]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1496 (
      {stage3_18[5]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1497 (
      {stage3_19[7]},
      {stage4_19[2]}
   );
   gpc1_1 gpc1498 (
      {stage3_21[5]},
      {stage4_21[2]}
   );
   gpc1_1 gpc1499 (
      {stage3_21[6]},
      {stage4_21[3]}
   );
   gpc1_1 gpc1500 (
      {stage3_25[7]},
      {stage4_25[2]}
   );
   gpc1_1 gpc1501 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1502 (
      {stage3_27[1]},
      {stage4_27[2]}
   );
   gpc1_1 gpc1503 (
      {stage3_27[2]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1504 (
      {stage3_27[3]},
      {stage4_27[4]}
   );
   gpc1_1 gpc1505 (
      {stage3_27[4]},
      {stage4_27[5]}
   );
   gpc1_1 gpc1506 (
      {stage3_29[9]},
      {stage4_29[3]}
   );
   gpc1_1 gpc1507 (
      {stage3_29[10]},
      {stage4_29[4]}
   );
   gpc1_1 gpc1508 (
      {stage3_29[11]},
      {stage4_29[5]}
   );
   gpc1_1 gpc1509 (
      {stage3_35[3]},
      {stage4_35[3]}
   );
   gpc1_1 gpc1510 (
      {stage3_37[5]},
      {stage4_37[4]}
   );
   gpc1_1 gpc1511 (
      {stage3_37[6]},
      {stage4_37[5]}
   );
   gpc1_1 gpc1512 (
      {stage3_38[1]},
      {stage4_38[1]}
   );
   gpc1_1 gpc1513 (
      {stage3_38[2]},
      {stage4_38[2]}
   );
   gpc1_1 gpc1514 (
      {stage3_38[3]},
      {stage4_38[3]}
   );
   gpc1_1 gpc1515 (
      {stage3_38[4]},
      {stage4_38[4]}
   );
   gpc1_1 gpc1516 (
      {stage3_38[5]},
      {stage4_38[5]}
   );
   gpc1_1 gpc1517 (
      {stage3_38[6]},
      {stage4_38[6]}
   );
   gpc1_1 gpc1518 (
      {stage3_40[6]},
      {stage4_40[2]}
   );
   gpc1_1 gpc1519 (
      {stage3_43[7]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1520 (
      {stage3_44[6]},
      {stage4_44[4]}
   );
   gpc1_1 gpc1521 (
      {stage3_44[7]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1522 (
      {stage3_47[8]},
      {stage4_47[3]}
   );
   gpc1_1 gpc1523 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1524 (
      {stage3_56[8]},
      {stage4_56[3]}
   );
   gpc1_1 gpc1525 (
      {stage3_56[9]},
      {stage4_56[4]}
   );
   gpc1_1 gpc1526 (
      {stage3_56[10]},
      {stage4_56[5]}
   );
   gpc1_1 gpc1527 (
      {stage3_59[12]},
      {stage4_59[4]}
   );
   gpc1_1 gpc1528 (
      {stage3_59[13]},
      {stage4_59[5]}
   );
   gpc1_1 gpc1529 (
      {stage3_61[7]},
      {stage4_61[3]}
   );
   gpc1_1 gpc1530 (
      {stage3_61[8]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1531 (
      {stage3_61[9]},
      {stage4_61[5]}
   );
   gpc1_1 gpc1532 (
      {stage3_63[8]},
      {stage4_63[4]}
   );
   gpc1_1 gpc1533 (
      {stage3_63[9]},
      {stage4_63[5]}
   );
   gpc1_1 gpc1534 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc207_4 gpc1535 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], 1'b0},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0]}
   );
   gpc623_5 gpc1536 (
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[2], stage4_6[3]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc135_4 gpc1537 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], 1'b0},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc1343_5 gpc1538 (
      {stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1343_5 gpc1539 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1]}
   );
   gpc7_3 gpc1540 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1343_5 gpc1541 (
      {stage4_19[0], stage4_19[1], stage4_19[2]},
      {stage4_20[0], stage4_20[1], stage4_20[2], 1'b0},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc23_3 gpc1542 (
      {stage4_23[0], stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[0],stage5_23[1]}
   );
   gpc1343_5 gpc1543 (
      {stage4_24[2], 1'b0, 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2], 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc615_5 gpc1544 (
      {stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[1]}
   );
   gpc223_4 gpc1545 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0], stage4_31[1]},
      {stage4_32[0], stage4_32[1]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[1]}
   );
   gpc606_5 gpc1546 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], 1'b0, 1'b0},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[0],stage5_33[1]}
   );
   gpc3_2 gpc1547 (
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage5_35[1],stage5_34[1]}
   );
   gpc1163_5 gpc1548 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc606_5 gpc1549 (
      {stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0, 1'b0, 1'b0},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1550 (
      {stage4_41[0], stage4_41[1], stage4_41[2]},
      {stage4_42[0], stage4_42[1], stage4_42[2], 1'b0},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1551 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], 1'b0},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1552 (
      {stage4_46[1], stage4_46[2], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1343_5 gpc1553 (
      {stage4_49[1], stage4_49[2], 1'b0},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3]},
      {stage4_51[0], stage4_51[1], stage4_51[2]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc1343_5 gpc1554 (
      {stage4_51[3], stage4_51[4], 1'b0},
      {stage4_52[1], stage4_52[2], stage4_52[3], 1'b0},
      {stage4_53[0], stage4_53[1], stage4_53[2]},
      {stage4_54[0]},
      {stage5_55[0],stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc1343_5 gpc1555 (
      {stage4_54[1], stage4_54[2], 1'b0},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3]},
      {stage4_56[0], stage4_56[1], stage4_56[2]},
      {stage4_57[0]},
      {stage5_58[0],stage5_57[0],stage5_56[0],stage5_55[1],stage5_54[1]}
   );
   gpc1343_5 gpc1556 (
      {stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage4_57[1], stage4_57[2], 1'b0, 1'b0},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[1],stage5_56[1]}
   );
   gpc135_4 gpc1557 (
      {stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[0], stage4_60[1], stage4_60[2]},
      {stage4_61[0]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1]}
   );
   gpc2135_5 gpc1558 (
      {stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc615_5 gpc1559 (
      {stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_64[2]},
      {stage4_65[0], stage4_65[1], stage4_65[2], 1'b0, 1'b0, 1'b0},
      {stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1],stage5_63[1]}
   );
   gpc2135_5 gpc1560 (
      {stage4_66[0], stage4_66[1], stage4_66[2], 1'b0, 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2]},
      {stage4_68[0]},
      {1'b0, 1'b0},
      {stage5_69[0],stage5_68[0],stage5_67[1],stage5_66[1]}
   );
   gpc1_1 gpc1561 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1562 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1563 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1564 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1565 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc1566 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc1567 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc1568 (
      {stage4_12[3]},
      {stage5_12[1]}
   );
   gpc1_1 gpc1569 (
      {stage4_13[1]},
      {stage5_13[1]}
   );
   gpc1_1 gpc1570 (
      {stage4_15[4]},
      {stage5_15[1]}
   );
   gpc1_1 gpc1571 (
      {stage4_16[3]},
      {stage5_16[1]}
   );
   gpc1_1 gpc1572 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc1573 (
      {stage4_21[3]},
      {stage5_21[1]}
   );
   gpc1_1 gpc1574 (
      {stage4_22[1]},
      {stage5_22[1]}
   );
   gpc1_1 gpc1575 (
      {stage4_26[3]},
      {stage5_26[1]}
   );
   gpc1_1 gpc1576 (
      {stage4_32[2]},
      {stage5_32[1]}
   );
   gpc1_1 gpc1577 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1578 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor_CLA54_64 compressor_CLA54_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf557993b258c583d6b470edca4cdc9e7a9eea5e8eecc9fb6f666c123854fb126fd1e05f7914f22046a285bea887fe84ff3ba30c0c9349787c2b60401c400af6ad16ec82e200d336813510dda5a77c55e3c460e498fabc7e91b60c3ded2477018594a212724a11f79716495f332596342b063e6eb6ae2248ba1e962146a63539b498eb44d71d3bd19ef3860224e9fffd2d12a44c55913b4b3c4702a1e0d09c9897a154f3c2594136d79be8b48a82612d8dc5f56e7ee710b90a40e888a52cc2d50d264989177adc5151838e24fbb6b5528c5cc56c676c9458cc6ce8b1bebc1e09b157941a2a00900d8173a7642ce836aef2c218489f91a11f09d592b84fdec73759c39f98ede0bac27e4b8cd1c4cfedaf02e1b96530ba9c3e3f15a2f71598088ff2bdeece631cb49f72f23da10659e6ca9b1b375b4ce2a0c4840335909a60cfdb654fb7c67b7b92e75172b4e21c675b45f272641e3ae63e813f2f868247227a5a34cdad9964a71a86c214b374b4283d6548a875f7568e4353cf3b0f740663f344a9c31e533acb15f3f8fdbf671146b97b0b0a9999b7323a92bf8d6d15e22b13f12f84c0e0c53889ab45398aa34f4ce27c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcd7fc3a15d2e5bea10e2bf273f0e65b6c0ccce895593738b1812cbbe594d1e23027d1531959eaf8e0b55ccd861225feaeae873cbb9e63cf730b9902db335a687ad816a71cdafa9c8343a390725ece7fd38f9aaa32a37a59b0de79aa3d59bd68645f81637489892135cfa67b3d65b299d024112b2e3c0450c5d0ecee43440099b90122ecd9dfeb2b0a20916c145b32096374db3e8fc7c91522bc7da861f9a522ea1d0b808f4f289dc664164eae42fc4c11b0f73c6be30d828fd495609a55a06588a52a48e2481d797d8618ab64248c856122c3b378c7e22cbb3c347bd306662a73f12c48ebc2b496b843c5c823998df0b00d9de7eb316e6d9e395ceb4fabb2c1de05c48da2506b524c61c664f982c9e1d7ea405c73cd0cb9dc63251450efc16bb1ab48110d49bbf5d19dd07b07a0f5669c3c4b8fb4b6128864a7e545bc324fd12efeb9c89ffcccbb04dac15644dd2df413eb60dfa419f99f93ecd02647f39044d5e23c94f7c2ee78194a1c349abb58e2e6e8f248fa5ceb5df07ad17593c500525f3a5e3e5359063b26cfbeb97908a0463695442cd603a01465f41c15dbefaa1b951ec1a3ac4d0dc8259a31b68f4a8f07c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf2b0286714e08e8abd18423c3da17173c33428744aba48bdfaf6034999923f890a37cc3e46ba954375312b62d9030366457c4c089a1101e42c6e3e294193aa0cb94d65fd86e3e4114c74d64411a4ac8c234de4cfaa92038e1733e2ec338306093967cd8f87c8ff311979357b345229c561ee4acbbcf60b005ffa8f161079c3d899b940d45997bc62452dbc1734911d98c5d643a63ce4f1d10c82f6fdc84641bcf2b4df423376eb922deacead5e87dcef7025cffbf58e8350ac77c8e0eab828013c620e9bd11bbb999fc1d2e42f14d1a749a36a623d4bba679edc2cefb884da943eb16cd75f1c1f2d59f69918814aba498513d0ae58f8b81bc4eba7eb29253aa01f092d0953dcc19c2c435c1d50c477a27d069e4ec52c2101c2c4e4471a129da893545df637d2cd0f30db4825d5355beff4043ade668f257bf990c3394dcd4dc94f1128e3e6294f4b2735bfe5bbdc9db960672bb6b187ad4d8907c67d2d91d975be08b16a88748f8d45d32fc03b6b8e2723829d2427544612916ef62f1f70b45a48c832456628f04214ca07d214ece0d2907eedacd060d62589905e8f4dd07578d828dbc37ce464ed18fb1c0f9f7a1656;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdeaa7d8101ed341e5c02c3a913f5bf666d6b258a507195ef1672bc067cd4ccb7ecc789a78bbd536a158ca57e3e910d29d8c3a9bcb21eee326457370f6a0102b1561f9c633a576cee8b26ad9911fe4054705ddd232c370aeef7d6c7730b0c90775ddbb2df1d5d6bf86d344e13eeaae5a713d60c5f204fdf759987c6db44eed8b0636f17b7e130746578f358f1ca30500ddaac43079b38346f2822366aa03b546c67269d86081bf4a80188bc5d9edd25762c139b320d422e54a6cf93a605c53284a4a2ee0ce9a67bbc976c71ca31469754426ba470d511b355833aca628cb3081a651da6c13f0d9efedf2d194488a4a2c68d2d0a6c4a239ff2b0cf6545518ff3a0a7218a8a09d840df743263ad2549a68eefea0482473b7988ede654984636a21c8ca02a01bcf3eb6c176ae2baf79394ab031d6b69219e7fcdf5cae1480f0310f83811a5783b50e7c291da347e9a7c1fbf6b9bb223d3710a49b53772206a470e957baac56376b7dafb00200110331ea30542a8f5a48a9d1a481ecdb124fa672baf1c9a895a2a98735366673390956af5d17265274f276c2fd01e7a5e5766314ac4d0466b01960db02071d2c10c81066e60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc75a4bbd1c93f1ad304afaccebef0e57e9a42bc8b747dea58c443e7e687d1a6da269b5ff37559a8454e0266760ee3e8e3bfe680f9f79d52f9ecb5badb602fe0aa6c8e46e08d56f28589be5d082c82cfca69ac7b0d97e2918be0fce11c27a63acdb1d8912e9959be7bea1bec4ee6ed394fc4459a10a2f462de844dd289adec435df33fb11abd3bbe6be426aec6a768c62f1a77a15c0e189197b1ed8ecf74d949346f7fab792599d93d3eafd7dc225b6c8f0d0e2d7b4e92d738b705b2764beaabcc80a214d2f8fec8611eefad55cd4d9a11ad41f2cc911beb27487dd0ae962030019fca7d81dce0684563b99504ceddf07fb6384d9e427e1b586814cf1e1c42d4f5349c3304f9beb588770973b52d416b7e697983ea69763b8553e815b688d7eca5efe2bd8ff2d886db677036650f9e04b4ca0734280f3861ecc6d420513ddac0a16df7438da19f5bd67b1d079c678e07f9dbf48aad1e478a4a551336ab3389977aaefa4abb4196b9c246bf7ba99572b8d2a821ffa8f769a260272234ee4aaa0c2b7984dae98a3a06099589d4e4afdc3ec9966506260b0024c488dd6c3f0ba4f21d80e8d6c97712b939ecd1d35eb1156bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h58aebd6e9175ee37469d39c67442d38d0eef9c6acbcd90afb21aaa5a4eac01e31249be3495697a1da8b83048a0bccb8fa94c68be38bc3473f900aa96254e67445523a9428607cdab03793638972e90ed448106fbeed199a46497442b3249f08950d9d3663879bbe9405bccaa1f835ce0a9c7926ce2230dd90eb196a5063167a5bf98d84c65ed97155d2e22daf84e47c3e6b0fd19d6c6af1d3ef06fe2eefce23da8219e8cdb490ded160205b88c19618be9ac2b941275635e2e8f6baa14d7a08e95c09bcf842e191fd50fe00256268a836ebad6b762868aa33d4657702f0d9fbd03ececdb3726f8177097c78fa30bb68c815c05983c1b21fee9af76d24eae0efb85a7e69084aed57de4b200a852314707120615b1d48de315f28375e7e8aed412b3957541024ce7b4a79bee73734037712bd30cfd1e941522220321006f710044dc26ae31f94b21b24232a1f1d9b2ff87b5e31908b2824c076be5d4b3128f0f6aec3e665d57cc1e110526c6a95216866dbc83b63e6cfb11454dda485f6e37df390ead3a1b71b6314994bacae3b2d4bef5f47c6f91fbc25d6e0f3706bb488228a395c1b25408d8050cb68a0be978bb9b83;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha8f187d2255f1ddbe021eafa3e832d9344a9391b339575ef218e3d2d9c1e05ea5a63c9b1768db6907d43892baa05e9b52bc5cc4895e7a3f2d2afe1edc922b6229d430a78314a7602a868ded4b2e08df071ec69208bc628223f15fda99cc08ddefd5d4e0b46a6be18a4115d4d20fc9bab95660e5f9615db17a066b2aecd994858160082636c94f4f904bb4cdacd97850c3caea72ac361b226215653213a50a1bceb0adce47112ead7c5a8154f6e74671bc81902e448462a5f80f81ff4e10740434b4668571be5d353e9ef4d8bed61ada019f286d1fb278ee0dead3bb2f3fa6265d661eff1093dcfd8560bd6533ad030bf69852388a2b311f086666093c1a3d092b7365f8f2a21fe5cc14aab94a6319acb06543bdf2ba68bb8ede86498e27a53ff236db4cd76cbf97cb0d443a3cae0dabd8a5b266841e5bc39ed84a8d4aafaba6e88451ede233c2c48be4724a4d19e340437affef96ce26a6c0f951c079c171f260b03cd16850ae6ec6d401d4a52ad925b8e980e8ab7c984ab436befe6046da96f04555ccbf526fa32c4df093bae6ae5e0bc00fc64dfa5c3ab208457a9391f1e87eb3e8792727ff30c7b5be979eb70ff8d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdb4e5db1e8ec39447ae30583058378e860f54ea833dba34f5c39ddbc51652851e994107a0a8adaf3be15cd8066e8e6ffd11328f9f01c967433d16bbf778e5d7bd0bf8b6c17d99f73fdbc8dcbe65a8c522afe71cf504c344127c694bf13803efd5965e3478b78e5e6b0b27cef707842b783142ca63eb704182152d0a909dcfd466fd4c5eae396dbf8ac8c739078d4f20b2ad5d951d88d5acac2d5a4830f08a71770231e8d18be395e3082e3c2d9ff04521b5d45ef748a24641eceeb841fd77e454d2555e07a904da36ef3965480953380f40e2bd99d1eef46fa74a004ac42f2e7dfc543ccf85d70881c7dd70f6dafe602ae7ec92977873a833df43936b517874d051de8eab8b221b67c0c0f5b3bbae8f9a598bc642c850ff53aaf7c249b8880f166f2682f6f44557ab476edb27433f5993c802243cd23dd5874f0803afe3cebc9a6c949f65f2112e862a5ef16875d5c4e5eaa2228e7d80f59564807f0a88e13f3002bbeccabd496d34799ad356cd3b84e8c581075634b33e7200af6118c63a4d9d343483b26f396d675cab218e04415c567fce30913c8195180233e91400a749e4b5859dda576a306d2038f36641d78f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8c1b524316f06b193544577054993a54a33a36de3ba9e1e2019a8b1e6ab3f4cbfdfd6172b7a1ea2f4c3b3b321fa440662288381ed970ffb535016ea783aa270f464f117da7020edf4c6f5a2914fed32235ba963abac0af567ac2fd84e4f93890c467a8138ffc0ebcc7db28eebf12c4ae3b822a8225f1f3a98f159575e8fac6aad45a19e528e0522952d95cc2204794b2f5c1d317c0026cfd94100b6f044223c1613fa297e9ca62c349449838811bce53bce6d7c890923b4b889ac3b5280887e65e77f5f337d0a1c76dfdcf0e9aca675bbd83d23cfb833084d02fe6fbb1479928588e7bd255b15ddff5f83f917d5fad5ff8a120ff8facdf1f1f1fcc6789fe270129662bf32764e724e6228cf7778e850bdb0765b990b79361266f687f90ed233aef7a5b0758044c79fac8d74240d0fcddcf1920c826a2ccb3831bde5287493b10524c30ea5dd2032794379c394489e2982feb56b2243ca77298f152ec861cfe132dfa96fa109e453eab4da310caebc11ce4a85dae2c44fc10ac301b13b75902173155812f504ea05260fc02e89b7e8e682fbeb67b658f8993567201ff58a897762516894e90e96fc115c6bc7780b42e98;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4975f5ad26f9960aed281f9d45df9203256ed416871c0cdf69fbad69737ae4fe4f3580609130ff7799c496002f09a342eeb3863844a5a1f0de0f39096b3556ad312fe4cfe82583b3678adad208de3af70b3d7683e5d142c976a8d2bd4d86b39474b6028630cd696f0903cd0547a69904afcad48899e3e5aea565ef1f56ac95e3466fcc11050c6b41f36abc472a358f11b0fbb2e349ef1d3d0ee90e0623077da7c7a636706d11fd78dcf1bab05059223c0d6bdb6357947714f0168e5e41117bc461702d81e1c99b8207946b355074e32929816810fbaa76daacfa68002eb7a4530a51da82c838811532858c6ddb2aa67c2a439be922c71f0ac23d72ae800af101cd51610489528cf1467b1913fa7512b39cd694b43dcbf3df28ad247a2a9a58d8e5723690f3a8fe4d2fe648b8b392235e3b91b0477c8c0eb51acdd422acd618be64f70bbe3dd92cefa24ef221a0d4968fbdce1500cf2aa3ac87c9970bef779c4aef974082b2f098eaef9eceeb425d2bb263c621e8446027d1563482e3274cef7005dd4fc9bb92bd7ca5a4451ad76b01216b963ff14b8d0f031282583aa814a5481a95195619e4bd1c1a23a0fa35ff876b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdb3237bdad85f3b8103382f0d88eb55ede86c3ab2b984478905a96d2240e8bf970792bcc8683e85a0127c2020d61e6915a35f911a91c7503cf645527cdb43706511f999d71851484e6622b48925db18d23fad383621d875a3becb57917abf951f2e5644a721389b702d130a486f9465e39e71c3ce00beaed4b82fc849806192d499f23714bb9b43d7c5a5678a915dc2a96d4cb76fff83b8edfeb7e372f83700c85312e4093b585079231a4549f9030b3216e02f5f66da304d0617f5dc38b695a148c59274dab55af108de40fdb9a3c5e9419233891391c2f37a6ee1f5258eec95469d5179fd1a1162cf4931a5b151f39a6703082448cdf58e40a95894d3e2a9bd6267470960b54c4209542e3dd7d02b77c70c3b85035f073f746ad2bdbc57b0320e830d8148a5ee740478ad40010646d67be678c00d5666cfff623d073b737ae76bfa25a26c38f338e28b7de331d68fbaf43830923f6c87d14ef708144275c466dbd469d807c1d52c3fa050850f4e0a14a14d6376ad15ac305c8f502233ab70beb4dc3cfbb675b75a23674782c81d9b83f61fa1b9799bb7bb4c721d4ff07dbda0531c7e314ce54a71fcaab16ddb34870;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6cf7ed6ab33c0993d6f705333b833604301322330aed5c54607eed114fc1832984a3fc464ec7436f3d26df3bb167fc963feb38c20055470d85b18f6cb1603922df38aefb538f33dd322590f6f5140cd9a62a6cd3460ff27516ade74cce9ad712c11a259b8452707479496a5af675278b36dda8b3422ff605e9e20a2b5ac3409198a40b8715136a54cb41c2910264de94ccb873191abf4a1a280ba76eafe4f33937e675a464fa11f5b9474f81e6d4a69fe1c5b0311bea17f8ec7878d2f5dc973afd6e4c46d1441f73f1eed43219c9fd22dd8c1908c4fcfa764853b7602e3b8ab558df7b63054083c4e13b96f7207341ffc8fc71618f6527a033d58ae707cdf34acec009dd659638dc75adcb3f67486fb8f8d7b3af8297a053ab2cd555e5bcb1e4da02fb4c029ee8eed76d6270e096e83bfcdb211d4dc9d5de7c57f117d0a0b3ce239d9f61690be1f07891c946608183d85aa7b667d66fc9f9ebd855c512df5bd4033981dbd928e569a0972e91316494ac6aafd3cb144875cd259a4f83878ec937bc324504dad1c531b75c6ef734cdfd2be38755b78067765f564ed284dd494543a8ed1303f7e9cd539b81ffc375b72d4a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h60d04aa9216c6197e3c2ed9fbafccafe184befbb12158ad621eab556e853ca277cb6d1a711e6f483f9a23ffa5facb3a010b8162e1b218677ccac7912a7089d2f4f10f28385b67861c2e88bb6dc61844b80c45b98481828f24755fb95f3b517cda5783187a5e7b256f064dc13193967be4f08c15cc03259b323bb836aa3de2dca6e7ed77b96975c82d5814b58164242e0ab3c732d32101dbeddaa2bcd1f5f667d8d76b8f094f1c47fa65912e095ffeaa624de270740a1918462516c1f4a991585a09e5dfe2d5b29eb2199d3fd925ed7397af3c0733b693d34882a859fc9a473650a341f18aefd4872045106737bbb3c1ed5a001c4f1cbc78166fd21cd832630caa5cab9f88c56ad2875bb5780b5d1cc618facf8082857e810ba9f218dea02c3c34c8d2f1b71abc543aca9194c46f3e54fca5c0d6106f7645fbf0fc0d2f1811a5fbd9d5be476804412972b06087af4b33d525911e2625aa450eedd583d8bd0796162fbc54ed7b3b3dc2c1bdacd5cbf9768fdac06dfbad5074e162428ff06f890dc4f400fab1794893e32d4462fec36d647733543c8e361e8fd4e9253bb6d16ce8c59fa070c90f5bb307d07013404367e3b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd461a7ea9c49b9f65d875a1924844d8266f8243b9c9422e53743bde7a12f6822b198d031d2409b6442b97af15ddea01c9b952f3de4c76bfee6e005d733de2cb47a239a07af587efb1ebe67df3b846614ae138d5c5881d1d133d507838d2fae22fcc90c1b5d535eacd13b6e7711b6d014dca56a0a5627c784680310781cc01365dc0da1d3c0a00cf576229ba26555fdcad0be3246a859e0d67c9e6c14b70dd88c17ad260b3a47b1725ec0105e703d790a4d3fec8d74df1d675cbb3d5b5828dedda1b9fbfe41203ab741f9cba740278f8339140528a8c61008b460702154e417ef4eb2af76c899ee2af31e55ad3cb7f7f31a6b70f41bc32e304b74bbba60ef7f0f97e01c19ea0e98a21b6380ac58a6f3f1dccb84f3a0dbf9b095dbe07a2cea3835593db1e323df59ba370fe69f6ad50ad488a4b3d7e8bde101c67abfcb8df96469814b0b9aadfffbdce1275bddfd70abd06a09ce28d91ba266647c22020b1ff737e6635d478d104df1abe177205da8fc93aa71e8ed40130c02236400188dd95a655bd7d7eadc99ac55a647c93038553da1ac892a63237c8eeb1e6f03aa5b168d8e499e54c33096032a8949bc01b1d4be74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h443b3c2c6f150b4b24e78171244fc7ab7a3e82d9bfe3d9d7cfb23870035203c3bbb3226182b3b24b3eaf80530b015418fc2c3bd774f243d9598156aee191c0428e37565b155606c3d0773c1fb2587c4cc760bacd664925febffc584c3ef3e260271dbaf6cdc7432aec6926953466f58e25174afad9c77fb9fba30a62a41c318a8f95ee5154b132db5f0969474dc9280e9f6d01b33f2331fa5c5acb69e9b5b379144e81f34c8a593c66336b341df0ef0b854b3db952dd2b1984fc5226433abfa85ce174b320a55c2df92567752637ed27b093d49e2b691f1af9a7122e56f3f204b6fc7ddf20e7e9c13ecdc078d6eff32fb785a305ff533c0d6a4fac5c8e4f31e840064d2f805fb9a4aa0accd2c8fd712797b03931bc0d32749ea9b7374d7e213d13a08c306ab6ec081407c19e508bd0d96cae4b1a0539445c3f8988f39764f29b99119a03577c9df469494164d3fa0850804da495bed188899ee7c67571de454f2ab1926184a6fe74e164efc1aca7261facac3e1cd079c5933859979ef3c741b39874ca2516fceb4677f9d502ba27360c786d11757d45a8e01580f0474dde5e7f7de25c67d3a1763a22f679fab2c84b20;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h259a0849f5a5d907d8bfda7624024d85f700570db2768fdac82fc0de045ece6bdc58e5c5e4a859a2c43c26642c154f08dd9cb32e64c54a28b812b2029b115dc89805c828ebeae20db30733e28b0ce698a954b71902d5c7536f85cdaefa0432671eaaf0db431254e52367b2d55ebb4a498f37af851a017dad2e0e0069a7d063fff11131f487b1ea93d58a78671495a3158cd0aa2de2ada5fc5349b2d118dc07c2db2bff213c4a22979ecaeff6ac7dd17037c02af5ccc21d3e4b98762afc574eaf63e5271eaca0171caec745a2e38335a181067aaa6440476c5d108f2cdb2e344bd0710856a121a155a380e3738960784e6d4c01aa7a84a2d5a09799172089ffada13ef82bf787311e2c0d54f766289129f046075035b8d080a00b7669bdfa4f1eebeba6748646be4f91fa1fc5ec856b87397b342b17f2b4d66294f0b27e8bdba1d24eb6dfe4ae7f9e837d844103383a0c63ba29ce1242c7eb39b10a3a14840ab3d649bf21e375fe7411e4e0cd4ad1bcbc66e31075e199df812cb36671b4069f215dc6093f43159fa83cab9e44fa50ebacf66887da22908c0fc684ed1561064b04701565e47bcd2d6f13f5d94537073f34;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcea5f08d5e4c31699cc09d07368c86c2a0416eacd8c7032faf0c4546b0395022d43967e91e214fb3369327be654ce9fbe70e640c8594fb7879d8cc7480f8d65685c1ade93902315703b5cb06ee9a909a916d555fb5604c8a423c1e490523f253040f851e681933bc14e12e1173de05a2a7ffdefff1f14a14e41ac0cd7565569c3a17415f5518ee56e157e3968a730fda00cba01da8afd0d7a126f227af76f86f16a4155689d830ec8e9727d0630976e5189a8ad6282343b4f061f676661a1c9df7474a2b36ad3f0581ed86b1e65f6d32ac0d750e946d70eb7b706ca24add9c7fbc66c86c1a7ca48c43bbff00e98cb3bae14deff6d8d511167a3d49567dc938d63a3c996dae337277d8f8b1fb9a962c7be59447ce09dde58171e65ab8424cc892158e21cc44b813b0d451ca56077ca2b10e33aee0c8c2b9490d493d13afd225da7d4e063fe4e58f377c18471ffdfe1c11f6f25a36b3aec8c09afa7d20c0e048d7ceb80cf141239acef355b3939b3b47f1c77eb825f2403f1ee7f90233b17f3ef9a7b1424d9a678499639c425a7a8d4cfc19b9fb0e690f109166049da871909589b04134926ffe6d638088184e789caa02;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdf460d6becceff416eb704e6a35dcc8454672f1fe441098cc787244a67942ba2c6f88f4f9ecc8cc45f56b4866e91704e31de62694e3f031b8cbf62266bbdf23deeb86b998bd0e7fcb2da4ffffb9fa2db6e9561fa913585cd741088f6112609429d261a43e42a844d97474cd81de8e7f51a1db518802ead2ca7fd731a76c8f8b472702d3d275d2257b233683ac2cde3c165c6f764353d32fa10924c02bce413280405cc1cb0fe0a1abe4858421af1a85d0660398622cc887304e2af1190b600dfead1db715f70d40a0ee67613db4fd35318819ebb1f90880652e48de93b4068e6c2ab64e420eb0ea3727e95743f84b71b4af0e84537f607491439e2651a03080e8a50fe6d2ca8bffdd11cb5ef946b664b7d73940c705da246fea26fa83d372a981904377efc091d6c407e35fab0a7c4c2aed28efeb730de289f3cfbc206ff66614b4b45a2e9bf0c8588faec4434e7f835c72ad651a150840c5470335150361541508f8c6cd15ed796211193f4e9cab0ecdfcb4c098b525ec750edb6055a934a96e9d6e0f06f0b28dd8cdc44b73b5294c1013e8823a26eba3af31ba8d88a12099e4a66a1b2e6d9ef16245d4bb240ce3f79;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hae3fe1c2e11864b17c9d06b342156e6882b7374cbce3e151f8c9877ba8b71b5cd7417dc69340c814106e7ca2640dcbaae31bb2538b3f78cafb2d968ca380d379f9f43f0d58e92354c3c770f030f943d8e8180536cae58bc838c37dc46ad34546d256e2006b2ea1317b36b5fd567f8849acf8cd2c13fdaafdc6e8c1a2c83ad2f5cef002161a4729a077b6a92b48197e26e8a5ed07a508c2d4e44b60311f5a85ec220dd1638387fac22cc1901713db22b617734ac9166c8e95fa75a98d7e18b68115803ae8113b31aa7091ee47ed5afc0859e6301933db8b22ba8d19075f488b15ba3f75f6173ea5e287e398a1cf6ba664779333d03b7e2dbf0547ad68ceccd1c201e1c76765c0292af44dd0607d361f5294001daa36763685ef1de25e139e35cf695acda5ea7102f1aaf3e2111cf0bda78caaed5aff9f856cb6176ad75d0eb022c715a5a0b5e923c0f48b4dd7f946e2a053b609a8f5e2fa015a7d8fb4131505fdba4e0352ba649bd0af10b974b6a145be25ec1739435726ee74c5675a4440c7508a546e0148549254fd0a49b811907094fcf40f62421dfb7393204a07e54ac25fd883028e1419d7978c95b31de9759760;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb1e1d6c44c64a7c22380e665843c610b87dcc6ac1c596bfe74e8a5788e756ed79d4d75f04aee12bb13f55158f7a879e884cadfe84d5a51a08af4fa1089b3b55540fc6e9604e43920a8c8d41a90ac2942b19a3076477eb8efdcd69f137478662a8218485c03aec9f66462fb93321d1e5cf15e54779cbceb33a4c6ae60ed42673736cb452c2b9ef40e7b1cfc2666daacd79eca70324fb5fbbbcf03fee474d7a967a8a2c8da8feb92a20c5feff7d4b41e0ec33b830a32ca43aa658b1e3a3d434732ee97111c8826bcf8a09930a86550e1c78a0c54e97a41452022c13623d80d0778b0b01883c4c9df12569b5f2444bc397719747b98dafd3cd2e39aec5bbd4ca3e6c64a91d03b9b94937b071000e29e4c2b3265aeff0f42d72c1b21e32afd5b44ae2616ad955d1194cd04bea57b1510deb6f5f99c0c51729c243c2c84dcc1055ff5a1cf6133d0709ae1519993546120b9e087b08488a6f813f059c75aef4b44cc8c206c31de21a770fd1d738511bfb68e10183a96540bfd7a8991656e996adc5bee0d5d2602756c89d163f6ac1147d28f9653c2672b87446941fa7222b61c9aa5b8a08657a387ea75a4aca81c20306606b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3bce41e642e29ef7add9a2678d1a85ddb4d8329797aaa3f098d40b9fa9e2e8543c90820864418537f2217a9f5d0c3cc4ced8120b6cdca4e9ff236e643aced3648bf792eb590fbac4dd8a84aed47926dc0dc3923f959f1a8f56e67236a5b83f3110a3beb48759fe8a8911794050ebbc6c02c720be36c94918b8d757c8cdbac1d6cc85c49bd17f63fd3a251464dd5cb82a1fdf38e276fd58acbe52249d57e5c2aac502ee8c3b96ce03d76ea9a02719754d12ca9eeff2eeed874fff4153a86f98a12bb5db7ca594b0aef442e7e82a3020e2fc7c461801196c2cb9ba3f566df2ff785d29215cb9543309c757cdbe77e9c9f32f370eb7a8bff4f09f7a9d6bfc6f39f2e6dbf43e2e846e48e2e687d5949d51b473aaab10c20fa500d1d025cdef32a5085a3b4d7408b79a635145c57da7909ee5cb69f98c186bcf7355f3c5635ac8831a771533354f1e1a1538c598f1f6e793bc9dc2fb87df137720573d67a77c1ed58abf0c8d67b62f0bffcbe3203b2efa2eb45b1f514a66e5c718c9c9f1cfd03fa05435a0238b9380bd4a95239b2e341e380ceeee93777c85410f8c1763b029df2f3a1870dce27085b7e344078021de426e10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h61d665e7b1e6ca68a096d2d3ba9cfbde018316a30271ab6c70b1758f055acb13c89c21f50a5aa9f76bd616930de66ee257e3d98bdaf334425bf4c468d90a359385ee531623ae5c3671572cf84c902bc6fa34f1b058ca3d4ac5d8cbbede4fcb950929a1e6e18833e5b90c895924abaaf2db6399587e0016301664250456a1f83be5f8485e5d73c666d7370546210116a0b6ed4d6720f283e205e65d75074de567a373a32565c4ae0c1ef1bc464328b2742a03dcc10cfa5f13d14de86fb25eabcc1cf201e748f87409f21c85de70201f733f03e0282829f7035598c00657f178fd51602bf57af295bb8adf0dcad1dfdb932fbb439f0ccc88b71845a34be007df9a8cd5797027a09db3c8998bd4a8feeaae780e522e929d41104ada9cf4236f952eb765adcac7a18c66b57a8d5c892dce6c7c35f4575d43cd256ad92ee51f1acfc3145067c5bc4d7953a9e5a9061155454923e0df1beb78f9d3399ca80c907aefae224f956537c46ee7c5a1efcaf3943eaf274a66378c7dc03c1a67c4afdd22e413683411fb2610b00d7d9c9bb3d18ef4a215482a7650cfd84f08cacc0d5bfd5f1129b55f606d07ac8e3881ede2cf7a627d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h79e24cf14f0d208dca0a679fdcfd3f34b6a1a145d340c5fff24a6e5488f1c68ca517e39167314266eb7c099f034f6c4d8bbadefd6e7489ed3af59325820fbd0799c07113b6875b3cd8c51d2794e4289886e9ecf614f3bbf877dfa4947ebc74d73584053629318b37c7b3099d148b45119fc72912c2de6bcc8ca020fac174cc5e41b85a6d7a73db0e9085af2b3e29ff5baea87720977c8be7c86d670d6ec094817083289e4f011a48f029a2a8f86e813e81fc28fdd860fa5c4d517bb5d2680518341ad7795e5b9e0b645a884b0a47351539275ca11682e9b16529f20075b487aeb1a8f350ed6fed67df2a273b9268e19b46522d3e36ef724074b9cb4f47e5ca78fe03ab8c7e467a663f73fe58d7c8241076ece5f45ffbd329f87cc1a8fb4b77cec177713d441dcc77d9350b667624cfa6dcb8865d365858d4d6cdc06a47343bb9560977b17bb2307cbbc79c6fbea44b55f04306320ac5453cfd1396d960b968712b92fea074f11d2cc3a7e72b9ebe33be5849f08e56900404bb488408a83d7456d9299fd165b191070c929e8fed6fd16311fff2479576edbcb755a2f851bc0eab9b9c3211850e889625909cc5eefb0621;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h91a276095cfa8ce1dffe110f346dd61f43c85f2fbfe00a9ff283e1d16d9069595d0ee26ba5ef12db7040c7e49ee39dfd184d6fec447196027342fcb667753c93b29a429fd4123c736b98194b323c71f47db8f184c3f273726bf7267fd0eb7eccd86ee4a219285380d85f9f4e2b7e8140ce3c1c8fdb5a191a87dd0d4fae2d5a02da703aac89e0873b7f31b9323f448f21ce8f70f482e1695ad940318e9b8a29efe063be1d4c0144f6bf91797f78a80b7b7b5080f8fc653c759a52817d9117810a3b1b51bcc51688d6a51fa7eb7640304dcb9c3815528f55515077813ee180d480a80e898a2353d78139de8c784b1521c1d226aa1436e924bf3ead74c7adaacae7bb3ec3a62ee4c00aa963968cdb63746061fbe0bec4fb26797b15b7321bf73ef1cbd6f2b64316ade4d19dc5f2e3152257649d20dbc60d5d884f28e39434c2081a593c54e57e166b161f55ffe108a73a860abee7f4c9bef844b163c7bc8779ca0c5d71f67b1bfdeafad0e5075cf0e064a08a71549bd2f82339ad6e1a0329f415906a5719c9a8f3c036ddc1729d7bd6e6c8a11a03369c4324b5cad5c86f0119f318f9f8f41f23cb834ce60d4211ee0dd152;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h82200473595eab6d5bf2ef0606d4194376f95edeb9a93b0e9e2a59b9d1713fd2e28966e332e540eab810660ff9a55c5d4697b18dfad60a47a4a9a7303c6ede967196d81db6679a49ce7242118b1071443360f446461f35bde635682f19e6b82aff99d99d325c659f6d8a26f7583236792be953a88690c3185aecf0fc2695111a324db11b45d8c17e6f2833aaab1b4b73bb7b057e84bb1e28d26d2ae50e78bdd9ba3bfc8fd011fee211a92ced47954de189c21e2ec0366468302a8a28d9f3d0da51e0bb94465bda3703625781f9bb4b332259f4efe12975d149087f15e867cb6dae7b800526b438d48224a25bf91ac0803edae16fbdfd00a1d89592e9a779f9bae7fa9ea79e461b567d3b9962853c9f3e84e90444df2f18c6eaa3159af06023f015cfc4428665e000ee2dc2a0c5eb1bf53472d99e77db5819e4a0fb3c027d7e24f5df410995be547e487948dc6b41043db3e80d784d59cf4cf149901e5173e7f0fd89a14bb11831370edfd6deaf54dc78e27acd638b5415876a9a2af481c410fe288d12192e5e4895d38ee48c92d9064e581e645c1e351e07b3df058e0df4e427020263ebc7f81a19c892d0d579f1770b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb3acbbdbb9cfe14c4d889ad7ed1da7a6bd859071cb08107f9c36c3e1fc54666244aa1bf63e491b51f5daf78345871fd631ce0039b7c0876294fecf0b3c5bbc07be4e20f616859eb581741333f1abb2fc9207fa6d7b022bb9989c933574e92b240e2b33303a5081d2ba4d9630cfeb42598a7f6e0cec8c76aaf30f39dfea0e085cb671869a53e2cc68a8dfbc31b259affdd1eb71402237ee9e72d73702899adc21f112688e8e08f338eee1e622729d15a7ff85f80653d327891ba3931bad0ea5c4eb7234d3834e552dc2377f5bb03f0fbdd076348e4618947fef23ac289118199f6e209bc1bdd066d088144f64ae8493e5fd26db686d93e5f990ab94d27f94c01203b518133770909c1c563b759ff562474395dabdae1115e2319303bf0d0a217ab406435ab9c0e31d1e7bfc6be4426d85d1da0ac9df23669779c567b8339e4c2e7cb5134cf3f7cdcfb98e997d9c4277a11ffb97bcc16cd936fc6e4094761de38e6471ec5942cb10d739c81851c5eeb7c1ff1ae5da67d867068d8b76139b70fdfea22d2bccac571c3a7359f3ea5177440f48ad8c9ca1b3f9d7cc97b62003f28d6c00c83a807b3edeac6235265819f3654d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc54f69b5320c60aa522252db4ec446e0e95178f3c8006fa4fbd7dc6d3825f1753f665963e75ca433e18841351fe330976bb14aef446ffd2e92127b10eb497a92c7bffd5d11a941a8cc7ecbb9a195b4c140af279d2879a7ffba1bd94352f8ab9e576b6a54148b0d09bfe3846e6c1c1ff465223007376f1c9b2ac70987bf19589932f5be17e11a75115b0861a68941f7c43888ee0034b605dee3f48f121c9243ca74cdc91e2b18f8a8d91f358fbcda36c1074973f8d1a4d8997203c610284c49351e011c0419bba9f0fdedeb81b58eb94078a3d43218ed9b80d1a9dbaf5a0a0774d058389b6973634e1feb886b9c6883b858d9137f46f5dfff489480f31c38c9e9ac6da6769652e5b5f655cae09ddd471d5104f214a5536ab240937910e7e1ce9b5fe03dae3d61c6eff6718155ccfe4ca5d5d4520c13c07c9db810a0b1776be8c6d5a8884840097cf17db0697c531eb7fbdd6255f81a94a2832950226e69ac67345f5fd7a5eaa6b842692b992e0a8b4fb0c260a60c8f64f1448b4ba1e51aea295ce6d2dba0bd439a9e1bdce25d7a82416b2fb6df9e0b90b69c38bb4baf93748769ee26a8132efde46949a10853df89b492;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcce363f1c2091d57b3381e8cbbcad57e65730ddbc41af13ca62230cfc9a0f2c36a50a667f59ba2ed414fa8883037b400addd652f45d4c1a06ea2989aabb4df80c614b3855f9b15edbc508a1f4fa8fbce13a6dfdc57cca10ed40267a159616cc9de5d10d7560270db3bc57d218c129b5708ac5e6f6e918d706880ba60b890e98371deb14f5bf93455f86a88d1bdfcd727136e68bab94f92c3063a9065b990a4889abfc6d3ccaab625355fae414e44041798935f49cba048a4a87d625423da52fa2e76a518f43fb92efb6d21e6aff755334a55fd120e5c5fa36cdb84155d5b0a607d51af07bd97fb6161641d1560483068d0be7ca0f04267d85373d953a31384fd53e92e5d4d5b9a96a62f4364839b797773740281e8c739c381c7cc89d025401bb285f1195a6b78daccba37f695654fab1d62a46f0f6d17737affc38085f69fb4a5d42cfce14487f2a31c8f26e1ee6c94fa0fcec9b2ec8e334b824d7006b425c1bb804f7aaedbba246f1a418e9198ed96986c66f675f385b921a30e295a0901967a20ab66dad7baf5c3dcfe0386d9ed09ba7243a95813cdfdfff009a80e19ea78f1cda9df6a501c2bfcd99fda1da8f7db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3a4dfc51a4b4499b1ae2ecc166fcd05cd94f85d420e3fc83853453bca340cf20b16528a9bd799f5defb8619dce35abee842410286deecd3fd0cbffacfdacfb28c21b0f0f1ff5f22e60aeb9f211ba1ea0b090df047e88ea288c820428c5dd890f6d410b6243a9aa1c8e6ff3d86eb8bf459e2fe843ba7ddaa8e4d45b4d01d2b9a292593f0e70c7d76a0090a28949779bdd5520fcac5425277e70e9371ec15170793ac86ab6867a9f888b3f1ea774296672f6e2c33b0744d8923b79dd5c1f52c4372b504918d2caea9a3e7fc5c79f18af00ff1861bf18a6472aa8732da2e7ad04a134f690b2b4acabdaba9b5357b5aba9798c56f6b274ca97f594609f291e50247067cf67e741daa13f23e819ecc7787df79414d566dd5580458137ea9d3a1837f4c07bc46b51aaf3f6a973acf46785ed38626cbb6934ed4c798ff0a540e913b7e521aec4f06529f5693f0943d39497688134ba7d63bdc1db6bd94c9350adf2e4f1311802c7063891bcc62e2774404fb92d53cc601513a1460b99cffe7594ea5f39092f50639d8c78322c88b9d4a85181d6d52aac0ca0eacbda7c2ded012d0085d5a9049695828d6bc3c54f0a5e9241a0af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2017eb8a624ee861e2f0716673e628bda5a0b4fa4ea499b78b1887f77f0ba57ac8eeb8baf3de849af952358983a265a1bf2a52f165c7b1181c19a2c64dd15086294dc86dc5f6967b284280927cd0671a32dd9d504f2a11bd587e2a3543fa169339e92c5c028c5244049c8f93233205eef3ba71a79d36db5a129bf296268d8a4113d0129033a8db9ca612c7eff513ed7f01b87b018356da59b28554fdce21a15a86d2109416ffe67cbf0afbe212795c0f7cf1a3b4fe7f185a95a888fc9a180409f5d556db8bdd71efc51db211f39294ae11f9958b95f0f0b0f03d74eb248acc9a036a70750aa6a1aa68e7e9ce8acf15a2916fb2c7f433b140c8d72d6b435dcdbf387d3a4b9ee7a7f226a6df2c4977c0e7577a834ceb1969b4f91459cb5d48c1d7e33f305de1f762fab3644489a1e05cc266dbe1ab5847c6eb18e0ceaee48fcae2309f7540d0c0948ed135cfe739c4f230e707d5af2947b0a4113e6fc723c043e1a7a3a81748549847478d5f2a10f96d1339960c2b6e8e52d6a86d915e0c93f1bc0500265e4e21c21cf88c7c1a0b76a33db2bc172c36073ff41921da8588e9b1efb331e03da238655a9b304b59d3544923;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7f4e1a64dabc99113290f1d1a1923653761957293067294f9a504fbe6b2056e5ff5a5a44f41073ae4170ddf12da131fa4df2a012fab8021ec7e8779c7a89c46bc2bcc401aa86f2d1bf92eea61efc01fedfee74fd85ca0adb48f890dc1365c014cd8f50c0473ffa72bd6ded6e4401298accb0586335fffb06c2c23070dce788d3982be6db6249e15e6732e6341f643213b78086e159efe16e3a76b5e93e09d1dd1061109132d69ce23b5c0789b72e49f25f2a05d4706685d488bdb4dda285760f08c14896ec074fa0017e7056fae609509fbbb509e852b9d1fb5ff89ac9eaee5fd997d5241336643b62a85b45655d428d2d7a67931440d8c943a02918df09f6208232a2d26f13df70a365ba0318ff44e1d0b8477a44ffd5cffb889ece55b69fcd0ee0b04855f3fe0fe72a9f6c7a93fa791179d6a9e5321f8fafd4ae1e52fda17dc3b8518de8d0d9a3e1f01092e87b14f29c0b17d96fbbc7270daf383eb624626ca7e2d244f02ca8d6c771d9113eae72460e700e49fa08df36199a3a4980db54eb8691b6f7f9862febb9c65f9d066d81eb979a64e2d0b75fc468e1b84ae52ae51bc3c4844170cf8c5498a1084d145caf3f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4e272d57cd74e9bc83a931a2cf2a78c303a7a19b3b9f90b9c074d2eb6ea376c9188ddd6bd3db19a21c7959594ede0113169e0016720ef6e6d75192d0d9af57b5d4d3c9d68d002d2079a47f4ec2f59e889884e47bbf42b3142d0559153c55174d4526a7c6bde31e4c433b2f581e3a4ae5d862277365f93d8218e7eb5574b507774f8b0705a166b609535d2826a9190513b2db150d7c26cef1c35c70b7d78dab43261c4523781f1a9c843a05b54abc66e63e3c02daec099e1637beb34751c8d1e5ce8874cde52d0229d9405266a67ebea56ed2e9aade323b91512599b8dd36379520adaf1ff7b44aa39c618587ebdc932006d4325134a873ad057cc7969020a2c166d462a31f427256609c04cf0a27623b38b21c4716a4a760743f44774f296bdf02b2a0c0cefdec24ac4333a1401b321f6538d341e9b62c6017d8f1375f24a0676a740b86d5a9efe097cb230d7ae94181db8bfc4b0b6865292617999cba6062609ee190587ca949ac15dcd7340a1b9481b2b0802f13db57d6d9801847c14bd0cc1131e8d27f0949b33d917ae93be5bea3917707af7b14cb549e57ce1c1ade787509c1df12bd6ed895cddacfdd63708a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he93e95fc1f800de7b6d85220fce87b2e58f09f1e0a3fa57a61925f2a665039e5055b0699821baa613bfb3a990fe0e1a300454af24fed8ab6efbb6845cae5befecaa90d983563edefce11bedd551015fd4be346ae0df5b438ec9d5317d7baaaca27c797aab243e4af623463481479f21eecdf3729299e85b8bfb320dc007061fd4dc41256455005d1eabb6215e8f1617b2b1d597faafdece264d1a8a493a0d756397d4a688ab0a025310e96127a96563befb68b02c6ec3d6fe3b1f653370ac425c975f56600c47b16439345d69f72fb3544403f5943b4667ba31e94c923d7fa278545d8c0bea66bdd0cf57f7499ea70c352d48af41014637c495e0cfc9c4bb8ee9ecda6b0e3ceec07bc80746e6ccfff00ad4fa20458c2c6f1b5847860f880becfbde6512d794aac168929a216f919503a8257a35d88cd7e4f49cc79393f2ea07e9944a61e9e2be7cfca857f991cc321dfec2ac8836dd9dcc09cabbe11e6cdd7b61b0dd01745192a1c8b59f59b36aaa287d76782610df4e693c12d1369579e5de96115139bb9bea82d05877b72af690e6aa6d9d1787146acdac3de730b9bdeba1c9cbecaa0f119fa353a1b3b1c596c662d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h12e45d077d583f320eb775930e7a79847f9700da1aa00fe570c15298b713683112b0c17c5a717cb02f1c59269f011047e564df66eeec1747fadd3658e51755c345df2ff0b7b037cc1d2ad549873970e45dcdf5e993e200eb92c2e287cb226f69fd32b81c780333382070d9e4883b06ba5be414033d5e0712fc7b20205a7f559ee5bfde604871e54aa73bc694c3089aa1c4e9e013696288b10193cbd6b8898d9140fce1b159d00fb99b47d29a71b55d2187a49b5e19df3c07d5330ffed09fb05df2bb4f42399c4272fd168dada6ceca003cb8e397ea31796a0278d83a0e7e4e0edf9df39a8d91b22600b67692a18d5358abea9a5647dbb06ac09c7d596989c899ceba34508c2cd99aeeb545274c0da8fac7afe6dbf0638ec3af589a81c3a0298581ba22b03b02fc486c9af55a6dff1338fd8f3abef2091b8b0a8d2a82413d6ce187c058000b2434ab11e12868d09d4097c0de10b7510a314dcc8a4a905c6ee716b8278aab8be254e5192ce1c6cfb0dbe3963bcbc1a7a9f4dd5421f0f6912ada8e69a0f302ed1542cef1b8e6d57b5bde29fcfca76ee7d3e18e1de2a63f07338aab83eb58c48dd9287d8ea128b16878c4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfdb76d6b80823c42ccce797859964ffa079c800200ec313eee4b20cb48027cf61ce4e3c8255b5d28b91f8cf5f63220de070cbd4cbb760924f70c66ccdd5f3a4f2d9bcb030b87e744ced0d37e02bddbf04d6beae21420f20b816e5dd831e0d20bd57145c3c5f5265583a8de317dda38de4019cbe54d77e254ce9d450700d2a1d25d17806b0b48ba06a7fdfdd4ba056b667e0b8e94d7a84707612f75b1eeace15acd246457c07f355db3816da0a4ad8a27084bf248f93853ad0d03c2e519bca41ef5832be71060d4ea6de354cf661229804b6ccc460c7a24f8909cbded2b7dbba9322f469d0d4dea8776863a27b0e3ebf022e8e1eb11a1aa20d8fa84dbbd98bff55a3cd7287fc211e8de5941db4d67a075c51af2228cec5facc90351cacde5f944521662e370d08b18a7b16dcd843db358ba8eaaf1d9c8d1a154d744d2ac6085259da2755dd614b3eb667e42c421b5505cf8c69560154e8b282ef61725813f183883d14b3130e95a546d38d86ced59718f6fe691272cb878b77f04974872381cc74181587957f05c9f2d962b5edce8c163d0cd45f86f6d48ca4a910062598c778f2d78de4c9be42e961b4ea6b34c2e1288;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfd83b8140ac3c4e8ac8cc2db5731d4b77ac69c04170464ce0af52de121047402f2f44ea842bb25adf75538c65f3339d70cbb25363cc32ea31250362399ce0ea76c9abfa9145cb3868a58144f42b1fc4578ee6c556dd71cd398a4e7aedc72373c6a6568799029e4015f28c221f75d8a58080e5ff7b7456b8194aaa7ce507a545028b02ef43bd667b0460329786bdc33e5b078bbdf8e4edca03b35cb1cbb7663a71776a5e3ea2dd1837e3db51d6e541c354b5847dde718d4d60d26af29528377f0c5712e461b9a42b4f81f4e6ae23d052db8aae254af5b53a8c612b4879d344449ae8801132e8a18dc9f5cc70e0b075b1331bd90b0384f46b99a7bb2ec2c21414fd8920a2a68ff6666a6e270ab96001328ba2d073afa4ea5585382dbcc685c3ecebd3716c965c8b568199621fd3db3b2e21ce21af382a3f665bfd2987f609c432ebf8d4236c46547739efab23c2d857d9574397cd2ca5c1c27617623b1cdde8d1b347813d4bc1033d70875f9af9d22881473179f946ea216b61f7240699069e1442d72e6bf6f5acbe0192578bdd2c4191d990a7a85473e58c637c091903456a9beb75a11b6e07d7fc1fc652f1ec73da364;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h22e739e2229865c766e9750f2c2fb3af15b51d41841b25f746da252a293a4470e52c7cb3c90ad1837ea1cfd4b33ec913b8ad43cef6807ef5f0c7559ee5c24298cc23fd31c12b3e5fb627fa4e57269d8bd3725c1cf715b5bdb96a971255e30f9ad402d12a65d09beae51e9eee6674823bcfce6a1a725b819e2a87c2333590fb24b17fe8196c93ac4291423deaced8986c1f949e4a6ca20ff23e8197a461efab20443b39c65b3deb9a8c45403b19c8c80dc19a8b445887e27bfb0550b7f95702c09714c78ea3f1106964b7acdbb069fc27e0adc345c30de6da252c42cade406ea0181467d73b3db68cf9ac75a53b85fa74b397bb8d8c04c72daceb32976016dceba418a655d83f7b06ef3f3a3359d08da039c0a5fc4ed6a2beb565d919f850a3ac472c539494d87122fd887924d724f8ba99f96f86babdbf9122ce4008fcad47c80c2dc99fe2e885dcb189949495d5fe5ffac6500188c8884b186f96fa034144b9f51a7bc90d13b48c0b45d351e7df1db9674d1eb40f3c384af6e45407d391ecb3360ee2e6a292d88ff6ebf08a56cc088449fcaea747abef5284a5a210c6dd138662989afd5925d4f686712ab5f3d53afb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9e01c7f25115b0e10f9bac80b9d461b8dd9c7597b5a049d1b3a2e43d7057acad40b828086c005bd21ca34f4c0314d74eff8e3215fdb425308c14338b420575b83830dc68424ccf5f716b22521726dd4caebdbdc916af034d4539424c300c0e00a107607b9cd24e685a1db4dd7db4947926ae4a956448163b88f621fe1da82ccf1eba1ab3af8941955003f85f641e30a69b5d738b93cb88e0c0e0a336927bae5c11de38da283d219faaf0853d3b6ffd62a610ac00665547ceb410a4ca1c1535776a19122fdfd8690753cff78db482eb90aada1d620b92767ce2230032133718af2f0e4c2676c35a5b08f13bce50ec094f9ed82efecdb3294ab9193a50133b19d1a01f3617320a78ca20684ca2634bd8485be449d42fea1838fc891621ef80d2ec1f0c28ef425f6014cd372c72404db99ad78381c1c405e6a305bc50aee5ec5a6882832610f73ccf68420272faca8036b9118cc340fa279a9904a16f25b88afd65f21f8d2dfc71b41b015dd8bc6dfb345df9dd48d08603049ee6c57f530487e250bba6e556610f6ed0941301402f4c4a65a762af1cc8dff99c629ec610350493fac4f0a3cd4a3cc8cd3fa9237d65f30a2c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd2c01abb367be9bd66d93a65e3086233200a304be2b3910f975fc97372b685843506ece8401726177aceb37383e7e004c8cd4b76564d83b6771faf6a5e67effaa81527b7474c00271d8d5ca5bd2340117a634c1970308263339a8976a2104a6ed465981d6e6e74bcfa84209dc5c50e49d00159035893f13a31704a2f252f9907b7820a8f02539cb46abe80d7a92280901c1befc42d0963746700bc7f68052736382b5517dd722560f076d3e9adfe6a43538145452b0831f3f4ac447cc5cf0558dc71f52125c8c9f93fa133f5ecadbd89dee7a34c7f4a0f56cc8373373f208a4602507c207275ff0df0a87826d568172680ccfb7ce2d2831dc32923f78bb73764ea4e7f18eabee428d6cac72406a3ef29feca6150a7dc6afcbdbef284ba81cbc259eb35b14b19ef658b779285341aeee6bab34c6f3efdafd7b30c70208893fcf7f5f8955771ec95b517c0330dfcb8df152e123d4c8d81feef59a10cfbf80ecade2ed9277b6e6352b4e152f7b44188fce1f0bcaf0e8e82fe46ec45087eb9f25c17bfad6753c70cc7a4b8c13893871cf97e1d92cbf3ed3fcaebba7fde62d599a002adfacbba1bbd34928f850cb2b43deed3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6e9973e9de100e18c10d2782799114a1302ff7ada7849c7a1957ad7dd4fd5b6e7f6cc56e7bc3ba8caa52d096253be185a405a727de80324cbaf3d6cc642dd8fa6458fc5c6eba601f561090629090e286f88b9b93a9509f8540d784b5b5e9e33b77780f3cec716a1b26b980ab3792b427d876a29297dce1375a13086b87b283fb587f1fea9fb08091570caf4ee46925cdef01e19502654bf9dedd0b245e66037aacc25ac91f3902f915cd700ee1039898018875ba1bf1ff94e1f8d03fc68225c20d7ecef5b46ece8c893904471ae1fa0e18a1f65d141a30135515d50340058f61d3e1553c60ac6ea64a339d58f344300681cb51d114da810e32fb015c22f7d4b405a0e140fc808063c9e5cbf9dd204d80955334e6373aeaa715811c4eab42a4b6c38fa289e14aabe19a9a496f1168893c0e024051be07daf5e75f0f3820e1729f6968a7f4954ca9876697c0d7c5e8e92b517990ff9bab9700b304bf32895325badf87154db13eb96e022999551e648fbbbb85bcd60dd0de33ba5724cd98ed7e04c35ab5b1f3898d758d5cd61af4aae9720cf1a219e3878c27ab678d26a60dc197eab8f11f355498535c63f9faed81351d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd541adc97550bd9fd3a13ff8a513161431ecfba3bd5ff8447f3074a828b39de34d800b0ffca2369b2e418706763ddcebdabc4e352db14c0b5ad525c8f8bbd6d9a379363e338fa1c66ae85199c9d82ec84185188f9441adb7e53ffa3d4c3e781cb905469f4b6d29701052010b96d917a1e2643e715e31cc7328bacd3e5984a111f9346281583542e3a5729d3222cf094973a9b9e3dc7c7106b912e5b9be54661da3d5c9de5fc4ded26f204fcd181da8098490b0038b1b9fc647fc04cc70e7abd1d77f74058462df374c86b0b506480bf4aae99c666b3e0556922351b99bbf19f15f0bad8ad8cddf31ab55354ee29712f36e53d61bea3b27ac767993dc703a192fddb148fcdfbf32a34dbf04ab3aa5bc34ebc7713d11f840d64a98611841571c18ee5d39b3c12d2aea04a46ea45fa2e178b5361e6f0eeb66db4c0a7cd54fa4ab8872bccc899a439b4298910ff9c906d01e03b7c70e667e9a3935cc1f806e5cc20f1ae81c3c6b7c581b13c32343ecf1641ff504b7f3caa907c195c43eab5288c70f0420f5b1f83839ea8f550daa28593519c392e8d33608964f2b32523f7898904d2b72b26f91357257e05eeabbbc1a920b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h556dfd55129ff3a1963024f8e0a42c9e4625276d289502f3a0b485debc6fea4c102d528e21684b55f85d469deb47d508ba032ab2939cfa58f3da1aed46e521c648e01e03db7d02ea05471ddd2ad63b8d92049ed27746797518567013f8ad7331e0f73e4ecf929a531b3e3eedab586d10efffeedfa279b5faf105ad2e73bed39829599db54711eacc8df0d8c69855f9c9ec17addfc97f906fe1e3cea958c9f5e899d0a7e7330e369af5d516f07a3e38c7ecf3890ae32847f594feb965c6b50b26723d61531533924c5ab0a8d1e9befbff52154e4759da326c89086cdf1c35663f808083fe8e2c5f3bc24e5130826fd4b772423880870f29e1965a500e44956123f3b98cdc6d1b56be9d97c20e57b8da2360f3b3ab348501131aa4b87df9b0985f9183f1b2438444749df74342acd933bfad612d3985232ea5a9e076ef461312b77a868fda0b069530ed5930638f7bd0cd15e0cc6e49b7e4b2010aace12474addd022ffd60d19f555ae990e3ea28260c3acb2466f80ca020473d32daf3d6dbf36fe39c95c7576edd22d9a5eb3b495be3f948c5495b0bc38e1ce680bfbd8953ba928c3600f868fcb188438d81fbe2361464;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h974c54c031f3d5a35d5fac22ee7b33975d647d83861ee1ffff82090f15c6cd996ddc2014f4d3bb3d74906486705965f2cbbd4efd1487ec4bd536398495c19aa1676fb981592a4be4d442fa51991f9f2694b17df14c71995746acd4b96c81eaf99732c6f0d6211732b42cac80705211f5e05838cdc9f0f160335f3c92db665cbb46ec4e1d2631434418e1821418b143dc4eadf5aa316e2db3adfaa0ba4b86d91aadbc94a31b4dfd3df61bf178f493e9f72a659c0491df5d47353e39d977875035c7d4757c05fa7abeb70dfd2372cfb3f24eb765654d6fcd78cb58dff1f71e894c7053af61318593a54fbc130026ef6d722bd4efa90b5b571007bce69f5f1e8f74cc5e4c65e57d3a6f5cebb9e5a3121a8d08de35366e53328f0f7f35c17b52961c57d9dfaf7c956cf78dcd5fb320ba9bb1b97770325baaa2903b8cd1d9b9e0b31466f81f4f7a2f0d6e55d48a55f998adad450840c81ee82f120c9b8cefce2b0a72974d02690557a3d4a8f15b8a8968a37f2cac7591fe99041eac88cfda96f9bba9352dd6256ef5baab544196b8fbc623ca60994425cf8398a4e911746b7f26bb43df0f0df86fc5618a64b7aadec0b08f38;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc80b92f54b5544bf33164a019339c0d2a1c625b92875a5923cc3c16296ec53ce185c6ee2bfd55c57bb9998f847ae462ec2f29ea14957c79b5d5caed4ce7d229f0de94abac607085677a0d272e18f7af980e6eb85cd02177a403769b88ad0f1cc7024d776c91d5a4f9c21b9b65b43f13dace36a61ed6f8c2d0bd12e6e06a46c83fa0a2ac06d6c6ba41bef5615378677e674c45c12f82f0632740ad3d527b5b4eb93c87252f1edea7dca64d80c53253570ee1727f1a7ec9be8bba4444e00a9d3c6e89e8d38e679c739f1f0701baa7ddc3c6b367d558496bdbca55cadd98c73eefa45e53d2f34fd2df975d2077a8571e6d40c24b5a609a838d6b0d003dcf841800c430fccad2719ae16d8e3a768b44d01951120d92cc06eb1c2be630c03f9cab81f67267ff0d12b28ff10c797f7486e2d86cd4c8b28a351b110293a2b375d96b3d3a3457ad4981d86ffcc7caf3dfcf405e63a5ae6fc12dd61d5e91dbf669da2f0fa2d68eddf0434e96f1d2aa55ff9a331a6964ef8a5b8492784e2194b0f642064bce469b8898095bf61c257d8b17a0cb761ee4cda6b64464d9b62cdf36cfd018bcfb7acb7fb381b3b4a3014f3e57555ad83;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3b0adf35bd93e255d029aff03393d6d5a7ada5f10273817487ea8172a7fdfc99fbe4766e3f1a3af0d2fae0c05101bb04c9b5f4409bf4af7ecca9f361442e381dd48486b78782f4fd6d0e2dd1e7d9a426eb7ff22512be4ac6672fca7bde695696edd02acaa9478a3e746ca43addf90f35f60206d0972d1471bb681b93621145c4cc9812199f84fb7ff6b60d0ffafa844761db281edc8d09ae6f6672d937c771ec2c3def46966706d0113e8379344d6370f178002f2a5637a46250bda7902f7d273f16e5fbed11e7c80af0a599becab6a73f302cfd507200ed73e158f7de47df614016982f1c317e847efefe6ad994d725b9e7b16d9b830f07656c48b5915e5130a81e9fc54ba3ea5da6b5db5e30b896a068eec293b541ed75e3bd56d84c62dd27b98cecd127f7496e736d37c70cf1b324a67270ec8482e782b214a7a83858e5f2ba7439d03f3ec53790f19b81f6c541784585039b269bbddc82a748b051b50910acc31fee7f04bf6ffce0fb74770b88ef92609a48570f6a7b885d4c19a64fa4e4a4dee8869117cb7db4ecb06668c48856a4c3807bd90d2239fd089407d12e3490f264692583153176e0a64963a5c64d87;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbb665853c2695b784a473923611c0e5f13965e10fbd4112c3c34605cbeed52eb98ab6d55ab469ad35b933866944423d0fce3a24e47567b3c629343a274e2021a40fad9339a652c0e5816cb8d57c1edbc3afa474e078b1847a860dc938457ad1d0e3a00b009029c262028baa07bbc2b61c9f8d06ce46ad4949d590b188ede8c057fddd6a823848bc499986c8a430692aeec8864959078ebdf1eab5d94b8badd4eebd5890263cefd29c555ab8acfed45f77816f58a1ec27364ff78812f2bd1368093cfb214ce6eb9560f026c6bd129aee3742cd174c213c2bcdd1993738558b0dbeca3b387b95b229e32fb8ca88812d85187da5fc065b67f4edc01113fac55f7f2d2232d26aea0602739fab57838dcc64dcccf10cf7b2b607cb6bdcfdcb741f404346d2e4379096cbcceda300114a99c675046c6d8db81dc4849cc44439f6d6a0eaba544e0972a22224ed2b773c9b496e39851ee3636e6a2e9ea2619101bd08bb9ef8161d8bd4c04f99facde8ed98c5d2dff29be182af2ccb026a99fc1375e2bf6a9277d1693e0677f7ce751d3de41191707b92cf79855106871f79244f5335b044dca0e8fe1314b46d4075d0b516049d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hff941ccf0a0de9d833f3f0767407c087da1ce998116c14cf4f422759a1a8aabce08502b1409eddfb5d9bca65e070a39dea490249ac63080c082e010b3a9c628bd3e781e5642694b944c8c43c536c65e03eacac7db8b71c667f0cbb9ab6833837ad51ed516a4c2f3ac2270bd2e19466f38228d8e3c2f46d722d4c84aa4c1fca9e5d422e5e07174f9c5732196b219a06b9d4001c94d641dcb3597e35244be67e26eb75726491af2b83fea6835ab566ee488bed567c6b60a6e6527ef1107ceeda8aa4c0a09357c8c08e7edccdba9f985fb6889dced43a91a2e9482c1701a3befbc90b087b109355ff571fddc104a9807a2bb6bf4b71896da0997daa5517cade27e7095312a5c58e3b2883795d143f3f794c3191b9b38758498d55cb05ceb38e59bbf9ca4c83ac89263b5a2f2af6b92ccfde870768abb23930c1639ac770274cec52b93e0b7d5509f2dcc67881bcd6c2f212ac5dff5d69b9222ba20b1a637b8041ffce43bd7d67b6960626b7616b47e5eb3d326f3c8a65bf3217f2b4ed65913aa0458d064b2451ca997aa0b854eb7cc4532c4435ddb269a9eb3a1611151ab55477f284c3966faca73dafba76068fe877c237;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8dc7337f201b9e3f7e9aff1b592f62ce96e9a19c0d7dcd1810de976c8bd22c0daac784700ac9a84283dcd4444d5544adb640cdc6d14ff861130bb29aae35c9a82788afc08e9b2fa9776f4d4524f7da63d842f63b90f89665c4fee944919639bf80ee0c56cff6449fe23f3a9438fd8a6453c476049e173ca8b6a5fa3b0b12ddd1be898ad0f894c3c19cfbaf434058aa861f2e5e7e8cd987deaa04c0a1325a3f5edb3bba74b2f83bacdd4d7c4e9f52b380c5d9a223d55c9e2caba20a2ee7e613bcda71f7d9d7e815a83797e8f843d19e4193191eaa7fb24f9b5d2bd5cbc2818720973d99aba8ce37843ece78ace8dcb6659bcbbf6730e90efea0eca008529c2fad5cc59f5b38eedbea4c47b54a99e2a5b5ad2369905dfd0fc8e300ef0b7fbedc24ceb5ac34c052813b53dd40fe2a927a51aa3fab360feb0d2bd315c299a653c3d46193883f0c5b62661d39b4a2c6ae51e16e1e7dad5c70c63e1ab3b21ad5e3f7f9a35c6ea8656b60261ebd8b248ff2bcabd5fa9b96bec75663b38e3c8df01523dbd8556aaf31287725dd2e66583bf7da48487ccbb4c92338d0a740765251a4fc82d02fa0d8cee3d33159cc6cc8964f58f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5b91713a6537804bcf8e50d3445b416e112455ae6482d52a5bbffe7ac81f990bc0c42b0637a6b17212b36e8f9d0b18066003d1e58f95f5959afeb706c8e1610340f3631e668e37334fb3fd4bdaeb85cb52225f73597c8882bfd6a5b026f1280d37a8b78e160e33c5da1b97a90ae5129cbcdb9d00a0eba394223477b648b95c3056948bc70b019981ac7d16bab59a2d1f2b233622310426d61d6a99007a623c95179b3db9ac6427606ba81169488e1108b46a9c9f64e9b0901216d2e308b15461671aaae47ba8fb797f4a411b8b0ab334fa9e23e50963e0f24dafa4116aff44df6961b5ec2737bba9e8c7e4aba72269d1e7e5c1fc466dc25e4dc5b655ecca098d536d460543b238edeb7d31af3a37c78aad5b0454250b78989b34a8e9140e5b42b6261fcdb624425adf0c71f1006972e1c6446a45bda0f1d42cf82d93d91623a9407137e224dc1c81a21ddf24500a9b292fed63cf8d11ef13abaf0cd9667c2e96f1bd7527fb0be0137450e6bb093ea3fe185d176b290866b533108a7a614c9c5cc555bea7e010f5fb00cbd1e52d14076fb68e3cd12bf0234d3bce811251c1ba87975c3ef1805d424889a7323415c0a8e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h55ac4dca745d1a0e018dc0dffef271574c7049c4d5172593e56f37efca5d971d852c78c83c23bd397fbeb8e455097d75ad0d9ceae1fc516ae8c146ca6eb9808c294d5b8d6000214b2a3c85f2d0dae389051950d750ee552a60d035ede4be3a232f46c820b7fa06a7ce12daaa10e6a489c197f541348e89872c55e9fadda741fe29c92d2b6be6e65a8215e881c97f72dd05275a5114189e33c549a69e388dd9ce487250908d9aa853aed1ebec7b7ff6ea6506edb3bab0ccacbfd576a393e221790604c7d2c0936e0f896c60efb2603a50e3b28ce927990d28b0bdcd89293d78ee7924746b0ad1e0073cd000126ef79aa0656448bb4f623d43d2003bafc8965bc57fd9f1c8e1e745dcfba8277f2570dbda445892637dee0a90d196b7dcb0c06a7a31275f41e4a303746cb6997f2beac0b8594f3c92c3dbbf10d51140fc1cbd1c961e79def4c62ca19d345f6aa3db204d961ce0910f33336e18c3b5e30427340be45e130e70c540fe0c096deabd76434b6a0c576f7c7038625b7bd48dfdacfd34316d9a21845b45b2680bfe6fc7074a87830abc19dc9b4de8bdba3da8afe919c855809cf24b8fc333b87330495ede9e4547;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h61a4aeb9849aacccaa504bc99955acb68c5670bd03579a3dac2057dfb13cf20f652bb6ea82348465f349519560ac99ac8ec4388f30b89f40645a84ef5866b0883bc3f51b2be91c591aed1beca69c9d150b137301e5ce904fd1634490107c36d5afebc83d66ac009d0606af97141e466772f926a0a4ab43e552194f43d4c816a8c6ad25ead8ea11a9fa0432a6898976943a2de48dba0abb0c31d1b09155887e3f8f7c4b848b79cbd6f69f6a387f0091b9397ac1c071a29258654c002295285a712c6a39f5a74ef98d8ef98e813fa17a5c4c9cd039783215e4ff43cb6bf7bd232e704fb7e81eaea847050f664a3f4c8011576aa60e83db29750328b09b5e3861ec7a488cda5fe34dbc1584da242fe8e77c0e8eeabf4de5400233f338a0e8494c9ee1ff2ba409f02d700172e038c0a2b952d6d5f688d11d514da0939c17490c5cf113b78e1a27b4581ecd3782a1392444ca57bd8c04e93e96e2387e56df5b5081f80c90adf633cccde67cba5b6ef8bc1dc6fc7cd836e20cdcf41fb05ea80eb6fddc4de1c069acb1277242d0c59c3424b6b7bdbdadba16b68b24e2aa94b4cd8257009197f1f572624b8df2b91213c7f69369;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha090155757e66ed5becbf0ca311676467841415e821689efd739ba52a62183a84affc9c6d08334be2fda1a2593f66c8583a34c8d5e5339114637b0f9e1e7ad38112939420d5e63885b6a355e9ded4a4e9e084e90a879a70090d3fd9505ca133e63deb32cf5a93722e136b175cb0f1310d57536c7edc1e35450279971ddf82ce73dfa0526d375ff09e3bf5f99ff67c1643133c306ed4bad49a1fc8c5c6a7065870d534e91d24bf867a15a331e50f02894b1ba29635322b4ee17ff9d0196ed055e4c54db7e8152d13cef05ee81b5f88dbe2b7e58e81725b9c3e73a9f252d58272a047efb67bb65de2151d5cc38d76ef2dae7e7533568368208cfc6087e2145065e78a6b719aa53721c5d571af1c8706917bd0ee9bd0f721b196ab122babef55ecbb74142326355e8916237661b3ef8f74398ec17706acc2f149040dde86f390e2bbd0602ea3622ad281406ae9a30d05fadad4bb261b98aff6f4ad32da9cf7841551a32fa3da1db6fbeb2556768ab916231d4ab0aa59a6fb8c5cd6d4aa9b00ebf1e62de3d1af87970a04cf1da5d01bd85be26e4bbc34e6f2fc360dd15ab1295a4aca37e9bf44c0a7c76ea3ce7900ed181c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3541c291057fb63396b383abf4b83610240d94970ec88d93bc06035a08ceecd09745da97104c5c5360b654f5928463d22e0ab28b2bc0cfc90b761066caba678783eb9124c3e1da07fb64713a73b5f10129e6ba3f3b705878af73647cc52c638b6618cde28e108e49c28a8a0cb55866f35b92e8d8801397ade300e932e7e628f27d6de1bb118a6234f1d6bbdf94303edbe1689bd6a5648cca1fa23c3199bd2924bdbfe236492864da697e6d63ccb4d1f8797448ce2d1362839bfc07981bd2a71dfefb6881b8877ba35377baba4c2631107336e925dac0888b5078607c17d556fad6e7db49960358a04c7abef83f46305ca5ead569ea3858988adb590ace69d2417b14e973886270b9ab5d7e2bc953b7cca9b8f5bde5ef68da57ac69ea464dd6e5a78513012138b6529d43feaa359228bd5ec53a887564d6eed287b7015b237b9be4f4af152da402130b76801225bb679ec1ec6e97656081aa11c9f9e615f432ab08f90f9b395b9978edb5ec15888619d1dc2abb30d84a861e2c062344927e4b01d57eb1cadee30d4a953662d27621f97dcb3d0584de4a815dff5f6faf719ec841958e479c6ab90a027bdc471ad6af6777;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h252823c1f89080bcfc771b532736feb6f0707d2c67dc2c6666f48181d0016da28ab1c7617ad8f65f48909db78ff8e29f888a530e636188aacfbcdddf6dacac9a1a466f87996f62031b64ec6350a3bb6ec8cae773bbc03c6f933c2bce28e3bf401c91e73c6341793f57dd98e7196ff127e399a8276f63a30df5886715698eb97459e0304eb7d422ff00b506e8f7d4e6b034a57188ac877dd3913356ad6985a8eefe258894f35146f64d09b51c14e9ad7cd7e4aa603d07d36f0179278a980e6da015c534e24d4a3c15724778bfddafb17ef2022d351900defeacde57afffbbd24e738f3a67b8cc4ab09a255ccc52a167264089ca5b9e73ff5166ed3d742bb3091038912ce38c13e168fe9e702dd1bb6ecb0b82a7a0b14a5bd1a5ebbdbf6077d16c6da6a9ad4f364641882eee6eb6db13e85ab706cf6c9a7f3cc5320e771e9f7b5bc214b9c112cf153eab117547bf1991dd6cf7fc2d70824211cd33292aa99d02da16208c6f22843742d123d75a8148a9afdf7002b2d23d243f7527d88038324c3c1f6fdd754d39ba488a0babff501e35a4ab660e8e22c8e8c5ac4eeb0ba98c5842fbb2d7c2becca94038eef15347bb366d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb46656c9865e6696f90f74c2d2a4f999835d9151e901d833e0b12c7990601f99f9eb1dacdd7aaf62e2abb6af552da0c71bb56269a7052fd5573a5cda3ee4416f444c14351777fc0bb38cea8efd12879e7adc5ec30245e13c2435cc2c5d2b7be796a7c539c5879cfb47e051aefcd4d273f888d4e6b3cc6360120ef7426bc426f1c71aa09a112a6b612d3fd62ff9fda4c9a4f22859916b7a2e54a406856680f7d7d6bd403c78c7565abde594bbdfb05190b8ae14934ce130ee7d741c0a3c2c3c9484593053f653aa8c5c69dbc1815a30cd67c33f2e189d3f379abf87f2abbc35a8199ee0638c389fac0cbcfaef7aca6af3d0a6db936d405aafe56b40a74675cc91cc19fb8b36e5e408c2cd95ab535705299e57ccf8d9320f0a6974c5b8916cb23508d6239529bda9c5283c68ec0a34cfd1e000d1f2227c0c200232a093ea00b5854dd0038f7e26c4ab9a8626355dd53544ae60fd3a67867dbecdd0edfa09216e05f9402c72f8153789f3ef7dc084ef46013315a9877404232ef37fa40920159065e6f1de82cbb8f7c0525e0e8873691ca8910be9f8799d9b9c0ca94de53ee9c4f1bfeb944cac62c3ede9bed2ca651992d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h1922d4aa50599ddbfffe1fbc031243b12b984a59a632b1ad811ec7d25203a5d030f023b794780b30ec5cec7b94214b9ad487cb987cd0c98daf6174456754222e727bc9cb286c49666dd31c2509ad4c4c565de63eb310b6870b81d6d28dc19f2e1d432ac7cae11d5e4052700d7a2f511907dd1f1557928dd7c6740c3b65a30e82feaf03560a3e0af11df17cc1ead5fe2ad09fce8de6ff98265e812c66361f58777370fb42dbff7344c53719ea3591a4c83a17a19758013ae7e0ff9d98439ffd2e60f554798bb0abeea0ac52f9d86b7ce0491bd0b61c98da4be78e2980d830ffacfcac96f7ad6f5396073cd41ad6993b862ae1d6ec965eb587ddb6e88fcead0327809fc62e6e3e97576a1825c43af485234325fbbbcbbce8210de9027bb2cacbeb0894223d32a9519a0700c0ecafb34bc1c4f60cf1b167d661bde11f4e6a97813be393c495bb55d54e9c0b2058a36f8942ca6b0779552ac62920b69b7325788f5c400611534b0800f2fb7e3d6d8dc4bfe40b3dea7684a933e2c58789a4918152071176b5a5df31e5f2d9fc25e01e8ed31ead3a1ce73e18fddc7ecf0b8ff163d11b787c63445a20b9d22d97f267ac2f1acc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdc376a7ea2b47cbf2797a79cc7ded381f4bdd1debe9b8bf6c00c69395dbcc162bda12def1cad4c2d8369a687cde252a9217d2715e522f4c4edaf114b5bf64a7b9ceaba788cd76e341ccc593f30b55285f8281fc7579b705127c539f0edae4a6d2632b0b7eca0848c976009193e2a7fd0dd32b161c3bcd82878786ebdd0c2640e917e361b3800012d5315203f1e0e035bb0c8baccfd22b802172a87b28d24c12ecf8c86c19f594f6856f2d57636a4f39d6c5cc8a61e4ec724f07262215e84131298c0b64244fcbbdb484893c4936c64655fc785b3833ae5b55b8cea4629aa9f5127aa57ddd5867ef4956bc2568ec46f94b63d64d528b2ca1df3e9b3e61ab7348caab151375d33fd35e653d4db5f5b1adcb20615f97801b2d38d1b4fbd84ea4fa7eb7a0b44beb68b200220c53b9932e96f98c7c5381c19fd2bb586769e5abed1a28a3c2fb77ea127a0dfdc4b6768b9252a4920a61495746a60f82a802a5414baccd335c52aa48dc0866e8e91980ab6ba845359d2077d920ecf9d94bb42542cab42303e570ce41c577baf1abccdeb3cb73885b929ebb2f16edd26ca28fdf46c445e881ff976128f17621d05830c255e935b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he5ca8e3cc23916891e66605f75c2964b809b823e48cb9ca4d479c30df651e998dce8c1a21e96d1d26e99e67395b7dc346b79b81788113b40655740cdc1d98464b0c816f4cfe2c07377c9fea83af1892bb9377b2680b80c903eba816a4738514d957dbd767ea9dbc279c9d4c1ee16b735c42cac7a48921b05685e041878a38ec5b5e5b7040aa74628f3f01baaa7f3debaa5320466cd50c354391f4d61439ded75e881c27b5ab1fa579d5a44a5d6177d3f8593deaf116b996950e48b0956ca0922851c9b688276df8d9c5a4de84b5da7d9d8cce9950164cd0ce37c6f4dd09171699ebd93c1026b505e53095e1d5f0325977757206909b31fcb7d91c872cc1a02a7463695668cceaae1c8a78b34495509e75d66bde191ee86cf2f449228ad499240f329b0a0ca733a5daba873682b2d91271af0bfcfe0019fe485351db07268e1fdc9ab760ed9bfe573f5646cdf6c8c87f61fa983fe1b73d52ef0b6c342b7de123c9fc0755043cf23ae7efb33dd13be5379dd792cb1c3bfe544fa70db99219e9f11aed093c7a166f09fecc71bc3d91e07f083e05c5270b29b8addf45a8f9cc7d96f9035fa3d7e86d8f2ccb45e1776903c45;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb93375f303c9d9aabd77e44eb4125085f64b39603392d6343db1e1012529424658fe3e1bfd7b0c5b265fe8c787ffbbca56e20443f54d044c86930a50fe13832ab6e0ded4ad2710a0df449bea8966e1784a529dde1f6a64c0531531ecf7d239f5a149091f714b7d859287017063b0d6f69e476cc5f37cf7b0a63f3d89db861f627ff634831650b517d15f35b204ab6bd8c43de90872a028b67d9e4654c4c8452b3aeee5417aae793f7f7431ec25a3dd2113bd479e3b1946a016205711ca52f2f9d06523aeaa1342b760933cec7ed9be9fed1697abec4ceb96420648ff10f17ea6042e593f316101f505422b794d496e485599dabce18c7d38af0a5b5f275a25e2cae9c962d49a936cdf0ccd72b027b6f2d93b7e59d572db3cfc91b2d2ca1ec1b673976d515de313c0967434a788c9a7321179af0879cdd438b467dedf2d000345d49f8647d8ec4ead37686c37634578efe14d24398ee1cf38e9a1fa42e34011d1795206f9cd46a8ba16d18223842c32d383bbcaf964c8d9c3706dcad8d297df9bf1eb9723bad8e93ea6484660e6f423c64ab6f028ba45d25d170212c6f50522c4d2a0b63840df0cc88fb13c831d39de58;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h20bc9e8aaa057f1b73d027d58f8d3827efd0f59da6f331e1bc938c4e9a2ad874f354d3714d8a66f0b53efef118b7565edefb76593c57cadb3727601f708ee827b076f01edfdfaafe0439a942b8c957dc389e9e40638c61f2159ec61e7995e9b59bda3020543c6171821c48e514dbfe78dbfeafb75ee19dbd78fc17a665be2a9aec2551a284d64a983df6049d63574085787ee05fca5701dcca1cb09ba777269482284121eddcf0420d3b3c52c59fe6d8da9896c21cf602349ed6f263ffcba4336b75a0dbbe7bc4191455706069b50667f1415258417e067806d0e298ac032724325ae4a0e1c3a52cdcf119a77daed64d0a2f6c3eac361ba38ef8d1325c0b8c83a67ee9cf02d9be0f6eaa8b69064a6228f9adeddda8f443ec5e644856fdbb7afe8b3d4bd11e555018d3e4bd301536b014885e4ff7bad2eb222b8c38b003f7ffb0cc5c46f07f985e0af30ea67852974e6a260382beca0fb38337bef80fea4f247feca217ca2a5b8be705b22ab5f7c0fb2c01fc10cef5e4839579e35790193317d39cfc7c3701723f598d06f2747722ccc400ea544478d450ae799ff327264a5920cae2b2c6bbbac48431c048c1d42a4e7e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf029efcd92f2ed9aef0d98b571e1cdbe85ecb39a5b7edb7b0a44bb46ac7781ae783a44e04bf5a09d72b70c5fe21148a0ee42a3a2cd68a671be2136ee2fb9cdcfe1a11f4d641114831881545a60d0049ddc7b1b67f500c0b0a4307b7a94903837c769e4f284d4ea09add99f2ed180fd050d83b87fe5b100cbc726b99b40207f4afc89cd10575b1b066638447401046eaf69ba3658bb3a4addc7f77d38207748affc6449bdc61bf2b1bbaf1c0b3254862efba75c39a1899a92c03d0ba853bed3318b527387493fcf8e1ddcf4be3a30a58b777e2565fcbea92b71d5fbee2fa7233aac0eb67334a9e3d72dd652c76e383121f94db0ea8d470cbd7ba8cbe7e7f81e3d29acc22522bbe90a9569929cb2f4523e9ca9aca4ec5424b0613413f95262b1b7b9786d9cf58f1454c796ec0dec3761270b1db4bd8e88add2db8a6c0e013bafc1976b6f7904e98f4488687d76d32dd6ed14a7d22ef2ed0fc0dd85d08f3aaa841df9dc54d94acb42ea72255cab96f13c135c59729b5113143370f56fb732d8882bae56450661689d5d998b0a721c339bbec957d9fcf2d5fa72a2a748833f8c90d4164690583872a91ca2be92a3c9065ce2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc629e16e145701248438eea8d13e3ce5b308260d90ef42265533ae6625544ac152f70bed65a663c8b002f4dd3c5cf7ab173515015d7fa072f2b2e91d54fb43fd1e85140c2d380c48f80e880c047067235203608909bac5850ede60093f55fc0e246a03d0595c851cdff6fe55489935c6767b08f88d18ed5ce3abe7412f66cec5bbd99d7c5d0a5c22a979bb0bd0cb4210716bd274b5d16466b3192670b2af5bee9104e16b85f1452b6cf40de7a15d032ed6cf2e59d1acea692d44785de7c2fa1320f2e66b9464120380dd499e0f14b3b6d523c2e52cea243e8b50cd80a133b83eb5cb01f90944576b9b48806e780e6ebc525730720ec56a10aa743c482b2f210a7dece4d5e351e23fa18282a9eb59903a9bf6e437a17e19b54ba71a2c89b157db357a052303baaaa292e75c4731d8a5c3f3e3a304ad5943b98b0882557b5f102ff6554f137edbf0bbb245b70c4d9ed640af7113a4b1a924b3613e6594310ef00f5c4bc17be8bee69134b1f0a393755ed426a8894865e0a4328c1b9d0e9f200f56bf6905b826a4b53e457debf66ee8dbede3cabc8604495ead5960c34142642ce1365ac45a237223f4562c6e3d6d95a195;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6e639e982c5974051fd9b2c82678d0f4e2a65e98f513aa9576863458e41ed6744b7ee876a002603c7970fe51dc51a3c7fbcd95d38de227c70237fed1131eb0b9a0f3e91d256695d4f4b2b85b8574f8464c5e2cf92d0eade2d88d717bf9dbbe8ffa56cbc48ebc9a4022dd921281e134acff9882f5acbb47ed3a1c485ade7b6e7da2de740486cc4d8b849873f7b5201f76774d43b643e5e114c4f4cea07f0ffcb6769a2d24eb4776baf632401b7438daa27693c346b2b47dde4c5b4b59a2e5240ca559447251d8037f607edfc22a943c27448afe2a6c8bb9ac7bdcdeb6af0394173d7bd378ee2618282413275457ba84332e04fa06a898d86922ce65570c0647ee8f20b0b1ee8173ad44a5452a0c6c7e093feedea86acac61c42a0f675c00d315a12b1fd48fa40f8526279deca5eb96e534a3c2970e6b85d4316205e63be87e1d579218961dc3ec3f43c1d7e795d2398da354438ea390fae1ad71e46def2a5f8d51335e219129e7827d342750856c6cff47f665fa6d83325f8efdc3be4781d3cbe41fd666b0a24686a93ee34219336799378c69bbb20380e33ca64b36ff3ffda3f9ba2ea276c63ef64fafc0d4efa9b016f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h32143e896c850ec026e06b4f055c78ea73a793a18c20669e3f709f16772e688e4e8065d919f0d54f3ec592dbc1df6b178dbc58fdfa9fca9b95b103aa2a2dc11f10e525b496fc1d34203c9d697f9f6851dd23c2ff367dd47ab535dcda09c11d1b8ad4b7048baffab0a1b6eb32712d938ae89e63e29f7a42ae0115cb84ca09252ef79bb21a2dde285851fde4aedcc0a51ba56304b136d6030238435a099b09615d74414f9efa63f7d0fa7718cc7a2fe8022f72eb1da087b79a74dbb52981185dedf91b214dc170c52ee98be32bfe0c51161efbddb28f09fb249a7b1e8ed47283c163d8222f48e6e50c761753127980b6921415da35dc7e7b9b4af9238ee0850caff8eae718e621a5bb5232a993067eebfc97c34b615245efa6d0074915fc698d25acfb38695bb59c6cd967af16711eda7c86ea225f36d8f2a99e686e3e61734be2aeaab01749d45926c625670b267108b21e4d420f0040d956337da26c2daff5004bba69101b94eed77c64fb67be97054a131221a2985efa1e524e535aeab6e4ad0eb597dab76c9c9fece3d5c7d437d58308d38d864fbed2f5a398a7fa33bfcb29bd848c20961a11738889c3eb4e889dcd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9a090be6c65fabb1cf3ab4dd5d2d56dcd46cd8a262358fbe8377f00d20b511e02f3b16d2ee6a10f6e43a332f61527a1f503496f66b03b6e4ee61627dcd2a31f53ebd8e4a04f38fbc8012dcec5c7ade4b00c975665e66c246e16d5a59a87be698109ac493e856ad494ef1c5333da9e863745548348d1ad424188e4536c531e4b751d0f6c7cf3997c4f2c3e66ee8e2db24df790f16055884cd36dc0b26dee8a34da643bda99af4b62fda275fb5b4378f4adf3d0829482e54432734d724102751e6ca231e689e3d56508bdc12c5582c99456048ceaa5086aeb2f3047b19d89dfca62662bf6860a38a2aafaf633093ed20385746da1f5d2c18de81c5c798eac502c811b87455ac0cb729ff4e377f9467cfda0ef9d97d5322394232ef1e2b97f089b5aec2122ad8f175e8f5be22e455b336ebff0226a684307eb46cdf95ae62fa0edb1f7cf3bb5c3b4fcf4b95bcfb2761c6c8990dceaf136d470b50d30a078430de2643087686e12f7851026eaaed0cfd311b0dc47146afa594511f3659c9a2f99402568b4fddfeb79c1375cacc261d63a07eea09a0f88c6f88b516145ebffbc1da80ec1b364accfdf3320d424f1932fcb100;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hefca20cf9c113bff7147a4b50ec54927d17fb81c9dd0d81b0606c775b36e9b023dd28d03e7069430c432576009975125905f3a981f7b1be3f89266922c4b92f04b85dd29478e6fb0d2bf2a38c3786f006539c4a8fc0a8bf79c6dc3418374f079b895abf150a4c7229fe5d3b107dc0743d7075353468b77f230f21a359f45e421dd09a9d0d2391fe44d71852ecd75c6aa4a23cb68974e66cf54c64ba7b00675f5603495853e4d6ee740d7949ba18463492d056b04193f7ef095ffa84190bb1a0eb193f160c39c920e0aaedb6c680566f11623510d519f0422e73b08c28d3f5d9c268645f5ac2be7b4dca262815e43f71afc1a6164e3dc1c49c33768b56f5300d7d0814de8fdc61dd2c06e0703b03876536f4c309437bab9f914474ac7c65628791cc5144ca3ec28a782e330372f8634fc0be4c01980aa76b7556d616b3cbf96f93cdb24e834534485f850e2b8ebacaa1178a6841fadf025183a20ed56cbcd8f1fb60cd7ad9adaa183cd3b89c6965286edf3d50af5cd4ff2d2373bd209fa28d373ebbe7fa406cf12729e94e0134e029c04ef259b5bcec8407d9065674b690fe60c12cfd81a8fb645188a84869c99c8c641;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h678e2c89876683ea54d293a3246c93b4859663d0627c5c7797407bfca0d6dade1476a0d79382fd8206421e314a1a62b078d21037ea5a8732a83cb1984b8f0c3a79ac6b8dc2937ea5756c395d430faabaa02da4e4e8bf28a80465bcf9ca228817d94dcafe81f8f1264c181258518bcab8f012dfbcbbf90e9fdd79d876a28a0dd6c3544a028be196daa39768d8daf0d289ea8c641ab6f871a43343eb9fc5931f04cf5ec643bdc9a05cdea9318ebde42317843cd9885643d3f2d7c0874e00b1d44bf071108b0e00a1523f33c35c90cd870381c11f4e9109a5fe79219c49aa8a3dd2f857af1de37deab81156ae6c49cca39a1765f88f3a85d3964f779b09d1779f7654923e9db7c64e16c13d97fa40d9a67bcc361f239ef01cbfcb70b7b80a509d8b36997e3a0972249a57db43cbaf056a32ba4a60b646c386c22bd4a5266aa0c660f713386144fda95578299ed7185ef517d31881bbdc09f93ba2f270c15e752cd3b4745f51de0a8a30b2410a60eb7bd76f5cdb9a7711926faf7752f2f79efb3ef86394a98820acab58ac97240068ecc8fe41baa7d2603465ac48fb2574cb2e98c257796ce5bb2aea18862c7820f777ad69;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he7e92b693d45e37bcf0112e61962555146ffcf7fef8d6a65e50bf1b6483772cbe6da5e1e16c57c4e751f08e866436381faad95afd35f3e8e9d6e87207c28bfd9884bd76332a056ecfdea7aa42f3682a561de93ed6b3dda839c6f0227d7ef34e7141c7142618af231ea0b2217d1b8802299448c7b02c0804fd0edd5b9552feec6d75084cbb25639ed55d99ed55d0f03abc272900062fca5bc1ad411ba35f00a050ab79f15f0c8f8a52568abc84c385c376b4ee27c3443466f9270f9cc77fdba5c315918d5b7fa47958bb9076f646a3065cc6151ccbf70324fe99fe2bab60c581537ef55baa8cdc27713ef2ffc8a3ef0f44e1bb626b457e3b78b7d39054dabd3509186119578a662bc9cc9b0575e4baca6761702b84debf3d37a5a342c87fe40369e76679e9dcfbcb79c7a64df248e4e284f839adc00f276ca4895b09d39795a7099482d65f17d51a8e1eb59c3d69c764fe4d17a00f6c54f3445087e55f3bca3749f2571db8d77a52d58dbcc53cafce4931b495025af1b5982a34a872739b5706d6f450ebe5ac95468a4ed9915e257640f52184aa9b21a1ebed60679ba226dbe669230b88674078a40d2f268dce22d02a9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4bf00852159fa9a3e64676a613324f4005e3993e8e732253bc031a0181b0cb2ff26ab7f885881603d1d41cc31e0ea2c3d53a0846a6f2217c4b9a5db37bb41f61ad53aa6d4f96f485e0300b6c4d14b58616585e7b867fe6df0776dbd07fda13872baf3ff3b0b56869c7f2c300c41cbfa1151412515c545cc3fc5232430263800e2730655ef43fd423d2cb4995167095726a6287a920f71444ade52c8e0e1f9bca51c5df3683c7b27a5ade17f3f6f0ace58a79fb1afdee96a582005adead23a9c0974dd276db8fcf2519bb69cbb61c61a970da7cce53844d8f02d9623916ce7f241dc32e7d52d9dfb8139b00d42f621f0f01dd7aa40ebba2c4e51c0d5ca87e150d3a71de49ffca1f7b105666556c4704c19096cb84b59b9cecb2145f5bbd878f30125d95c7ccf71c8437c607e84076dfb7323aea88589e9c0ab53638006522f9426d706de278e58899d83047b5940b39752728b550012d81bc69cb8420068a228edeae6d3f8c20b718c011c92614cdcaf725a05347bec24de898c6048c0471c7bbeb8cb819b63c02d3aa0b09fe3a5b969e0e2ac7f62ff70e4792b0c211dd193378fc5db8908ab4bb97f93f66c8ac5a1893;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfe36d65edd0fd4e8abfaead695420f65f3d9741ac47510e004bd4234bc56533f0026fd08259f2a986525e8edac217e3d7d6d92b29e3a3e33664dc1420ad8dea34b158bf8fd1660e5d340f7f5fb3ce0533346131ffcae089cb77b66100228d6947cbb3421feb20fe588cb868a523c95e70ceb315a80cf2cfe7d5f99c3db712795e292a1ce57d66416f3aa33b3ebefb6c54b400e6da997c0d403655411967a5db563c0bfc0e4f9559679059ffb8a3a345cdb032d9da2086fe59731c28d44ee006f12a517cf789f5c4be650b57254f272d64e1d6329d48cb8e7042b452ce09840ffb911c3eddadfba0c4635098fd297d5dd7a6ea169f497bd21e498d4455f0b7a73f397345a839e31c5868060f35fdc159e8bd36b138679cce582d94782bfd2a78f15d449367d274deafe9211743bb5e0d5e5f4a2bbeddc00d0eb76b81d3afd2ae2c9e13ec914bc88443656084a1285098332dd5c740f4db5f14ba044955fedaa2576d7e732eba57c156c24d35b087b788bdc71856c95e379564e59cf8f640455d1590708a522e90b71f5375419d7649fad99825666640dc39b68a984b592c8997ac548a4a59db6819b095650bdb673242b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha932f1079fa5be135d6b8f24e1b2b2dcc12dc1464d291ee342a24df816dc392834d3c199fea1b5f67bc7d8d763cce0c5ead22e416bd2fee144e3ce496f698ad8573c08cd66ccb4ddea26ebff4df3ec54084c001028050ea859a4227178223dbaca7d700054bdd9db237bb650868f03faa444523f43e57bd597ec4c48ef1acd34d9e8cbab93f0788e033eef2610b9b812a336fbffb36e6d9a6357c39a7ace867522bb90588e437355ea19bba118d308594026c73139d371510a403266ea614fe5d9c861c6d15b8bbf32f3928d67a2beb8987f43ed1b4850258a60ed058d76b93eabf9c7974c7988c30ed98ec7db798d329afb44874a23b0a6586fa806edad4f268596bec6ed84eb7ea2bada9424e4190b4b70ec6e05a16faf4457ca27da859e1e60dfbced374898432498a5a294d6accf18ba7bd02c1dddc9921c49affcb479894b89565cf23c34439cac4c1306193707165c6aa6dcf0560c431922e790c1189286348d2c3bbc0bcf7ecd9f6cf4686e6300afcd95d42b9988c43e2c45e9eb3079c390b70528b70f7195f6737f1ccb0640fc0f33bd800f54ca590e05531f534ef7f7300804da5f93a4250f2927fa2ed46a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2d820f95da960d03be3c30e8d65ea3f744b9cc021a6710d464d01af0cc2b3b6e1a25a2538ce1cdff88a33437be3df959f7746893ee502bb6154db20a1950ab0fc0c7bd0606f0c6684b5cc463906535d35b1878261df3b8cb5c2b63e127c5d3ce04b9e687a1236ab04e5634ca3767bc96d13578a93a131dc5d00b34804b32aba01d02bbf1fa356a10a534022c998627425df040b4893b34d5686e30f9734bf28f5e160503d9f47506f98d58601c3a2879e9c7f31ff090bfda47c6c28a4e40e96848ce5fcc6e36f10de8bfccab7e2051f4f152865e89927ddc24d2a058f11d8168bd03b1d90a2d9ad996f99e8ca1d1deacd61cc5365ac3b11646d93400e1f66c2c6d9dcaef43816599f4ef2c4b1446ce50f7b1c7cd68d6cc3028137e2bc33c528ab3caf7f445c17d4232e7713881ddec930520948d0a78eca8a5608059b8ba692c25cf64038ade6980f14b3fe582ca317cee9e8d555a64bad6f828de23eb682a6872cf11915c9827728f3e49dbec74541e54a09750a788a605d37a2eaabb493b04b6630bc54ac0aae572fe5e83d2aaaf7ddc8f2eca0fb2a10461d2b27cc451d0350bb23eada1c34891c116cafb22b15c64;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha7a5d1d0b3bcfefb0f51ccf050ecc2f098baa1a23e7ecabaa781e45cbc1eb99c05f232c751c62ed7f832cf03bcd5160a2f95ff06e4a3f64243562aa1a22f8ee0c77651dbac76b31c05cc716411cbf2206a4c3efce11277ba834e5428ed325257230279ccee138a1f00b5cec910b4c99fa4de320c8bef19a111f64650182e34e90b36f798ec316e1299bfa67b160435c0a40dfe89cdce7e394487e2bed46febe38c713db161b3f53adb86d70e6eff8738b760a0823970e391f3ac12c828fafa20682058a30139c810001434b2f8b8b4c99a8e5c47e5984ea99f63a50bc4ec12d11a089bd491a32faaf6c1b19a384c76cac9489162882a17f0d9ceadc197a5abd9c86ea90e7bb5a56f4e9e747fe69287db10d51480d35082a47e1c38646bbfb1bb72a7034668e7bf06bc5d55e4fad97d3c720635e72dfe6b8321304e5163a5cb849ac76a2f75f4a0939cb7360947b100eb51420ace227b4572b0dc9d108d0a46be32ae12701f7f5ca26b185cedd9b4c97f22f33039de467bf2e0b164f38b920a85c2ccf6b12c970fba2fea0244bf3335b2ce10ebe6b7fe65facabcf154141da66a6731b8ae30f5eb2caf7ce9cb9a83009a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha2efc703dafe5f6f195583b56ede6cbb7c1bcaa5c32530c4b1244862735800e6273a585f554c4a4a6df8ca38d53537de4bf4fda92ad983df1d42667520ad8989be64441a15ab08328930e81adb05d6dcbb24ed1a3c01ff5236f38d5f3dc3ff1b756b3f37f4d7d0cb41f78119f83bc9fb2de71eeb20467db2af78dd35a0979ae77eb0402aac1052ef976e6784cd719ff9321ca37319caab99bd5a2cd47c13350dd9d426f2a4f56f300807aeda195b5e45dc7afe2b4d579018c2a48e7f4e5d1acfbef2a155992aa370ce8b6792f56b673a47705a4c140797b5bd8b71c65627847e46a33af90661b67f6fc1441b9c5ae3ed36f66230ddded45e085497d063e0e046efb6263466e5ef1574c1af3173943543d0b4e00023d225553c888e458dcf1d1ba802fbc03a103cb2e2560c579515bc8e8b65a6f005d40a490cb025b9b13ea0079f59e92a8db9583d30553d365d9f346d4b81c6561a2dc25d33fe904d7260e3556550f293ac8b0731672acbae9237165ea463f251ece1291fa0c8c492314bc84b62ffaad739c45e353f96b49b274f02d922b1566c7f810748572838a365870916c07d3db6809c1a45f47bb69a7b3ffbd7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h50cc02d4c17bc1d3d3aca6a368b646eb81347854a156dff1b83def1311f3f88b9d39e491c799f3f4c23b105b8c9c5f29f687e55de40b2991bf268507471d53542681dd1eabc31dbeea00c47558af3350302e4e33b8fc166f7221ee956eec1c9f69dc8d76395f0ad955d49d81373b927e3091c5d1ba27ce8d9d63f23171a779e3c1403b1e56220ee494f14cd6f159a318c25162d54d494c517cbb831360a5a395929e9896bd434063ae92d93b16374c54b7e431f0f4aaa4a596622e4a8f343ba344d7b20089ec4c647d705047e87f950f0a87fe12c13e876fb22a1da56c21575dd7b9b5babe4d1ea8e2fb0dce6550c7d2ccaac0bb248f048f16efc85ed94a5d819c40a9b9200ec2d41d310a1c0974d022a0358dc10d54e899db6f036141ce0695a09213af3539f74d1fc42c89fd1f6a9bc097fb786b48b63baeaa2fafb1f20e1622b20fb7c91478483e48726a094229b539eea5fd79f95aef8b5846b33b33c4e799a58a279e53d8336997303e4883cef363a899e83ee225506f1c75a951a8032cfc1225581b290f02dfd6f7edb826d39ea76bee1a8ad090467e5f36a369b99d3a7cfe145750d6adfa33943b63f0800947;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9fc703e9feb6f26274052c78f8cb9d3a70f712c0243d17f93ad5dcf2db96df6d7c5a39a032a4a1eaf86670b09632d8dac758bd1d892779058d68dcd0f0e98c50f2db84526c1a171d486a31d8699d3fc663f8ec18caf2f26931b454904590b99ac17133e4339c7e1475cf85af7437456151dc059465b9d39391be86de7276b757bc51d8f0c0c9f7f1a900680ff5a6cbe4245bca223603849ba5825273c03945963d1ce02661fd7c3b16d96d1a35ed1f844dd64f0eb31c52b9c1321e3acaecf984b0363ef6c653edb57506340e88bb752489318f0db1e3c1bef9acb58542f97d608a59e8a59d2cfcd2c9ee6db2c8750f5936b05c7e12d0371d706ab36606bbfd2633d782c4b805eb921a05c2495c4022e885ff203cabed06567ac5e7d5454baff1f4d7f0e94993d93c0275fc87c878e581b4c24fc376bcedfe4620c9310b9437e9197ecd2b10d7dcd2f13b33b513bf73ab5abc3b6105131f7660994e0d7a109d4459cad24d8b9426ee64289227516bb729cfd2a4b5b2acdf1d0aab960f27fe68cae1c03f4022d15eb7163fa628b874eef299c69849625dad4684d70dc8450b99c17dbaeda8155db4ec8822d06a15ed6c00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7c00a1a43028a2a65a4f0597bf0b094d9119e0d036e6fd2e6923efd8dbc6f36a80b9f7187f36037e531db25c1b82d3f2b91bba033f436976409164a53a24fa7d5d97b21b8dc70ef1bff68a7064ede5f7fbdb95cec2cbcfec2fdf877e08e88ad0d423c16f1043c1716eecad303ae4fa78721d3882ddf5d812451f8fc557afeea41183adafb5b996324480d120fca66e004d74dad103b0c04c19dc5cbd5cd59fcddf0d685f65afc7783a7b7615e660fb9a8e4c6f8fcf41397a75e6f76e6153074678442385d7e22368cf172e0e4c70dfc49d0c8361fd636757ba08c39f7c4570685f624a9bace3a68d607c79d4c76daebb80fc3d49829027ecb64e96592a7f81cfb108d0b8209b93a858bed32ade25cb56debf2ef2a8eb6c8b0c29db8134eafd70e93c847ad1e2c01bf81bac6b2f9106f03b8fbed61adf105ab9f0ae51ab773156e31bb17d3c262d414b82c3223d2eb8638997bfe9432bfb99cb3da6eeb2b8bcbafb8326cd1cc8bc8982c0c73c80af71a539af62f0bc3b346b5bb826f282264bbfedca26773aebe51f22f83225d578e72da23e3966e6675a952ed2696003c74b4d180617fb56463f4915486e2571aee001;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdc1453e2d22e46ecff26754fb81b3210774fc5f72b2de028ac8b57ed794679566ab4cbb2461f5097db010e8a9e5559e8aa89257fc398f26ab923db1ff0c694aababf600ff05a321d164998c4884d7296f0de85f93b669ce2902181e3199beb257a78658416c4af28cad0a5ea0932f8e21aec6887caa872103e1c6e98f221900d5913904dd9e5103a17fe1a889c2a38302e6a0df45cb97f66a55d0a9693a45ebc8d69f23f0ebac3da7c67bf8a6e1be312dcd0aead2ef3e5d12d91a307435d43ef6a4557f48401aa86708633ad96f8aa78fd7a73601a3122aa3356535ff976ad86b8f17cea126b236d1ee706e860250e7fbc91e46feee24852c1fed9017e6b10a4b17442de4748e0b16be6c27f2e47db2df7233c64edc5bdbdcf7c61a45c1b0846ba401e41918750df66403704e37f32f755d1d9b8a8b364dcbe607268bd01f6b8c2dbb960e4220d6d1e3dcb631c75ccd80afa54bf069a741ff6d853826484df481d2b9edc7a66dd7627350ab5f48cb138d99ca8edaf06833fb89def977df949c5f6247abdd2e142ff0224843138619ffd7e47151d599cdf54ba341e863a6cd5436bb38c3e0034190cdfbd4a18d805734e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9f18dfb470475f795f1a6bf4d941d645c018c002d84e0c583897c2c31718c261b4870a9f92ffa7222401626b717573c3116c62d56766c91b4ea16d455e864aeda7a5313dd1bbd284d98b559f56180e96dad90e8abfe69596db4b485986a731d45e106ab69fc6659c152177f47f8b89dfee44885c62f476586c9bd9e169a7d73c384340a566dc8d6d898115e1a6a0f73d6863fddce3e0e78413c990513ee48e7c785ecc769a905c7a217d6ae08b1bac38acf8ff04182e7852111a7cabe2ea760248ba52fa8342437c7a7e91f9d1365b1ecef60c9783f3b40fec9eebaed170c872113775f524df12b0fd00e0262334dc6c445bc6a64156e4131843d16bda813bffdf9854ba03494721f19c70a1e32dac8781e1064c9f18b49a7ba6a53926c85bb24fdce866e4bb5f90c17e9ba5943e9fad13b77cc9c502a3569f7deb62518caa5977205050e262ac19c5969bb336d6ead53d8b35533ca640522bebfc35ff935dfccd6851d5465e0c07d14d7d8e9a8ede8d89b79bceeed377cea5e50f063a5753ffa6a530cfc65cded03f6f9980ffa8d278dc7cfd4f81e7b4167cecc905d52689513d521646d840550cf182027dbb150f26;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he5750c58c3302908848ace17d2727c9f3559524c7b0bb592c3df86cbbcfb2d78e5041f350a3f6d81bab7b4b98082d39903a56e8bfab3d9d1e9f826802a2a97c14e4e99cf9d8f9704378312fef8aecb4cfc7501a81b219b5892ee0dfc39837331f2292841d92a6aa256cabc8b29884156ceef68992aed0abeb5351be81e4c988db64b712e88a6edcb6a6421bedf9b5b192eddfc69165e4bb3d61d16e0c962759e464fd24bd7871cd4f0ec02ca14f0e8913c06c1b9ce068bbd18872217350b2b6652fe363307cafbd7cf4fbea2eb462aa35e461e772a07bdd7cb78e97a53fa23f87ec3c568667f804e459d9dc07ba2962b997bdfb78c8f7bdddc474936d9f5dec2a51a3eac2dc790a57a4838756688883c587395b47cfea87f1b2562d68a2eb43fc85364cc08ef8df93185a3a7f747127f557021f5d978613cd0f8df5afee5ec23e8f792b74ff0909cd1a3f0dacaeee0c56b640e5a852eae135712b27364dc1f816e9d7dd24033cea4a91ac9de6adbf0ec52ebed4eb146b4713b7a1b111da5ddf8a38c6ce4120d642dbef3299ea0b60b03d29e29f36e246ccc2fd9dc82aed9df601ed8c133b2531fa7427a0722373854c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he6b89b33b7a74832e17dc494c3a0d930356422082dce46a1585959098577a0defc15db590387447da428c394d5857674c6e18b055d26e822ea043354f5d70715bfef77db74a2c369fa50356a8d802da14e08884c954bf55160fa3e484922d485ae8acac9d37ea7d2be9a34a2f163a167e14a5be329397c31237d4ef8cd17dccbb939a567f476ea318012581caadca74eb7b35a97f9a102c5a232d4ad9a8f048d26ef4e9169a1a75318063831261062fdeaf2c8c66a54d10d1692de591a19947b56073e9050126fe56c3a4fc91eb46c1d778791b36694d07252b8d444fd33ef3f02b0181d313651455e3ade4003e632dd5b68343a6866f05e7226efa96f2b24aa3d2464541eafde65eb30c2624134e0f9db4ed6c8421ebad8b63350dfd61ad2fced175249827a2d15102c18665cd04af00717da0f20cbc2b80968fee4335fd40b9358b57f8b69ea25bc1d4a887d44bb516c4dd10243612f887b328f014e256b22d06fe963eb00ca4ad55cf9de1b037e703073061dc5fdb53727175497c12d8ba2fee900f86d803e91a2d5607b50e78a7fa1eb226e9bbd707aa6025f5bfada07c2fca98db8daceebfb1caa46d89f6ce253;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8da0bed7ab5d23102e5c8b2e1607f49d3ba2e4a13871a058879afd419d53c6c2e7a649c63d44e66d7fcf9655ceee5ec564cd54a53443999c85326d9ef76281dda2d1e117de440705ab7cbe5fe2a0d84beffd746b2b4c9e2f265751ff5860d29fdec12fce7ec0ee94722e36cac31f3298651e4d891f650919296d3b16b428340560eb8e567c48409c2cfe020ca58aa7ab90e07c2993b0c7f856ff7b6f75245dc928572f6726587a516b4b82ed18ba5183bfce873d298c37856fa25cbd5740a2634ddcd095939e6983ede0dda50e1a2d5ab8182b60d7e05e3fcf2fe8a396324b2d2da2d87680ad3cdc2e03534709d1b9b328f6d053280e463eb036b52a957a6de2a56f65272352ed49c2a4ca0bd7d74eb57e33f186feb65969cc95492c2cfa307cb03e78fb4e4eebe205f897b5a6df9cc5da8bb17f84f4bbb36da1e6b736d9cfa781f8e54fe9f986e1fc52f92d79375759fc65fca4fed45a613330ba1e20ce2335051ecd8d1c14569e1937f79dc8a56e5a7ee1b0a6391fa66e4f1462b9bc65aa2da985066b3502f001dfbab51f9355ee867156a96e33c55cc80b9b64e3291ff68103980dd2765c07b4a5591ac9d70e6e36;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha3de7384d994ba6c6ea847c079b792d85f004e2d3e6fe05e0600b8650285be82c7777d8a7f3b8f6541f887cb98e706b94434a5bb58d8e9ac7f30d437fcf09d063f5d0252459b75e8410f00db86d623d4d73f3a54b43fdf1f26d992bd096587cd981c3fc14b18d412d6c27af21d8be6eca54d3c469433033803e2f59614a99fe00eae05e72c451b0bd84373d0b3761ed7e785c0889b57058cb3318c892ead7c2611d02bbf5335f48b377f97b8f82f6caf21e6a19783c2883bfebcc702bb8c382a7b73645b338621d03f74404623a33a7866f8c7189efb90d7a9e880518447e36614a2d24e785e8b00ac2876db7d17d7d68abb2fa7d990029b56f0f6d711ac78fd02d4a3170b4a214f7a1081df67720d3109c7a19ea89f9821e5b1a5374f9e902b292be7f06ad53a6e92f820d6ef37f5f4d1c4f84b4a3f5ba1621a3698e42eceb792c0c8c7224c8614f9ef2d78207a677c69cd59add88e8f92877b361f53f562779fc17e1baf1211e645abe2f46c733d6372d1531329974772a6a7ef572e1986fd1b0099814ef2c7d42edaea9c4010ed0a4ef02eb946061d26117251d987562d3f106ab72db5d2814e17d107e7d03a1abd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha5c330da9f021bf726a8a4df5fd189ebb07f4d606cba8fa67a238fff0508bc604e6144eb84cc20909577a0aa519ad8d20e95203c771be272e131a69353973234d473a9a9d1553455e91a5e2f48b91dffa8d173cbef0f35850d4013d8849fd017f5726d1e36d5cee8dd64ce15ea3bc160a7043857c123af2cf8896c7cecd2f9c871ad5a8128509e593a60096ad40a39b754f0e9ccceca88b3c3f77dad26528cee28d56de51d114daf573b649f12464b728c979a24571cee90d736108e338e01f65119b7c71b3eee422c72edeee241e69e073245788cab1466517470c59d389db051abb8fab6a0a58a8cada296f9a7a35e5019360798489bc742a97a3283bee3926db7d63860dfcce9a6bac3d2f396bdd09f5021cfa62b2a2e4ce9fd74a96964296cd4152a7b29f5fd8366301232fdfd3f850e0d3f70ce2997ed693d0f295a73da1d8ea27c51e82fb76ef7d201bef30352d807674f2e584e8e4353ba3dfe06d4da9f9ae21fa6dd00ff4a9bbab5b0773bd6dc97f55e041c823ffebb67c18e297be80671a907fce9aae2d135dc490d9798bc928dad698fdde7fa3b929916607cc24ff1461c388a7fc12edb8edc8457f501da;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd319bb5dce0df933e35c2ea7de143305e5f77b824ea38dbfc4e2804fbae85d6ca6c14db0a7f28df8ca61614c5466cb59b13bec28dc76cf723f893b12c3929600f1b22c92077ba80317a075b9fd65cf316182c97fecc5c89c75f39560aa36f376b9bfaf254676eab482964900158adeb3bf79ec92c8a7a00d7b3742cf5d325f3b91e548c19d42d0ef4fd5f2b7c485aefd9bdcefe020d193a61e63000037f07e9c5eb004b20f77c829f72dfa0b868a51438fabf0270c770b273c13a9f181411c3b6a4d53928b752a8de9456de27ea50b1919fb7608c386c3b965fbd0ff6751c02d1392366e21999752fbd0f3ed63db5d7fe856891a4ff59785b02267d3f19120b696c49bbde5812a5df61991a15f669958888e08215a817c51b644ec116995b4222fe1406064f55ec2404391de0c310ee95b013656d9b32c1e48969e5e49d51fefc5aa7713cfd57ae6d596940d42955eeebddaba4d0b50ad7862b6337ef3c6ed81a9b9ea0c68f58bb401c5e570d840f36e9eb8b695e383ea52cde627bb736e401fd180507a1b0d95e29d52c6e85a685a7ee2e57ad75e2262930167494c5470fe372684481dbaf5e21e92df6c3e638ed1ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfc50c001a62f96e9863c246881098fada132924074c6769a9517b0f77c0a327881a343b8b301f69a70d0d12b0131f1bfd68f36e4656fb23c5fc599f9f13e3717bf6898d6fc96b51f920c6be5fea0860a4b10fb7a730f75c84213a05eda37e7a781148cb93363d1cb524e577580071e8f00b0e528e8e752dabed7a6e6bdd4a9e0e627b046a69179b9e5f2b83c7b251db750d471f50e9efdf0948463b5055968926ecb591d0755d931abca779f3d978c457789ecfe03f9418aca368f973b5e264c03c4d396718a1e385068291cd5d6b0f32e3ec9e0a976f67f2d6f73eaba3270f0f8d22923a249d131ec02620ec09e2d8230d7516ed2166ffa8a429ceee46de2bff91f1b0f5c5abba24dc71314bf9d7f999d66aecab29a511e456f9ae2e810e826d867dc1c48cb1a2e28ab733a99b1d6e140c191378c98ae7b2e50017e7938e62f05d5a85b444bda14146c1dd13d0a0efadba221e75995aed6e91692cd105c64be84d40764c5bfb7a3bbe45d8ed30fba6e882c6b8e5c2546f280502703bb1a47e2a823dec79895dafc21e221c4261e81080859a2f01413819dcb0e314a7dfd5bf080269b8a24e83d74339cb57c60935f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8953303a58f0cd674ccb2f7479e492b9e4159dfd989c686995407a93391dad7c24506dfd5b4d67ef5934d89981e635c280762379f9bfb81fe206e9ce999daab1a7e84724e04f304ed8f43d616a196726c69183cb7aed0e5caf26d7db1022abf680c835bd35dd951d6eb6ac055be0b73ed9fde11ea0c88c79bc1678819d0eb06da28f851320bc2c1390414aa2728f6f9125d3a7ecf0874a2f8871e9a6bda620caa328e00f532b90aafb6e9a2b9a2bf46eaf3b169208a227ddfeda6e9bea17cf8d7222c532b77499c13f207331c8b097678e565ae5e9a309bf923e9f9766b1dac3f69fadb970a2c72ec4fdfbb0ad35ee85dc15c3ee68d32dca7f9b4c44623741339c04393a10ca571cb5ddec5edde99318a28cd73daba892bab2b2dbb029200b14f736957dae4dab4187b43abd3465601c0e73e895e86cb197b620e7dc4bf36e1ddda8dc3b2d098d4e6fbab691c41033a55f4e66957bffa2a17ca89f1563284ee3d0df885d9ee769e418a27f0c452ab5e025877bc5897f623f12c1f4508cbe5bc2ac62667cc7a1420ce30137b07a0a39c98c64027ea1d3e79cefd5d027a2de5eaa4c69d975f202fda0bd66c7dbe9e12044;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h287f291c936472d55e4b651325f5becec2e5147a1927ae3155e1f2a05eb81b607cfe3b9409fee9883f9c4aad1f6873c9fcdda4874affd524fd38588fc78bbbd4de89de52bcfabb5d2b508c13e72c103211317ba8e98db93febd4da3df861ef49727482324814a1ada07af6e77645e01adb0db124e6e0012e049c3b32797ceb99484c00734b0a3bbea9622c9b7a23ec95aa6289d2df90594447aa96d896d015cf7471aa6adade9ab5905bf9c33af406d7e3b2707f809d60498dbcda006a05b1ee1eaa6b6082d62af5deebc71a1fa5b6a3694b3d1690a7ba58550b37ae9374f40c2af1d0fe6b3423792ad5a79f538ff845ba9d91cb765e4e8a4b240af0a8ca38d338a3664e33d497a9990101cb41ecbc615a125ca8154bcd3d7a5176776ae20b9b2b2a2c3917279d7cd105c358a6f6b5c858815a2cdb8d69b49021610c75db45d78440c3e24c4406c847593590fa45e0e7a55aff3d20749fb0225ce6307eee071b7fff0ed6d082e909dc995880cb85f167989561e6242b0d506b60e0270ff84d0675814cb680bfe92e18a12e779147fa94c0d19760a4402549a4d8a6ceeb30fc9f3ee5481d771e3dfcd781b79a2d3f0181;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb74e63478fdfc08d049a74dded7062ea5fd5fb118d184d97b36a1a86f4911f7bff441324b75b7d0cd8a9d966af5a131526d02a336e0654d55d94832f01c4f3a7d57c46871f0929448fe7a1c0666b8bc644f1275b64d6950c8c1fbfb2dcb86ff370396152f688252f6aebe119e1dbb3ace77ed6f7a1552f7958fb59425fb57b231abf7d9fe508d671acab43bf3b09a181d95f69e4b0500916d4a2d4ec25ad96b684f2a9a7dc414198d0e6ac7510c8486cd5dc2694d940cd85986819d152310c3f38375261d10ad893601b4aa433a9240b60c80067ab27de36a8c7ded90fdad137bc7e39a2a873b141305b3eb1a09bef22ec7a2cffc2052021910ca5140e2be97eab9e81db8ead57b8e7756d3a038f218844e2eadd598549119bec9a14cc54877223821d37c5cde5177f62ba7ec14712bbd89452439ab13da3f6b10f419d299031ec359376d719aac1e63d4225b58246798582e35b23d9d70c9f5563572fc46396d76604dcbdfd73e8890d64ebc9f7abca4f3829c50be3d53324d7d13b208568e63d23219f0db4bc94aaa2a325fd98e8ef0b731488844c185773a9ce59d47128db88a1e28316951e8f8be437afc60538d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd4c477cfbbbf22e20ee5cfe9553b180163adaf9ca27045c2073752643a22fc8cb6bc75157500ee9045af9528d16c421a1d9d29f415095fa19e57241e16bee73cd77f774ea518f47e7d53dd912916cb008af7930c83f9dfd4ebd888774710e72c792cb634f4f3238477b96d844c0e0c836fe1c5b91a397b01503793033171acb18d01b6655691df9c7ad3923bd40bbb173395a6dc82bc5803baafe994a5fcf2d9519f7c80e52b4e25c174e9e6bef4bf38ccb7ec29fd6cc474d8281000760fd99f324e0a229c90c44977d20d84c0cbc6bcde972af4202a93a2a7651d07ffc9701d1f53ab46dedfdc7481129cc3f9ede667b4d7cfd8b0254d952c07b47d301481b801091830c7b291d92c5f134a2af5769f66ae9edc44fd697a916d228e8afbb072bb33f8d3f4f28f9734a3412d8c618fe637ac5c2e3afc1e9a97a6513265b6dfc141cb3af3170a957eb3a8cba8fe45eabdf98c61f0795d2648768f81baa168fb968c3e5e267d296a7f93938de06998b76b8978a010be04049cb6b2742c57a7a4380df25822cb5127ef8752501b069c5d6a74fd207dbecf1ef51d4bd73e799ef0838075ce28ce84dcee5c93bddb40c55304;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2560d8290ba383a1caf0cde3b62975588dd5beff3c7475912419282e12c5d8912bbf7558110a3f39761fc9c37c9ade92db369b5ce60da3e0fb5a618a734fe4e466b947c3ce8df37024e4ee6f842a6ee2d7c46784bdd442a5eb3b5099f5ebe99f09140a1d3eae7e73b5c9febabafaef812fe7eec6c328cf2cce3d51e0f1a234d4d8ac13c1f359790a8006436a4206ca937370da7f2e8a34346484d48a84480326d1a2b2f8eb9c431644371d2d8dea7c746905d0699d78f9836261b3785c896dcc48b2af5b5b20ba721c1415001f5706bbe06982a193a0c301a184fa83bf666c4891694b2dd0cfaa08fffbe4f6e2df861289f03fd562c7c7f857c853e028b51ddcab919aa154e990d9f39838599b8aa578fb6ce21731a53ef1bce4df43fd55ff334f2920fc6ea9e648ad1470aa4420b1d7c17de07e0bf3a5af6c453ff03b971d9b47d4080e6077d21312ab82026314c2210997d10478f72b251eaee39a12f6452a163a2070d64417e251b0aa7f9fdcd8a3ec0540d654db30f007c54fc4264e9415610a9427410017a20cea4be47b1159785b8b11974401ed391f1bb8c2fd60238f3a3eeacffef1e2a7c42a6246bd859db7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha11116c3986052335d04d213dadf9a2eaeb62bbae57186a1aa5ccc3dcce48feaa3a2e6d44893ffeadc9a900b0dfa8d72300c619b6652102a8a392c1de2c4fc8579cc8793e81725f7dee112aeafd3f77be0140cc6b4a74a686104131f00b59ccce44cf6b682fbcd5eec8d535ada4f138c2c9b2ca99ebcc2b54d4e2ce55f2f0b9ecdc82953e282b6da0530fc9e0c60f0cf06eca0a415db8c2c949370e825df9b7fa62d8e0b67322fca8f230b76e9504a2c3ae6564280aa6bda08d750bb7dad162ff003e1a27dc2300be06e2c38b6441ba5c47eb095ef1bb43a647ee71e39f31ec7479d4345d8ed26d38f46c25c801310e5cea357b53f60173759b0e8786fd9f91ac9f075cddd009a9a4bca1fc0fd1b5df799cd38554356bbc5d6c7019ae0771885536ef6cbb3fa54f0f5f89b7443f84ce3aeae27bed1c863e79311d7ebfbe338667ed6470e6fe2cc7e4266275d72818d0bec812caf5d27ffa0908a1e84ca4416277b620a855506412361c1dffae643df06585fd70cc2a8c87684d84e4fd9ec893709771ec72c455b52f465003dfc67996abdb5203fa0aba02caf262d79a00978ae03ddccc1d01ca0e4f3f1f88639f05233;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9e2d325d3cd2446fd3dd6043fbb1236a8da19a2a9ede0e34536852ad7bd72c1e367c27008d51dce4f9b727512bca5a14a72904d1f5cc60e2d0a96521390176d6425d2d8feb9e6587d0dc8d2779131d26c9e771f1fad7b6b53f9ec97ac8950ba54cda729538422309b48cf822e151f890ee9319c4a5eb280b4a2b4b55524767605c3dbb2eb17695ead0a993f9cffa2ffb1f7a120c2610caa142cb33fe15debcd553e6a05ac28adf37e42180bb35dfed7db29c1cddaad63612acdfeb1b28b69d8b104b4d0574a0d6c6f8aa411b3e15125e42d6be5444a659d84913d1c5e7a52f2dd6ab9095c04388870ac47953464f887ca6ad0adbf088230f0bd2621f56b15c0df348c4c7716adad94f1fdb00880f16b28c3d0e0c5eae9d245a8c14522ed2d9d96799564bfaff0dd60be2abfba112bd6cfe0fe8b084c0e312c1501509136124c44e91012e6ec91abb4c8a90e770db61cbb700f6b778c4724fa4a13af054f49548fc4c7965782a4fdd4052efd3947f4fd331f85a3f2903e2db7e5e2efd784b636a3c253456e44d213f9547e51784a5f059f1676483f9c936543e83c45da7a6332b441d35917b95267a3584ac08a6f4f538;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h430d8e87f54ca0ff3a77945308d4892bc592813925a234656c16d1d82b0822b63e767c1c4f213da14caf929771b886aec72b71316b5ac677e9a2dab841e61f5df8b0af539ee54945af6a080945b12429d71c2f115a5ae32d326cecf733b3f27c87c6f1eae7cbf0d0e87a22957c4ba67c53465747bae6ce29f104f46d1ffdccd8d8432256f5f6005b9b1dd2c0df5f761b8e5dc0ff66a5ff81a6257c06a073f33d1f6f3b997e15e374d34b88effbe3b4f5c9a3b315a13c5ec9deb80602178e56b988a3d8ed0ce6e7189060cede26b833532195e24c95f564934c3719df1c43b896539abf11154a02a240f1da1412541cdd72587d2b795193ee693b653601abf81fe38ff0e755a7fe816fead3062515fd6cf3be64b383de2d921263c416b2bd4f5764e6d52c29024f2f8d52b762b2471f4a8c84794643437b7cf3b2160e3e0b25c9db5e8735c60b00eff65e421a13d1a5342f8dfc1d57b4478a61818cb025f4a1d0b015a9bc414e5a404dc2b3b8cc8aed7551e9d2331a690b97645e9739d06425daf5376be7676f3fca7ee5c5387fcbae98c9693af983058e6bdf9cbf941f19f1acb74b55415c05ebb4ef67f88f8339757;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd387bd56483a795d6bb8fb17dfa49bc874cd9865cf3ff7bd4b92694b134a29400e4c1469855bee6e4893c463d1d23a6a5d073629cbec70cddee918b5ae2453f2e0dd2b0898ba01d887300c84363c74185fea39a0a61c7682ce1dda6994ad36e59d41b7cca216a7c9fd1a3866aadc0a7cdf4fe4ffa1a2085eb5cd791aa246acfb08eb2f062e93add95f5f0f7d32346bc58a687090e6729bf3b0d400554be15da5cd3d03b92b8d3d5ce2f1e72986e33bf92abc8bc04536a9f52667b8391d01f70e65fa47e03ddf67786b5881274640d0e20949f26261a16bca8d57983f333aa6efd7b6af8caa4a848577961c1a487d6c5695d9416fc7dc3523b37d6c7805b03686cd3292f388c94b90e19ba7b4e06bc695d284cbd649529871fa0c1b49b56ceb46b9a1c37baaac25e29eed6c7e20da532d3d7292d4df3a56327e42e34185d44bb41dd442162fc6c57b1b1b7f908cc513c8f62c7f6293e5117fce8975ab7ad389f184cb5bb6e592e4bb0d3691b11d8bda212dd4be6c2ce77d6a766266a43529746c2e5e2e4452e00db009f189550703749a80a43f8d4a2bc29c78a40b787ecd80ea41568cd1c80daba2a0df85e0b344e180;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9f7fbfd771ab74fe590da6c7553b988b2bf7fb41a6130da252817cec87130f43326b848418faec77eb8cb369bd60dee3c4f63898a675101d57f0c8b455fdc97cf464a5c9ed4224dcba6d022ea8f6b0401644341afa9f03a4226bad552179bd80bb935e292d69a33b8efb246bf4ed9f374acaac2511c581d2275071f403bdb44cc9bf36a5d9239f45417eef70e62cbedd7cf3f424e99f135ff10f4d57debd57a1aa0150e6d8702a73dc326af2dd7a2866a61f0c8d42ccce815567b2096cbbce9ff2b3106fa6d05df63f78c9fc83e35b2ddd8ff99ff098d802dd16124669b4105e8b699721d66a5d3e1fbb958d1f1240be1dc310ef10ef8ac2e7d01dc028d663538b2afa212d0cded636349413ed486d4962a50dd3fb1022635065f3feb9c0f8c9c048c2e958f83f2c0b7786b3df3eff323a274663b9e0b8b51658b5a0b74ff3249197d0a38ba4b615bb32cffdc8813ae9af33f9838cbad11fc8766e4b99d2f4ec192724c0089b5a580f533781a771e3320d1af9a4948711f160a59c761808d5d4f54e13a5fa8f81bfd9c94434d4c195494e4cbf611f66d6e0ee0579dff7dce9b1d582c8bf0c4456e981f8b9e4998c9de3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc6df71b82ac1fc2e3d944b4584ce0a185836d036d1656bea48adbdab51b2feb7f7e025a080bfb84bf39734486d1605405790f82a48dd501f59432e7d34f7a7427cb6098e95c5170020167b1e138c0e9aa1b3d135f1de3290d3d6c950b1894894d5af1da5267e92ca1dfbaaeb66ca5756a1cc59d2393cd619bab85e3521023d2dcdb298e1c5fe5b4942ba49a798fa9c04e24454b0d901d227b37e07474baf7f2438f3aac1e2153a49c889a8164a580bda2349b79b3ac2ba09a21c83f9ab3514fe2692ddbdf6ec5d64735612c18bf883644b8a66966d9aa2a77a9a988b78e8826b9c2d78ba1393678227a24d03a0280aea64ff0e68e34cfd3bc25ba3d2cc3c52af3c134ebfc6c125a253026a26f59df2bb8ad03dc827999df11fb5b2562ecf744d657bb86a94b374ccaf1306447e79e1499faba9c456c4484dd7baae1b50d12c8acc4ee3e835ec96eaeafdf24247232732c3fc77f5867efb43418e7a934226973036aeca856d0e238ac8b8893a489675c1bbbdd2cc6c1f07f2abcbd452755a710264e51219a0b614aa9c1b965768539c517fd2e9cc593c22a3e600c4adfdd48dde9330e779c6bc169f135c6bc3d35f72cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h152f1f0187632b01071688c6d3342d4eba75f8e5be527901dd6f99d45b1c4e299ef4212ee926744c6862cae3dcf138b6189ec0f3f585acbf501f57ff52ae02e58831a1979ba127475c8a6d5666798543055b3ea6b301ab10cd83afbc4701c74d2324747dcce9d724e6fad66011e1bfa72e820c04ec258ef2f03da2bc17fce52cad2bfa06e6d687daeee9a3ed38b082b254219636f5ec975886f56eb92d8c1dbe82d3e985f48d739cc34b6589a255a2afeb5ad9d428ff15eeea695617747e0437c32846799a40d87a9220e4d77dc89ee0107c359b22fbba2a726a41f2778e80605867b0aa9769f2471054838d51691522f47bc48b76600005725b3bf8149eb524869f2b879b30098f763bcf7782b2dcb52be3973be157e4b10dae7e6320820cb9e5a2739a613985e1952b4abbaae769c1cb1a6336b8bfab4c63da1d03fb6901b8424b1e454f87e9c50828a394318a2ef443ece6a512c43d1005300928d3b70356b94924728f31048d81bd11fb8aaef24b8b6d7ff08c87ea8f02346e75a9118f0efe7bd319b5d15f19bba621561311bc8b8793a02a8dfbe15f145beae95bc62a631c6b9f157e745122351610b243a078fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb2c2bef5945d0348ba30b32d395d8cbe3bef39a78647d9c76a4d55be6099f2e367f994c2958360693e66f0b0e6c1dd9a84ca5200707a47e11021afdfdf5b9255c50fe145f6483c1be38d018d8e632902dfa1d4849ae72284cd726f84a43a5c2d595b293134305f62beca2327fa4cb6af565dd534b8b82621ad2b9fb848f3650dd91f691c2eb055989a7a97cc4ab341df96f78288df99293aaed8bc81cb1001c1ede7d8bb215aaa2f6c70fc19cb60dc94afa67f5057c077aa9f6fe586f6cf96e65cd881f34431f73de77b41a295c405a18e2b701c77b1416a452bab19dd7bd32cd5c86d4e5b445c0b59889c09071fd3a595ac2ebbe22e6737e493fc6b7bc8191b2d78415ce71b3470d1f77b1c13f808eed2890a017660728092d32112d3b9060bcd5013a76ae2303106fe79892328a5127a30fed01fa4c26f1f684bdcf7bea11b32ec963350d28224d2bb261a583e10446a7bc1b535366fe87c3a30437f07e7fc0e5cf77e3850c922aed2711ab84945276567352545280784bc6c44f421b321facdaee882f19e77f4609f3cac5184532d6cdc49f626a5d826bef1ce1d9349f4d66b71cd77d31274b01b5c1e20b2f475aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h339f0982dfa886aa25b6790f6d68343594c5deb2e725a33ccdaa767b3b60177f1fc3c10c8c22042bda5657a23dca1b797384a1bc5ee80e005d77fd4bd93865f364deeddcdf2d2274f8ca2145316bef9819c0f774b7c33694e807cab1d613371abe88a2f6a5c7e1cfccf3791bfb36126e4eb8d2f8c2d25ec91be3746bd0fda833add35af809bd0fe471ba15cadb0cdfcbdc19685e0646a7806d64f8f1b52242617ce98ed4ce6bf17690f52fd4bfb5f6daf53cf9cd02dfa82be0a707f021a47c5eff8648c698618b9b7129a4fa4787ca56f2645eff86c89e8b1d7077ddd85c3c64812396d9326bfccbc92b9a3dfb46abb1bb9f6110734b568577a5300ec97c2b447db5347c849950bce829d8fc1bb329f09ae3649e9d4bb868ec72adf21284fe104ca4047fb812406b4b12b728ad215cdd706d30edfc3247d76c98fac40b3a67383807fa58d27b8ca9596c6073878b1f7c2be5942afdd78a3d8b23e20a22f76126911a9f7e86c97aa5cc8fa4a09383f6e0198f3f942f7d2d37dd560d66d557f57ed39482cf7f4d41f9e991619f5d44983ca4be69b075a1444dcb5b1d22f2b20eb12edd6ce2238afe4a34d2ee6e32687aaa;
        #1
        $finish();
    end
endmodule
