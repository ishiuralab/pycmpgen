module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9249185dc231e8536746d14e9bd3626ac7b085a4739e69c24bb2520aba986593;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b22edfbd180de4999fce59b68e9a11aec96a3fc5cadafe9b596dcd3af233986;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3f58ffb9d21a3835e76aa939e9be36d4961c4ecb00edc33a2e533a2acf260ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42a3636c7ffacd807d9aa3490b6fe69ac9d84439bb6d14998d923da86cbd59e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h968632867b9aebf7dd299090d82e32312c922cd7e42ea9d2c99cbd1a62fd654b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69882ccf9136c52d7158ba4b933fef9b2e3c58395e0670a3262b698b3504574;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe882f2d5245b8e1a821d8d20c31dfcdc98856a5b3d2c98c2198627447dd1c30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7c043f6d5e98dadb6753bd190aaea8766943469de57cdeddf3e518e775f9c2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h680391371347d50d3490616c2e96fcda5731ea6508925a4e848eb5ea2f2e5c35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h879cd448c74c2783640c7cda4fb14911f6079636adca920f953cc2af9438fb92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5ed911c3909c303dd7f6116fea16131ecd4627a7d015f5ea9e6bb5823ee6bdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h646490c676de486212a8a9aa9a44da1becff34f4e413c8544ad74be420363713;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66b0c5c777347f0be61226dfd45fa7ea4155880521de3e775d8dd1a0261e0271;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7af0acf25d9e27590560ecbeaaf37c89d4c12ebcf1392e132ca281fa422b91d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28bbd87a82bcb20c2005a8858ed581dbda13a9356d6a5d50cd22a95a57c08828;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f9ebd97581844c2f2cec5c1582df8389f109fcb4d6763178ef57d0f1b86e67b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45612ae16b21ca7a6e15f0631e3328882d2d068edf1bcee00d7eb16d07113f3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ca4025640cbd1b5cb9e94abeb8460933ca7b9d501fc540cee8a98ddaa52857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1eeac1ac056f6dc879967c7faa48cb12c9392ba138cd884d03449e376e91c8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85609b9b7f454812fb9cea03fc58f1fb8e434be1463220514d958b13e0198878;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ff26135085237bf99af4616ea10c223f8af7ee4941be46f9d2fb62b8ef7b362;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha82ee9cc3d000ea7cc87547397a2d10a87435abdf35229b071f777194a6df491;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde32b6e2d8805ef7798080c23bed3da8080de86e05590e2518eebf89ee653047;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fcf54126275db1ec7eaf382f30b921276ab51e25b6a421612e38a45710ee009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52d241571cbb9e7615d0b0f2e8257741685fa9fc8ee87afe2e6989d39fffdb0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77dc28d2ae4516343dc24bb0ba62f2d096acb6e41b8d1c9432f5befdc1fb845b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b041cfe995d2fcff4ed854c449fdb35d23bff6f4be6b53dafc7b5a3672dc59a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa6c2bb0454149a22775b392c351bcabb11fe402b92c81eac27d6f86694e1f59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h497cd3d46127ad9c1e2181f6e80685fd10479bf65128d8aca5348cec15ab25c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b4345a018a83e0124b607353ea76163a2aca4fa0c6c27c185e0420917c5f3a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8905b5296082a33d5c67e0dbee0c51c8c9bf0456100971749d9d04ee85e30c40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed46ddc7f5e6c14e2698f3ac2a1b372005795b7b42fd96e60750038e6c18e669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf47229380ee6db98c24547a5c27ccd7be4a58e137eb72e89f9233d62b820af4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h361db4d2332a8200f75fc6431c6579ae3c66f29f069dc0b86e376d569f2d933a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8687f095795e511b500a404b1c40917f21872843a03f1b595e1373aed0f3136;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8634ed5ae0cba216051c1044ebaf14156378e545c2c7b2780ae75fbb7abd2995;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h648668ea17701f0e8021b126017573de09911f321b93ecb7a8b2b9db4a543a7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had591abc39bc56e1a12901c14b9214daaf3b67c3104977dc8f5080227416855e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26e0b348c3b441910d5f09c7318e78d347d69766e4fe643d44f0846222d884c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ea39927edde14f6a83bb6fb6a004ae5e31841ad400bcc4b200bfb8d28f2d0d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35f8a8992967183655c8d69212c85b34d82ee8d32a0499de844302157891f75d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2465986c6307813066c32d44c4be48a12ece911cd76d126516326b48024791f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccfa95ff77ea87bc2de81c9abb127d51c637b80533351ebb27ec52aa78808b5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41d1a08f7ca1270760709fda1b0f04f124579bb69bbc63fbbf3d48108765ba6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccfe9a56c8e0ca42a34e00b9261b444dd564f3af19c8877b14a27622697f74ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb457c9b03622dd0785eaaa3df168d208a4b4ba709286ab981277009e935a3330;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42e6ce5c4ce5f7923107e793feb095c664a4540be16971567e209967854284fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h373482f8d93d18e30c5ad3d81b9164b44ad1f237dc896389491c9ae8421fd43a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83e9ea44dd122166de8d282d2e5eff0c10d721bd4f23d3bbee0ddbee857bfe96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h814fb3cec56ffc0a0cdeb044e5e23ca1878bb493a09be4f008a7c9cd5d31a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7f6794fd7f2a4f384a5970bc3d1428bb8cea7b7509bbf5711ef4ed97d6e6b20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf411bc5c05bdcaa4b3e42363283d9b00fe96d8558a18ee75de0704ece2d2cb1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9603e47be11cedea67f43fa61586f65639aaa0825d0ffebbe2b5241953a96ec1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a3dcc75b807ca21812b07c2ac99ac7011905ea77258af3f5262247f0692947b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb43f0284050db8878fe02a0d430c504ff8dd51a4163ef91be7b504d39c8a07db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72f646e8d2f8093d3899dca7c4b04ffc43999092fdb1fe7a04e9429c70132f80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h478b51087f30de84e0cf8e318a5ed4a2a0c22a88105eebb3258009a5dc037b77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7fcc1fa93cf514cc06ab430c3f9271eed1c9c4badd613ed1c2b664fe298543c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f7f902480ceeb32f5adfa3c9e28e433e842f0a396db943da73ec259d1092998;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7813ba48c9af2692a283334b20970a9c2e4bdc97cb33a07d095142154d3a6e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h133427ff1d7b0a64ffeccfcba29abcf95781cbdd44b0bd26e7a23e2cc73edd56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he62855dc90f82e9f757e84a2054c60589d0f2f9555830a64d480f8e4dd7f8e96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h365bcc3d9a0ebb5f694a110833b9e19d5e8cf23521b2441921b5db264b1af17b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60db3e16691ec06a12fbf45451281ee056aaeb427d8b57e65d7c94a6e13de9fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd41cb93b4b8e0f1ad7493cba1ddf73ac0f6528a230a4eb7068a309ed08009e3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e6dec5493db1982f8dc7d8836a841f8c28c9deb22f269719156777e4b5cc1d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89b2415fb2b285a3d4588acef3efec169c589c15fa90b6b42b311ab5cb5da0e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c4b6cca41c351dc63c57c1394bb9cd05552a64d4933ae5f6f66b3bae43e6e0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha583248c5d35b7755fba0064170cfeea61c937de96e432900c4d55caab3a42df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5578340ffd75826d9791edaf7b9ae6edb2b256def608ea09d7f79c1a955fc5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10474eef756469231717da275d5deae5b46f9a5dd60bca62b78391034124ecfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e84ae4320de2dc6f8342a67919ae50ea53262bc4dd6321b393337a7734f8cf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba491660d60d6737c7fa3bc881f6cd31b76821a5e326f3f3f10942d3d105ebd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fd930c31d29beac969fb58c1094e7ec77c43ad151e7525507861c7b187f9319;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha91171d0646d9a7d0088be9e2495a2b629569ca1d2bd92982009fbdeb271334d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25650dce92e81d787f95d955fb4ca74a92005839aed47ec93bc5740524cb6b72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25eb298a4186983b8c0c1deb1263a3a7819d89df0b9dfb19eec3131fa0e8b2b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0d5e507b701fb0534a10b5ba221cb0c16b752c5ccb3b2213c219af85b1dd1ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1604d49d2a492178123071e31e3f3cebdc07fccee5211e3a6f071e91ba35670c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96ec28e348145ff88e795de93cd00cc8aa2f2b04c45424094a1692a7354aca02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4932cc82ff7b416758e61a9714a7f06450d42e95f6da021b036b294b4adc51d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbe269ab930f8211e7b07deccdf4fc3809603104cb1b2b77b777964cff1b278c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80410817b4544c980828cc2c527e90343d56b5c026d8d41ab856154ff9c33a74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3d065790e4e67d3a29d469fa4e2aac33261adad10dd7b09ec54829c18fb7531;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b3ee04d5b82ed93b2a5b331298b00bd269600ace823f4dfb5ea6ef879afe14a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca27d4467f851f3531fc12394056a9dda3e372a98dff99c74fcb8559e7dc3c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc110b9ef946b553e59c283cb39bf2919d7211cbdc4e3856a305dc1612010bb69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h287df63c6b0927537843b9335a18b6083774166d2793de3f46af460f165183fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28b6649b3638acad2459e29126763df9eff57ae08f0b4b1145c61dd18b06758c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf19e2819835cd06a2a141de253de6eb40038ab0eb6188c9a0196f04ee65bac01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbabba32ed74424e96db65bf20c6fe77f7b589ef28972d714f5e60b3acf0d2ce9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60440fa66e303fc86377b8b522856cd5a9a3b3c409100c1486e18288f559501a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37553080d0d81a564bd87ae018665e49b146bc38a7b814d3d494800d93467dc6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h758560901fe974624988327a1dc417c0e620811bbae734beabd4da9ecf087cee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he905c06e42dab55a9610bb0c21dac8fb887f0e15c3687598c0693bd2201d3a84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2af635a88e582a140afd6188dd8353247c71eab9d6e37a29fa872024c40799f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6c5c4bb45eff3b0cd0a3d0e277c7630bb04d4753912fc4fcd8af20577b22d3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaa167ba8e3487177e15b29e5b96387ced95e298bb762ae812923c6da81fc2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8dfbdf7fd4c476656baac5974bad792aae626b1f40dfd4cfdfb7c45b1584c6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefe5406eb89cf54d7b0f3947777218a24c579c135466f02d585b8887e8d042ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54dd47e69eebf43e17069731d15ce86bada5669c7546b756b77e56172d54dd50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c79214fdebeee558121ea74efad247ebc8603b55aeb7b4cc7166565cee88cf0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcc5b60d1d577baa4fbdf78dfa3a33d2cd49c250d6296f6060c325f659bdf13c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h518188b8194f32497139c1c52784d64c4ce2d12b4fa3bb0a5c6919235a27e371;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0d28e00faefb40c362ee316cda0627ae7d8b86e97b646dbd0ab35140589c4fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2ca4e409ce330b285e3397ef46e519b242394986763e9f82fbb9474fbb5b1d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb41bea3f0fe2f6140296e7bf9cd2e7de4dbf1a6de18bce97c499b73dcae9ba4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3013f552dd97e0375637bbf9fa1a16d866cf0e14f04cb5dde0f77c23d257435;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb825443a9134aa04a71db0d090da300827084c807de4db913f4240eb6f5fd99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ee3b5bac924586851ac74bd9811c81e635a4f7af4f1ae88115d788453481c93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7909d29376df89d4689e99e49fed9dcf55cfc582c7d531fcb527551406d19e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9947844117bd6c70bc5e5627c63d8d31059aa8a2a92d69f4319f04726420a8e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3330a92338aff0fcc250a344156336c7cda68ae3897b25f42bd567a85d5e1a28;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1514846b1ef17d4203a84c065aec0f28014b8c547acfa92d221c03abd46e4d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdff00072cdebff05b5c1460aaf2dfc87be440739d2899380bb9a75e1f2bfb8e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7cac1fc9f537dc7bc2c705355ea1326c26b4ad43d7ce84a325c99522a3b741a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37f74648748fd375f1ad9f16dd7750868466f9885998d2575e472b3b0cd13011;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hacabb9d7efd3253002e40943f06f630b240653f890f053c776235a16ebeaaf9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94fcc7a7b2031eaffaec433236adab1d43a85ff8b7d2fa3bd241683fa2a2c030;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d956236ed6993116dfd28abddaf7b66d876795fe93f955af725eb764de91f29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9621b9d4ef3d43e3b376864f428f44fa22102034f0b50981ab4d38cea61f20a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eb97e3b0fc8ab5ba972a09afcf58c39a7f1939e2ff8ed0cab4b505e80319c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3806a659466a052e92b0248c25da0d5529a287147bab1f0c8f1551156b8dba0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a1693fdf5433f3ba8b2474f13ab59f1629fe63c7a977dece3012debb483c538;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97244c4c81fc57985761d70a82ed8efe43c30caacfa260afd9c1018a1be08174;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h909f2d1ba363636d09aeba52aabcb78d03f75363163f1a7936ff0be6773fc756;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8946e784d8bf2b5cb66a77364f8ef80876e96c8bb76ba49ec8b42353d3f82f8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4dcecad51e16619f1e8cb34ca4033934b245d12935241c44a6202d1b29c50236;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57447cdeb2e76ee7c160890affe5f2c1a6d53393aeb44545bfaeed0624c60c37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h826f113f866f6ed68ae11096aba85edb6a9ce1dc8409db23fe3fb651c68b56d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1017a098865e31b91e0d16d63e3018695a3e098abd8846e44de7799da42ec7e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h769d6bf1683b0faade27b4572fc1a72e71ceb2258cabaccd78410bdc1b7f27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28c77b300cc2a93aa1ab6d27be1e66a1f7d81ad4c5c891864062160a85134668;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66c54e57212df7aaf1ff88f614bedfb0b792b2eeeec0c8ea8e5406a588ce0183;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha475b04eefa51a60dc829fae357917ad2fc162b122440ee63d9c8edb2e27d94b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cced7b3cb148e2002d5db7a2569016f03fc2f2b9fc164ee50592842c231a140;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f54ed78ff8f5ef86a820df219927adc20b3aa110525b6f7c27a36ac15cb9c21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a36b0d27c1bc948d2975752a8b15ff9f08c5257542ff3b66c7ca3cc87fce468;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a11ea784956da229cc360599a0fddf7673fb99e3e99e31f48dcf2dbe5481187;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9442e6188fddce06ac55aacda1dc30863feb08f986f40c7edab80e8add11d73d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9cc35ef5e79aacf5f677c2c5036139482275019085f6ceafe84dea4a8304923;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he841bbeac1aaf95cab82b8b26db2624173f503f3265e14d6734b997e32389c35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafe6ae3c8dd642472fdaa24b24e780b31c8f4f5203c7777024985b42c0dbc146;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha65ea83bc853365c2ddd3151ad8cf466c389d45e9e2a7eefb188901b6c803751;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b55cf9c7802f3e49ded4457787f7b3fe50b4541b0ff29e46abc10e4f33f9f19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93547a3b459f1c8afcda14af75504d60524148494b4da1f7850cd35690b0166f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f42a1be90848649675cd5a21b99964b2eeb20e10faab7b31aea26b02a1978e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf684311a862667722d8c74b98e5f36c30671ec29dac93bc0b4655cd45d5ffee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1d70c8f18c67d732175477785bf1a8a182463877b6a8924e1b7218479519453;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffb0b3d30e2f8b87abdef82fee5ef24f09d1459884602a0f9bdbaeecc383a97b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fa7ddb1810d73b3dde109412d458d34823d68c8a4050c2d65ffd10c5f6d4e5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64d85fddab9d8b842965da97c8be462454d25121e6999af16f080ca632286272;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b1bdd093447e661c5332d8b74c662a5b6241ba8289b228792dac664415bb0ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16bd6e933a4a4163a7e29b0c8f4c0a32528d46c9ec76a5f6b20a8f93dcf909f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb457a1b23e7bed90efa017b77725c71e3238c32a0e46fc4ebcfb777dafb74ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbad40191d016d74ec7a4a6f8e48fa7bad0c8259e80b7b1539a969d89f5010433;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha124083558fbaeb47ba71dada89f900b5d966116000f318da3df1896eb9edc40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf01926f33c9f31a61fe1916b88cdea8e25a000238dc2aafdfa6a3e512abcadd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1de3dab79f1bb945a158378a379828c25b777ae69747406e196b25e832e77d0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc28e4cc4b887e17f3293c7e1997b0ece7542662802ae3f91cbdf3911dd51acdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h376e433792a3b31b047a888ea65f1369f86242e937032c71b9fffb7ba48ceb43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb462be619c3ad61fcc69309ae48526f92e7c1a7204060f53e1765419117d763c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf38bc07e2d5d63e629d44dfa7a89d3f61f2a485ca32ebc3e8d5101e6126c66c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45834e68c0847ce01a8707bf61b1ed2526d0a74190b11815503a31471bff9293;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf3284bd87721efca4b6091210a6ce2217f69398b0bb6a8b734e002a3c84cdc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19f710655b2a70de2add2c84b2356466c0db34a979153ecff3a6948d808c25cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f4a4cb73236139b9b1f2fc3ae61a0cd9c304d31ff82da7ad89db3c43eeed93b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19a755c1ff20abff96719a0b11713105aaa3b3ebd1e2ab355fa0a4d30aa7288d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f5b6a43bb5c089414aec30f5ace5323da174f3c1243928af9d9654b34d7f062;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heda2dc4dee134b0b7bb00145127d878509c7080b9c46d2319a34b494714bf205;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21935a00e170775134d640e5d8c638d549988e145707d68be3f08c7d0a495a5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32f6dc2939a871c231dd953634d035231833f42515d6ab408d8b8e512b2bdc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2e529658fac1dfdc4983519e810de76ae34da61a4d99a7a37afe706eeb63ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b8d0a5170de326e1ba1fb7bb6c362ed69893dd0aab3959ad618f933bc83d0f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f72c7cce81e930099732515ebd28f2ea3e2a236922ff0653a1f3b9ed9dd121;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf5eb96d86585e93f238b232e386e474707c2e0f8c9aa4612feb17e6afae937c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10bcd53543e12f87c287ac23b8352b9012f250fad15530c2a9ab41d25391bd6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b02a2a610ad7c8e23a7d4a977f317388c130f682792a2a290d33d7b98320fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h947471755e5f5967a3f19837b47a7d868596640bd576be997e12525a807541b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b6d10f26eeb77c221cbeab3518630224e81dfa3ad44b5e222c457dfb4e51983;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd9649fb44a06def9e65208e27c2b0c5f4a48ef2372c3db87816cd696d59ca3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ad7a6845755aa37c14adc082e48461eff5f695aeb532b03f6450e7cb9c5cb20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3288b114a4d968be5aa6adb5bf73f8d8d0b4fdffc534f2f70717923a3a95f1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eda21c9c36dabae8eac8c793fd763cdb23f74ec7ff06355000cf3a660019314;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53fa8b78d3a0ac90e23899a4d5da5402003f68ec5de8f27a2e91ea0d8aea6fbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22df4398f670c08cb785e7e03eb68a4d641a410b06f26915d7fca28082551d7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c5d5a546a2e1612e15ad435ef3e87b6c395e71564b5feae7b95a109c0d64077;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h402394c50a0f524cae6597b749f358591db1a605acd09e7ee2b3b4c0d1fe697d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8b870694bf63c2fe1a2f9cffc0e3550f4d7b64814a934fe6b5d918927cab503;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b2f179afc96a1f1c81782d10d9c4783d7400687dcf6c87ee6c9a7e19311ceca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fe2af95a9c2a7c5bd921e922715e2fb1e0e3f70adf45127f06585630b8a5ce2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'headec2bf1b80b71a8f1bbdc83262306f71bedb7cf52dffd870e65d3fd833556b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98f37272fd314ca15920b75112dbb64d988721f183ca4492fcce6e8669925cbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b7fc6ea5890af710c087f277e39557a42db46e02134b1fed00c3fef8c29221c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h555540a44f771199c745b8beff647f115c4b206a304fe047a952ff6c4101d956;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a43b9d5082908e3079472f5ecc7a4ba3372f497e055d6f026ae531fabf8bc4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a6d70a88c0634ab47d86adf55a90d0253350dcd37e0ff1b341b54aeebd14c60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5c77417a24b57431063878f2085bcc484858316ecbc2f46d50dd903cbc023eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec2dd62bc089321e3c3855b0ae0c688520873740aa47d389366d0a27cb4783df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h155fae4fd29b4ee0c38e4f0b97ab498d3d6287e2dfe7fffa46edd541cb43f520;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2c0623c16965a462b0d9eb96e7a6319a471a62ce0b890ce8131b2ed529e106;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h598bcf02bea481524c4c59927510cd0c4464ba5f645eca2c44ba14c49f42aa1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc529109d1a9d53ac6ea18e7d6f48bccd3109d53f1ad3cb6c3fe9d3bf5bacc0d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cb3a2fec443e6484a900d2aed589c322dc0c0f4a36d25407b26db124836b040;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d6f54c767110982f766bc9a51f2eb80d1884ed717280f5fe8987bbc2a4add67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb622ea444c283742347a0ed6b2d7983868f8eaf601a4f4516344979c1ed2899;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25321a2842c8be9662e893a3589211dfd76900f6744e9d5e393e142e6dcc4d1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d1757f6d0ab3c532f6f3f8e28f6908c16888071506056521296b23c3c77bca4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52751ec60290d734e32c3ff9f1cee21747e139d9d78f9f1bc92335fab845f5f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5ab433fee3604549429e1c147909d889fadbc0dabcc5dd4ebec5b067a4b5256;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda3c64a1884c5748f9acec83032fb25b54de5ff18dc65020d3c1fae2eee5e320;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94d82eebd7e914e9e433869cea7bf59c759ca6d265aa29d76f80e84b8ff4029;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac25072ac2d058621e2c51ee53ea5af229a7992102c869eb09183526d8bd2fc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dfe4f221aa66fcf877ee9330b639b710d7870d58f0bc664cd8aec125b73647b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1262770b6b22a25737177e366ed2871da4325bf73e98d3fe230f342bc36d552f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2db26aca682ccc653a7ea88e5d805f33cdec4bec930a2b4b57a056ef70754da1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb989f7761037305b660d5fa28980a7ff645ec071f500d581810e7930b8b5fd88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf4c6dab0e2a792287e61289cc1913d2052b7e037c047f82a333500273cad17f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd066e8c31835e696625fa1da58dfff447e3783eb7188cce10b89f9c8ce1ce5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f3e59075dc428ee6a1c42a60cca8fbb255b7d0e6b8d9dfb01da58728ec51515;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22d0372e849350b31e5bd4b92fac865fd38d149836c25f25273581edbb9849ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haecc60206649ff6c8d62c4bbd84564fb9f91e6ead6daed3029070c8abe237554;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h952d4b0da692a9977652e2b7b0ce9f42df9d2e2773d124d7827c8bcec409292b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb8a7567e190cb86dc14dec9ae3a83a67f1b255a2e3c0831bd0bc7cd752cc380;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac3d45dac10167c5707517c4272e97fd1a726baec7c87cad443813d05cd8915f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95513e998d48af9f410c704da60016f2ae85e49cea052b37dfd2ae63f809eef6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha524bf8c7a06bb797ede0cf31ca36888fa7d50c7e9cf7c97b7e36cfadbf3162;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73c9f1c4c68fbb9d2109167df89db832d34918f8e0ba02ccce6f24eeadbb8980;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha46828cfd3963e8900ae64d9208ef16abc3ca8816598553bbc8c6b341845fff9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70fe3e7f86e7c307c1aec8494d53ae036c222f998010eed4cee8b7750e804b38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb645947762eec035f7f4b7c4ca90133af7c5e1851b9cc8217ce7f0fc8e93cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h871854df3564a426d3bc51da6961845dca7d27f55f5b173aab300188f8b54f6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha800e6cc8b8af2eeed4205effcff39dc583951bde8810644459197f8086e4485;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb28aab9e9f79204fad9c27a8ab82854687012e9657af8aab2fe2ce9e9f496a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h572b2aa70cfbc61a61bba646149e82201e2ff3f73d3a928ef62010773acca54d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ad19a3fb7ad4da484afe8c98e9b43760ddfaf903a2139821c73e2ea7b8ed241;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e5e80c046f8769719ccae007e191b7a01c6b0ba4dba42960fc6c48cc6e8aafe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0a4596e270041483598374049c5c91cde7d485efa60ab49500c6c965c0eef7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77db4cd04ac1e297953c607cdce3e4a6209d2542720cfed09b7dd41b53e4addf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h806e462af24d9f40b3786499de447ab701d22f7929220e58cea93ada3b3a875c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77eef86b55e13be25aa58072c5a256aa090949c749074cbefa7a449615a50f2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8e7d2f6c01ae14e762f5bafc2f73108d61a9218ba293f6ed116364ea0129fd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64213296b29e6b88b3d0a97813582a0afe472b0ade28cd99ae8d9e03df27168b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bd979f139cd988d74128f5e9f5d7f72ea7d28ee7dddcf6a56d04fba531b298b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac55bef9d555ef729ab37070d3ec99b23b066b281753d7b0f2cb149f371d4cbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'head434b62c7dbe36d004a23b5a04b0bf47c3a0c88029a38dda9de57ded246a89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbed74640fe4dab3b8dfac17eb9a52600a83b36163f5f9fd5894b4dd166151a5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d974c5d8631981e6316a9cd0cb5945f586a88ef7d867aff3af9ec89d6ca1090;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f013038b6cdd0acc952a07271c5adf5b0137eee99d2600c4bc00478e884937c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb7d6ca2ed71cc1a2048cfa2a8435e8d0b195ea9eaa148764c5491102fbcad33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h866c46fad274981b0cf223082d84033f406b1fcab9b01b62d2b5489321afc5a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h972c1d4972b7687273d963d93ec86ecb9cb46db7c9968ea74fed0cae76b216e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3104f611c5e32f1f2f053570ecc86e6690e438f078ba2a2cb1008ce40e6b852;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca3f924dec6f958040d290f098673b1af75cdca5d0f864363e0956324a537bc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8a57ae979be3c36ead55081a11466292cbfd9ed88ad9a78542e3d0f0b6e4c10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc228dd45824da74e6dba29d1ed37134f70946e6c57e09836ec886a70aea60c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6efb97f3e37873ce8f2a3350d76b0a1bd5cf3db1703e0efacf45cacdf251b23;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69e55d978323f4fbefa4672228cd5d2c9d2f491c48be215e9bcb82ccca358d45;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd51499d25230f58692878715e6736ee824bca53b30ae967a43e54b54df77c6e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h752fa1c5ff6e5a69778e41e9d1f03a934b83e51cb224b90060f0caf133e9a7e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4404c91ac75152d9c7c5994e8afdd1bc02ee25a9231f9a8421a5339cad6d33c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e175c079be5b5d5de12f3bcf819eb92eb331069ab4bb6cb12f058eb6bb0fede;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28bede5fb59aa9635900736d97f2e94ddbb821406a0a4d14697b39603ef3e337;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1e6fdff674e0d8a2ad268953cc1f7b3b1b3844a43e8b8754851c95a584ee6c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf03eb6fe37aa4015891aac275a9760af3a2dcc9f0a68cdbf1e22f182e351ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc210f1a89be736676ae6f05920ce66e571b9aa83c5d7f1371b8529875c7b9d88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a59823abd9730d9f761f1c6b2be65a261a90f07294c71b0ba91f8de20781854;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40c0f004c5e94c5dc1f4556caab18b0e19043ff61bd835f68127886f4784dd30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd13e0fadb2cf9bb008d97d7f8e52285b4428abc16f81cdae02187c1df4ed5b36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7083fe672e9a304c484772cac2d771cdd4e5407a8e5f3c7c102d630ab158959;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84be32b59462adef18b5ddddf51f611e22f8eec45026d1c01c4c0792df39cf01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1abf1d4696d551dcfa3c22822ba3a3bf91f3ab989eddc77e34aa521c70f8037f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4892f1620e82169a69b9e2d5b7309b861b739d3778baa14efa37cbb4306d47b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1058fcdba56d19ce32a85164445445fb6382e1c009b3132193e667a10d488a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4e52b4828ba55043d35e94c2c56a5f673bcedf9a8ceaacb5fe5c2ebafb7d291;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70874468456795ec2917ef53991b615aec0ce82f96bd8f4cd89be5b1a0bb38e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfaaa64adddff59eaeaa3157d2f786aeeb41146492504c39742d32aa22aa06ae6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3618a971e4acb425c4bcc921c1a9ac1d75d5d2083bdd5709287d5df1068ded99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39b2578656bacece22a393a584d22af66b0eecad8da51fd4530728e0313a4414;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4809c5dc5a90123d76bc2e2738a5ca326106ec6bf5e28e8863cbd3536cb83ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a8d52b2732af63553c819f070ed9e51c5f90701a24a24a1465711215d84c1da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h670fa5c1cf41a88157b53289fbe19aeb4cb2060a0589ddb2bbdc11082c9756e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f0504c16768f9512a756c20dc700d5e85fce0d0354a7bb9dc0e93446f6ae1fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8099b5ae973f82b578a444a2a22b99a4e27af673de60cb79b0fd05a9d37e55a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdbabc4ee5e033aeff04cfd50465e476531e0be3692d249b2dd00c399fe7c402;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6001f0159072903b27c44d89066cf86acd7945311cd5262d38c32d281acb59f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h309cf220401125639176b90e70052f284a67bcddc27de0c8e78b3abf2305e526;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d871ad19e97493252e37406990ceffd8f2c75c4083d54b2fadd1acd4b055396;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fb6b4d63ffaa4636cf989a51eb8dff0392891680f93566258b41b46ac5ca813;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16c8e9cc191d256b418e59d713ce05e51e31e6d44b4493f2b2617292cc3c3623;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82215a466cc5c3125849a0b850b1b7c1feaecffd4ff07251d6bb818cc58cf983;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6162623df2a8851b4621bbab361ca09e312e3dd8c196faa8697e104387c1363a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92ae3dec9e82c2d8d9dd268dfeeb53af0127a555318ca9405b29e67bee80da94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77104ee4b4c7e1f4cd1d74eb3891fbe7282e496c3afd700ecaaa449015a88cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28559f2ec6a37f225145eb77574923ecd754c419cb1a5f5d25f125bb5de740f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e973eeb15400d86a6559a81eabaa0914645d2a9c9ab5f9424d7fa8294f1227d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11c31f6c45f162742468693475b3dbf3e26a6d17e15e9b6b595ab217ee0ecc64;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce3067416855540194406f042dbab8944773120e78050c4598b20f836d928228;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdd7cf9e238bc8e37d54aa94ceed75bf999124a2548aa58979ab797b79279ee3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc32c3a9c15293d78c9e60f89dd3d68cbaecc34c6daf745cf716ef29737a0dfde;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha55fb1ad5c5ea34657b266d4e36b88ae895219f06453a8d7d358ccf0afc0dcc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2271ba2782c68454e9a1eaa0467ffb4ab88f50a0c8c6ad7f989eb86c89b6ce7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfc5fd3228d769b5a2ae4fc5b018178e0b018e832c92a7d7b78ae1415bc65f1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h369e0d53adf97d57716d5df7865a30de5e3ab215ed6bd3e1c9b209c69dd74661;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cdd2c1613d7a6e94b8feb439b7ed9fd3285610a490c7537418d68ee5bf7f994;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf32bed05d07cfa967bc0c7f630dbff2b8cffc656450d6571f699f835af4b85f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7116062b6dc4228228e3047084a36d21003cc0f2225e7f5151974a1a35dcbe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7484e2303b45395dd658ed3e69bb54493f86768db3e836426142aa84a29a046;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11583c6048d3de7a3807541049622032b8be5ea9b1238f98f0ee9c2567f148aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ed4841b76a2599b2811ec0d753fee91153ead655e664fb6ad8d01c3dd98aa24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha540cff59a9e8bdaff92e3b71659c432104b03380c29e5bac0c54d8af2da3668;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfab62b476ba8151891e3ea4a4ce753a443a93162a8a054e1c54e80a87877004b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h177e09988b381aa8ca1c35c284dbd05b3837905235f820386190fc1aa485db4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbeca76da69eea7d51b5b711576d4eb040eb24673864f954c855c6240d5b01177;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a1626f07661fff94caf4a43c3fcb55cf5c16b3d80afd3c1ca9b9a4a711a9c99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4ba0c6473b8c3b6226099985562073963e4d202a7aa5b5c711e842f4d4304ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fb81cb1f06c9d659ce737b75faa31343e1adb1d18cfec4d5e8a5a2e5ff5839a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f1960d37cadafe0d55cd9d876e9cecce50a7b72cddea21b34f27685a010ae70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ecb29951ac1518070f908ccc73f50fb219991f266229682d5aecc28e10e7d8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5be0c1cce963ada52c12fbe13ee85464be2330762d53cc1e5194f51c524005f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e52efba6d6e9f27bad13879ac48beaa875d43d3e3f5aebcc640151dad4c4a2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62410d8e5da62f78b80c0faa15ea83b087c869e98f8ef1d4b8a49db2c640a428;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5353baa5ace7e6976b9a8b25bee889edd5f9b7ebb309293f46ba61a9c36668a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34dda683b6f34974b9f7b33addb031f2553e235addc8d8b27ffbd28d802d2017;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39b361da72328138ae6f203768dd6cb35986879e0024eef5504708e275fcc70e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2468ea3cbca95e4fffdf8339dab75f682c306a4ff59439d60a21f4175de5038f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2988636f7fedab0d3639698d45ea21250524968ec14ef73d4bb52a290c9151ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf98540e6838e6b34c386c85ecdc603962aa1ce32dbf6578970c97fc996e59bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h563f4ce5a6d1db9301f31c7d8d4ebeaa9796e4e518873b1a8baa028b5a9bbbcd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h859858049a62530ff8849d0537ac662346be311d97ef6dcbbdaaac53832550bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2710254c32f0ac1903f97e189d263596b6b9526d18576c273e8311602a7ed793;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60300589c0ea8a67fd00f293bf72646ae23de01f904703edf92534ff062b4574;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca23379ba36e39f20ae68887d90768dd903cd8285fe2e871535554daa3833e67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40224319b8feade5e88d5233553ceda1adf066ee5ee68f7b86252996222fd798;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ba0a4d55c9f80055a5f98f7c243f66079fca187366e223a69dfc4a7d3f8606d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d67582521f1a543a2374c7fe324d15087a1f55233f9f1cabd2d5b0fb56f75f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h777e74871ff66026d8eb4170520c81b9ae05c36b16a034de6cfe912791e3e572;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e14e8719edefc24dd0343340e19998b663ad251557e3012a04d09a29351feff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h716848cb5d829c13c7e711e135a31a35a3d090d21fc4272ef7182fa268eb43ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf1ffcab55c411056eab74e30b5049711e221c369d06ea7a6162ea8d5873803a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda08f82b1f07b282298fb9da5ac23734c6ff9063de1637ab304db842c7fad100;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58d17ca8e7d72ce98d8148a4ccf2bc4e57fa4060a7d53335df7c75132c9b194e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b0124a129b832b180dec2ed5b2f1093301e9c653760e5e08ecd8721a99fe40d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he617b7a20064f71f2061a25e6835e4a4a2ba0d9e096aadbf80578bb45b659008;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e16c7668bccbaf0785a1d43fb62f643994a4d442a055e86f9e43fc1f71965e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h718558fab09cb36d491c065dc4dd666a672893bae3115458f4c9184657ea7294;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40991b06cbd905745ba2d1c152e69da3ae8938669fc30162afb1a20c3de8947e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5758702f4c1aa5b15d878d141a9bd36a152b0aee730cd2fb5c9031868fe949e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9815bfb1efdd4cdc243906d1f9182468c57caeb12be7b59409aeae372df028e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h802d3e7beb4a8fde8f7cecd6a0b9121754f3431337f8b7aa8b01f946b40472a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha00f32e6c2514729ca60858682bb41fa16c839e931c1bc757e56bba4725feed8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfdffc4388a8e2a713cf4c30e6d354baea3a1c84466a921b3c104e7563392424f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc5c780adf98c218a8cfd4dc7cf81fb9c723d29c1b143b5c64ea8a90adf413c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5194c9a4c5abaeb106ab0982efb350f66098c21b0748d939314a182df717be82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e9f99fbd23e409af67885f9efb021d0193d9b36a40e360fd33ad3fb449c4dca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h247fef3b43699551123d2f4e4abfe017b58fb4eeb3f894e6f5b33920044745e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a37de90d538bac41dab156cbde91995229f6651d83d0c6ab159788568d77ad9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4356bd07d4761441f68285303ae587981572c3d3bfebb145410acfd7211e12f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14828774d5928643054d1fb495ad34ed5d9bfd4ea58473c1732634cc8d68d2db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15692716a895b499194fa0a63311b4c9fa7bd4c2db5b7b5577d350b2e601e8c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d50e4503e265a9da4ec0a130650fd475d5d47ba80ef1fc9499b362db1d9196d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59af16b408bac2b2671901d103c59fc6f6191d16c011c9d225e6e984a246c97d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf16b2aa144e81fd7721990a47417304a9542e4eb76aec3cac58e1d685cc9c05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf8d4aa677844bdf50a1a52afde017e7366577890a403b06c992c824e346348c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7f3dc126d5d3322b94ba61b22a12d4b9161946ecd20bd18f1646dd179cb45f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfca8a66079fac29d1280f29330526785741ee29ce3aea927b3c71746780e93ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdce0f19fbabe8490797cdc8598241f8c4e29e390f8d3f40284b2f4ddc6f0ce70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha668cd3ed4cd48c8d27932adb13425d1bead34fa02dbdd7f04c672a5fcc54fbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2605d161317ff7d14a7ca4e6037c15f6d1d6bd3c958a6d0aabe55776f9a12df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8786386e2c39969b70333710b78afe85cc0f08725f9365e7cf1b108bd336f961;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a78f52fd1193028952a8209c46de3d55588d5547bb09d357f66148228c6e4f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c0fd2bb4a00f9b89ec0883802c9d04623cc05cdce2e05ceaae44f484b33e59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7b8cd1fb71a0006d2f85b860465e691654d133e85509e6d1d08e53c6e5dc70c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8c50db7562b98d9599388c18a1025193740ede3e733be9970a6e20f3d23d396;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfca88bef998374fb69c2fbdcfa477033d69f7bba520980a64742477c804558e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f52ae5f861dcf7271f3990229dbfa37eaf434281676a98e2ae3a4c871fb8685;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2de0c6dc83ba9221468ef1245ea6e1e5fb569994ca6943e24eb9979395aa0e10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b90e48bba36f2ef44cb0047849b6060cc52dcd0877288ae6016210141c61c0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbabe89affa9baaf5c51a2017780427fd1e619effa91571e6ae8e08343049ae21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2f1112dffe132718e2a948ae03cd94279ed27c5238d7a31cdc86c7eeed80203;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67f5a103ceaa68e1a9f47f6de1d11cc98f125c03f9da6c2f670cde2e7d30a04e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf28ca3e1de3e9ea89e63c327117f053313af080ddb39af5295be374a48491c63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0c498652a69c58c813bdccce6a029a4cec951dcb1c4d4cb50b2d05b45bf5e6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844ca2811c141457e9e384252c818f727795d308ae8326f81cc8ac7d3556104;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbad0eaf8ef22125e084b9254ce5ce6eda9250c25985464854b93da8e5a7e1bb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaa543f1dfddf242229a74b72c4f1550a6bc8bbb9521143d00fde76927708d45;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2aff829da99c30838770ba122a283febba59037a5aba834814f16184eb9ce39e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a6fb9e8fd04e915f1b338e6f0edcf63b1e910837c38be3f0e745bcb8f47b3ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84b12094af4012398fbae2466ecf181c59dea6c69049ed54f7088966ac70884b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h803e1f8c433ea67c2e4db8d68d80f5c0b187188dcc1a83c503d1a32d9bafaeb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9f41fcdf4e5eb1ec64d91f655257afaf2b758754f2d287725a610c651d212a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8de2440c4e694ff0e5d1951731662401910a649b3fb7bf04c92db558c8a81d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha134ae156177b63979360fd40e0befd042846e00301c0d9850a83784568c10b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2a646a5144f38755b47326a8dd9bfba20be2f488872c1a45688bb35bb5c0d65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1443542b16c007e3c375e89ffede1cf8e662d94a9e6edd093c174f6b268e7f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23669b895e88702a87b1f5ba178cdd28c946b3e48c626fb6cb363c0b8fd2127c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h951c92a9bfd17ee42fdb0b573f20542bfc22774b2cf7052b1b0e375d7c76428b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20a2ec389cd828fa3198177a43e18d8f49194d79f3d35e4a2c1359f9b28fe029;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ae8521b5c58bf730dacf994286087ed6af4901541f5d46186f40b78fcf540ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42c39d1e12374b9b729d83be8e17ef44670a8f7e20b5dc38f98fd2ac46d78f2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hece626f099809af27a11f079a349da09728d73f33f88ab944f4531ce059ffaf9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5b3a12b9db6834e6f28a1c1fcb93e311f5f8d3eb4e768716578c98b8b85bc9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82e1a376f455378b10e14917a83d84ca90a9e565f0c11370f028aacce54043a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88d8980294f5b5560cf4dab392480b412ef1d3a7cc007ada7c4119272cfe6248;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb839684a2a63e58cf2b2b319ae4856d2ebae3b19dca6eb3e75e2e6696b200f9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc09bfcb79d40de07cd7c7122ec257566d4f73d251a55a319c26a8c13b571ecdd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33611fbf0093fe28820547d95a9942b8d066d77c696e2f9abf15bd3465eb2798;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1557fcc9fea7624ce6823535fa5ec4e188949be6ff06d23a9d287530ce18647;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha05eb910eab2b43973b59605f76cfb71621abdbc26d45dcf4d32c9b1f4f59a2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2a99e190e2df713e7ee19a2c678a1f18f251139bf5f6d225de50944f184ae5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4419e789c394d9ba25ecdf3fc8d1ac936d9e0078136ce32c306e33d23b6d3e73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3e8af0d793a13dc28e90921ab4c202a5693058b2653e839b863f76ec9033420;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf638629efe419dd7cbdb6e0d9f2337210b34478df2da2ccdb47b3decae29315a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha08fdb7b18e125147bd5791dd783d5f48b90d1c86d531c1241712cf7e1ccfa5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9449f814a63fc8868b2e2360271bab7e9c96510cb997ab5f28c2ef633db98ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f875653605bede06588346782d93bce0224e34c18c75348cc3ace6c46aba914;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8e31fd25679a3ab18b376be98a8db888b731d3ecfea26f9927fbdb8c14751d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33132256666298d0580c1c419fd4fc44a605edc660decbe205e2d63188faac4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81fb7ad84b5d79ebe3cd4b5d26fbcffb556c3bda822a486d0d1d9219db8da3a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e0e506bf3b2539947de43c5f861262fec79b98bcb1061e65c6118d3f4ab84a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44a1341ce7f4be0ab1a8360c1a44602614df0bea3eaedae78320af307443adc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf29003ce4142394e6e163a25ba7f2f52e3329959b3850cb5f8ca2784a682bff5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3374eb4cf4817d2728fc386731ab83d2dc0d946ac958f39c26865ecee2a8ff4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedc4cf68a374ae2d3dd13c0b001758dfac006b17ea08d0bfcaebf3427b3bd266;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h225b2c570efd61f0db383ae03b8e21a3229f47db951d993aaa18e6518b8825c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a5130491bddf09fcf3b844569a82ca58ba87a63714a36c04f42e902b681e9ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca924ac13821015f58882b2b4dd23dfcdc897eb2c3b112a482d0f21a72ad192f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfda6d9852ca057d58c8985618dc564e879c1ec05a6d9164b67e1b7eaa907bb12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1de6b6cd3a14f2101d6d0d3e06a694448076d4ef8b12e5cc8c925fd1caee456;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h966700815f2306a7a026da187b6277b91bd6ac28e097b3016282b42e8a404568;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ea637332472da0717841f9a6e40baf8dfa63e6a8377fde48d831fa406b163c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b38eaf92f48089e6933e341e2ec2db343b6eac497dc71036852b72cd93b8078;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f15093700641bf4a1dd4ac457fbe49fc48e90d798418add7016a557b8de8ab8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7ca940966d0a8efd6fae6fc7264efad76632c079799ee4594002546748d4704;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ee81c8912dc917a709657020f8a67ad4798757bb315af57aaa12793e882404b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h672f2590d23fb0aee9258bdb0b9a1c970f174f44fd1487fbdd82f9ad60f9d5b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac2ec089c597b1aa2d054ccf7e953c316a96034a0010759da9ae6a5512ce0909;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8086dfcdaeabc6b0342856349bd4bc1ce5ba61074ad3d02dfd49be347bac55c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9519749717eb9feff7102db8ba5ca584e8506a43680f440c1ca14e3df7db8d84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6ab6ec1a4e761999da6d4bc77b096ea203b26761563d3f62834323e129ebf3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3914e5b2c1488028ec606b5b822c40594d319593cdcbbcdaad64fe15003a1d6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha13cacba343e0fa89d90ebf1994c5b97c594067871fb4e30f97b12f568d00439;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6dc88a70f6b64218eb64261c703178bb41e5e679137f670b135d8b6deea1e72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h481b0e46386c022f13b98a5981f318575f9c0be4b73200ca37f9fdad35f3c761;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a9d03f16a9e4bbb2627c5fb288276b9c9fb60b50eb143d543fc42b7058fb746;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaa7398f42458485c0964c001fab76aade67e31e687b3bc3f89cfb921248f334;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dc2027ec90292bafeaf42dcd88da403b113dacbe06f95ab140bc268352b81e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b3fe71dc27c3992252cc46ef013536274b8213fe9932b80a5b1bc7a510934a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f8b17a41587041ad0ecff0014fa2a189da42dc1e3accad4898ba0eb8eebe3c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h532f1ac59d8b12a7344226c7933d3b17ecfd0b1bf543142199457dfcdd666324;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b9163bfb0415426baafbd87c1c0f9bab6859a53582999011d5e233c5032c4b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc97ef0ee38061910cc444665276b268b04af828f33d161db9a536c56ba3d362;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd99dfb908df7a7e96a35c79f6b257893a34598530490fe6455515703c900f6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaf01e101fbcffc808b226be9137b2dd58fa53432927888bda243fe48c0f5f8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40b23b52569a4c26bc225d13621ff06a5cb6e28ba4b487b1644bf2228fc9b1a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he36af484d2466dd816490c26689bf6cc7293d652be008b4c01871f916a7b1a61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e562426e599ed45ef44420e4de02d111e0e6149bcf3057cc4fd54d182d02982;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c9ad373ce0a11263f0a69288ff074eb523854673b898c099cbb14222e2f59c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf921be9e16fdc2ff721bf81659a0141590dd8f7bc905755e32b53820a0cfa4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadaa27390996a27d9dbc340df94ce5211f2ae4e11ce01eaed7216918d55f5165;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc0770d6ceb437fc18327480f155d5cb82a3a5592f6152d03cf4d4e454d84f51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf23f209e3f0602de32a4613d5d8c12af508823c03310f6108a92a60c6ff9a698;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae11fc7997c0b421630f1d24608fa4df5d3b550de860afc9d7a1c10986b8b1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf90a323bb5da9ad7f7ae8cbb12c2d8bd6ab70d5a18c68a995bf5508c81ba2a78;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89d0a6ccbdddff9e1c16198f578457b1084092d23d9cacc0c4b65fc4751bc041;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b92b277759b124f929621f68550fa4df3be4245bc031c7274dedca004f8ef03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he34459b565ce7569d9de0432b22b4f6027f5cb6d424a96a349b2bc7e79dcbf9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h851bdd9486261723f1a3d1b23bcf36db2169c77c253f010789da119e8db7df71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70bf10facf68e123d0464824b4da57ba995f63cacbf73089ba937185c7fa0a95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7be8098ba98f83da3a6757a878c78a5e1f152e845d874c806543d902dad9ed35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha944363ed2ca924b1e5826ec5c1c4fe21fb51b590d19670252b66ae9fea26f84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he705d902bc85022312667bf06397eee7609f0f43922afeccf5167151f210fb77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7070becfdb869b9f74026b9b9af4fe760ee1a630a8c9f897d946abd6bb599cff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3079e012dd5b5ef73d93ca3be3864c454c1c64c48f8d1a39f8fad7e58e448e50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8210a57d2ebe876f0b963043913aaf79a110c53419b504a3ad4a85c1ad86bef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haef8f9683e8343d7098d147d2c30e5bd5b8cbdfcccc43ab09542487a7e624af9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h144d985e1ce2cb8066c6e65485d923071a90a5c5652f1a713a26316ecfd3990c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53481b88aeee24a7fc53a581b467d711e8aa5f2ecfca6c3427e7c4d1b809b794;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea5b0fb860bc53c41e25fceb8daf43ed065fdabd81f39c3c40c38069d370761e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h487b92fde3f2174fdf2c37d46dd05c428814ff1ead884c19a0707654a73cd5cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bbe0fc250e2472cb7fc5b116c0050b6401a43664a28eb58d3d4fc87da46bd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7db0dc32373965a802d17be2fc2ffd341c739168eb00e5a47c38652f283b178;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c9558cf7f8cfc7916b6614c7b84048c631e36f7d7a52f7868ead59d96423351;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf8e28f37aff81c2b899a35199651dbc11d25c713a9324c16c7aa6697169908c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91272a5269c38ffa16fbe375500be82c5c6a2b9bc53437c4166ce9516f11a285;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4057b3a9c2c655d56236d4e6bf8a74a64616b45d99dbbbe38e591bab32a3e7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5a84e6785843ec21e701e89dfe7fd45d9296812dd11d97d62d50555fb9c0d95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbef86a6a825868887b2703eed04b75f9bd04fd76bafdfcedb323a11b20601dfb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a9aafa17753f699eceb63571aed0a4df35e1da0e8bea8093b834ea415717dc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1aa8d3a04b1ce0ca2d235512c4d4cc6f8990973376f1b0e490de82e2256afa4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2416e88c703a69d1df058bfca316d459a3395f22c4aa1ce1da84606c96bc44a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c021687f1a4d38da4763fa79d3e6a76b458af94e2187bc3324f815b3269f1f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h186f5c716c88a5809e76930f06641c7ef98c1354a60bf3e6178831eeaf566e1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7d02be0e194d34a0b51ace6550cd95a56481cf6590eaea57f1851c9d9669eca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd4bd3052bfc8b53c5169539d879f3a321e72b59a9593d6e5f592f876e18f509;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h801655b81d249060f80792debfde66554b432e1216614f63d28da34ff19fc6d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc853b8eaf4b3e114f09b51aa2572814e0e38c101a43b0adac795922ed175e194;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee14fa9c0447ed9c6ab39881fc2b0e0ebed4949abbb97766dddbccb73a2a9eb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18a38ad7663603fd8b6976404e63939c36a931c5de7b176c85c4501bba3bb9cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9ff8d1d0215ccc88682d44dd45d56e1972f0385ba72a281a9b36aaf6ceaf568;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87a77d8aa684496eb5fbdc300e204cd1abe583dc39c1a5697ff3d3cd2f1a9fc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haccb2a4ba1f03b3474b7fe0d506934d9a5c3dffc8b42e8e09e60865fa6cea43d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a55d13cce7680b25e0ca1d6b933c5aae3ec43e6465825d3837a461f346da30e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb920270b056eb9f7788225047041b59125b5a5352b341b1ed1c6d2a6b72ea0d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec4e53d0b2a4134dafd2bed520f427aa831c24117bd9762c3d7950f1f455bd1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79f77f6bdb0864056309a71c5380bdeb2f2ba5816aa4673b90eaf5f7011e074d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24a12f3945c1201536c7802c96275f1c760e4e97f83f16b898a786bed2006c8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfcd7b6f1bcb8dd0732ef56812a8af82fae4935c1149ff9fa0ea34b223b981ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h472d354dd8adba8fd72ced2f6495b7d856b7a1408b458cb8f73fab4935bd27a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h956cff337418b6089b16f203adfe7306cd02bf4b12c190aa0a1e7969fca27a6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5825c398c437d46e3bfffc2c0b979a5f0e9e6b4f197dea836de53f0ae1b36415;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f9ae1bbf22b1756ea94ff52fe14ae7c4eaef4c04161675dfdeacc6118400841;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24d16d84a6fc23b7b0f3b13d0df447f4b17d8d414122263cdbc1978faadd9e44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d1f61f5307e3fdbeadb7534c733249543f2cb26a15758b0605e3e6e058532c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98c37d9cb6040ca0d6ccded3965af121d5905c02519362453043c48f88ed649;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h620098258c379b1335c979d756ea8a9fd34f75d6896c816682d667fbb35783d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e6458936eef81253783ca159fcdac09818d308d059c67120b1af06b7a18c740;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15e50c676ff49025b2470c7c16c025b6655940935ca990a4d5656d5e414d67d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f4e41eadf36666191ea900bca11e3ea3171418bbab76ccc0978c140e078ced2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bde5bf046e959d4e58a01e1a412c0884d070ac64242cbcef7b9fd03e5aa1c69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51272b38ca50dd30f90ed0d3cd6d42dc3f8c27b6e47aefe94f15a2325e69a2c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd30163dbf22c39f8ed8619a89d7649989ab5b9fa4a3c2544dbf23fd206f28aeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c1001cffaf3ed7935e6400fc11f34faa401e4ce5a0d772cf3e27418dab126fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96113db452bf2215a73cc9b60bda397093f3c6f3a91226351f1b54c775998fce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h323626603ab10e9e3a3b929ac3adb7443f383e37bab70007d758e3635b6e6ac1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ceb72bf25f3de28f6352eed2fac6cd478b59ea20c9b39fc006443809fb1919d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h586dd71f2a2e7a6bbf887be3b69b648c8202da27b10b40f1079876bac85f79e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb00f9bd93c2410eb31f6251a8deeddc49a5f612cb23c0c1966a44de24affebe3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e3a3967ccdbd1ead78f328b808e1429582e3afc4e3bf512990753966b018fc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf72637a5b9bbe67881d61a2bbf45ad97001b5c4e269200cbaeffda6f38999691;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ceef2ccaf3190cc10cfcc610bf68eee8975fd9d691e06059d744ea09cba415d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5adbda03e7bfeb39061382f1aa37208093f8dc37dd0657ce15d2ca22d2c9a19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cc6b607298eb060401419bce42228e7058d843e2177d7399e2714032a3d864c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0d9025331887cf651c3765f950447a2de7990cc2b650a897cbf226d8bba1eab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2be833ac4c3222027fc957207c45f845d89f06f53254d62314d7462b916006c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85c1d6a11d3132e56c34578ec5165bfca92ce161aaba988d3349ce23837e1250;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcca38427604bf606e0349b2ac9febc6caefba37d19aa9b511a4e270bdf13ef66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72075ceef94d361cc94a0a34ab5ce1b1cfc5dce70a1290e42dcfa791a9992353;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62af84bc32c464db42a59a3d715b74a25bd35ae422b5d1077c0ff5a76e7b87bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h888e602c6d751df137a917977c7c3aec08b31c21181eff9238ff70b69bc7f0e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb625ae81085cc8ed4f30b392eb08401de9d782d128b0b0752fe3d90383a6c5eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e78716a0ebc52a09bf1bc7de8f9fffe494715cad82358b75b2713c119be91f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78e324ddce353b4ad327dbcef273c916fa0930f828009b764347d151ca80ca2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64f216a3bae8c3734c148fbf44e69b3c1419af76327b0c0372549ca5c31418e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb564abe470f94efb5212444edabf28372ddb94cfd4b3de3541fcf7e47a95ae98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h542c4b80b5846c7d0e8404af1537c31551f2f9f1f99cdd7c8b5f6a1f58c658b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf266c274ffe7bcd8bedfe9779299f2e08f6b793dcff731a526872bf23cdb9c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50c014df9310db3b57ca471612c8d2d1197e44eb88ef47d433fe45b783341ad7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c3e7322d66ad24dc86f940fda14aae9b80a953a1e2a30b74a95ad73601ecb08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c6c11fff52f2ba08dffff65c7ec5091e1ff9a9293e1dc9975a207b96e16dbf7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84b27d7dc44a9c17b63f5dcb162b281e51a7a853ae43e9b48406818271d82132;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc10571d9427fbd7e134e824152e693c9259e85f2ccd772cc9a756485e00e47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb0fdc8eaed50079244105f070cb5e9b1bb7cd53d76272ca51e078cd40c56197;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d2fbabf4b270a4fd5b3355efcb37ae2fc92508cfe6776a00bd0f113a61f8c87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a7a76fe14243e4ad9ace5fce7b4fbae7783f02e4614b8dc53909fd39e62f4d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc77ddb018de887861c327fec761b98eba073aef841fc83cbca3ba2ae62d03e02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haac871d25ecbd1b13e5f6f6a7e1cfdfa595e91c07119f830093fedd380845aea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57e891d0b6daa83cfcca8560cfb7754886bb9b107e5e813df3fc54e303f40967;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h567ad02e22c08d1b6815bda7036d4256be228f464ed36f7dc98b117e82bc39b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2807a089bc8a095112fb0095a713eca1b2b6740f57ecc9a06a672119543bc679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1a0f8bb0ea2a4581d41c93b0acc5fc003ee6ab5742b31dd56e6bf8202ba0a90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3bcbc25a6b0623402258d43990f7da3dd1d9e83d6c65d5b91350381fdb49c0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a9cf933ead4df94c93fae2c5d6bc81192acabd49a9d5db34be529a6f0d8028a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35029f6f557a83921b2a441ea1fb48154b05e4072a4909814b522a8b54937179;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd49524a7605139310dcf6356c8cef29777021221822eafc707d4ff90baf40478;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb66049c93350f8e95fd07e92cd944f082ec3c4425a080db24fc913002097572;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb726a2de13fd6af166b9a7cc2f3279abf3ece159beff5e616f5f02ea8346aa22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha76436df4160f6b29e686db52da2c0a9b4c9b5fed345f95ba3875daa0388ef5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he68cd5dccacb600cafe29b167aee1be27a34c284d98631876e2bbf3a59de758f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38c7337efb7f46546694bf5a5192eebc3881bef4def3230baf26cc025a796f9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8165c6a40ef10de63cbeee9e7c2e747786a9068661d7fd182b5a617830448a42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fb150543a16f1a7485c565edc40c9f84c1bb3353f59ff38b3d8a9d5e14b9be7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7222b3e9eb134ae81adc6a92f3ced5ef6313aca264d55faaca53557da2594ef8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8da1d36409a2598dcc809c464c52502dc5a509fa278fecfa3d87bcdf63575d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed65d9c56aa67578e7b2dcc80ef95d3c42e46560dfa31cfdb6eae3239e5373a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11191fdd1ed23194ca098b26b5870c47d92307ec50cd6f5c44af88cb121e8009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e3cc5eb494c3a3442cea84a64a0a238eb7f40ad89013bf8c6c3d7eeb6c88910;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85f5d36e991b67681177e8cf94a9546435ab7544ffeedf0f61750cc6ea09f385;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h822cf9b6a88ee80492b5b54d99409febf360772e3bbbfd373a84dd50b0ee7906;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0b8310c447b832bceb6e2ff95caed051ba7970ee3d81daf4e38675008ba02c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf17d284f331cce2418ff087d4e9822eb07eefb9876c6667bbc76591e791cf2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11fee2443c99a216eb0262ce8fe26179e23a65bb8642a3845bbbcf168c2c7a8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92f8056b366fc0228cd0fb1eb9bf044bb1e91e1ef87896e0d2ad3f7aff392e30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7dcd09721d922217968c6a7119b9cd172a5de761f0dd40cfde4881360d4412e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69606d063b76e9a00d1a00af4bc464f76e69ab3ae38129ef157ebdf3a2117b9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9db80c8579ed5fc4a535bd3b13aa648abd1bcfdcdb0ec9298424fcd27c9a8ac6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha50bc765cb8a7d5220515197aab40470fe7b38323410c364fa457494eb65fafe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4c1dd8c9ee9c88833f0e74e80f77b37457583ce5ef6e35309bbc670919dabb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab768705a1f54df43931761ae9220530b9fcef4346cb360630f086bd45bfc4bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57e248489cb78a5b2a2a6dc247dc1a8aea20a053c817efdc256fbe61f7dfa53c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18f1f0e0e9071520c519d154e2e4b94b7d7569c9bda61a35da935d1d6eb7421c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a075004120492743d4f392f5fb30576b8fb6ad32f2130ef5df2e5ccc95708fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20b1545267c935cc7c92b86343a9b6243c0e16eb31396b12b64134f1072ca24f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ea391e57938b7405b0d6df4b31a16de86582be10f82158881c431d763d77e49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f68b910c41dd6577b3fdaf2ca6b9b9208367342019f4851a8cc0f738ae10d08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60871400df53aef8dc7f6e3d79b0d484bfcbe050e669a6543d53baf5c0a9bc21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20a7fcca6570c7fbb88162205ff0b062ca9888294941b8f94813a023f42f8d9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb05f3b66da974c99e01109d8e01b6a8b87d150082e85e625226e603de554a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h412d2ec649acc17719bc8c76a59c57c4da85192cf7e6543e792d2abe705cc9ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h289a884534dd878855995923da40b6db964714fe2823a6151e26534557e4e99d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eac7fce4516043891be95e3e814c6b52821f34e2ce06a5ab1aa022ccd389ff5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f9dce1fefe6d45b0ec4227aa6321c02010a3a06430b4ec4041c055afa2623f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha913d54bdcb488f12e3a15546344752d482669df0669132a326a9fb935966b35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h855ee8c842be5c718a3a314dabb145f35acf93fbebd8197ae8536d63081ffcad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4a05aa30ceeb3a655f73e50cbe8cdd6085505546ab5009471668a7454b0917f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eb70d5a7eaad4aad93207c5e96ba38bdd53eab9d0ae092c170bee19ed874c6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9b8c5f7e3293d98eeb387a61837a37cc6682174d2ba23b5ba323705c128c2b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f3ca4b06ae4dc0fefa32df6fdcded6a818e33e032ec317a4d131a9e1e26a1b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77be40331eafb497d43bffdfb38fb99a2dbd7172ed7bf729daded1a4bf7621a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49f1fa70b68ae5276c2d77de0db05a2982c338da1eba00cc5722b8a852e76f8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h203b2bf7c50efdb3c728ca1003cd6c90a171e192ed5c1f1f24e49bfade7f7536;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42a1a1d8847a43b47880e6cbd68a6e38f6db514ed89b7c6d2e9eeb943ea60bb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e64c285948d451d5308dd1509d990c82c03e9d5f9f9935d1d45db421e6c2679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf53a00353dd59bece148fd920bfc16c56e239938b85f4f77aa04579ca4dfb89c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf05b4b8aaf76ed10b1be43364f5fcedf597da3204613add0d10b9e5c9d4e8180;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11423eecf0c73f4ec1e08f991516ecc0c4801755f08fa849cce44ed42e928dac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd608a469f65340aa5a46f3f82450f87d10ec1b9589bc170692db662053263cb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35bde1f9e84fa5164d1306aa97ea590992506ccbe769e63da8eb613ff64299a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6326877cedf8e313100b292103c0d7700273900943e2735621f3456837e035c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33274d69032deb95bebb26d558ffa01e4173dbd11ffb44d75e4379ce6931647e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6394ee4273c59cf2c504af0f03e480d474fbe094534a6b72059112e4913d174;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heabb3453a0ecf83032a62260d22f5634b66199b6f0103f90d22db9498eb89827;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h357b58eb01f156eaeb9a282cfab7e10f51885d9741726f1f1e8abed3cc16275c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd553d7c365e3f718e619b44f8cb25143f2731993b15cbfb65f35fd85ab784ad6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha25a78ecaa3288d6037f8164c39cffe8392d3b92c1d3d70a1e30305069573c65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b509d75d354725a1ea61bd2ef8f53169d8c61b6df9d5c0f9d1ccd27791dedaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf79d954a8377343a9e2a803bd39fe4fcd491f2bfcdf111c8a5fb12d1ea413313;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1caf08ea9e984b9253660cd5b11a80a37233dd06fcb6debc4fae233f6e899259;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d7feb9b62038d9510ae4fb138d34657d543755edfb52a8103005164b631fa0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1eea4e9b29d944330ace479ca8ef2a115f8ef98933b62e81a3c6622015bf251d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c5743d5a487f97267804162d14453b7a1237c1d025914e28d4f0302f8dd23c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53e38f77518be66813c419e607a6578ff46bbefd8d4153bd03a0bce6a5b9a094;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h656c30e86ed05019eb5e5aef1587e5f3c0845891ad606902d4638be26a062e29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb32dab9f40553c902e26b47f1b1b0d0cb76b82b95b8c18bf3be5223cd1fedc75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h254b34d7188dedb861ec58d9e8e66141b1a0192866c2f88bfbf9ba8d8ecbf294;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha71b7734f63fe6e0a733b39af45c37a9cc63504808e1e16c97ccaefaae406020;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc39c617ff56ab86ab95ce0d1cbfc1a286006a45f769549138862f72a886209d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h913d026d20245faedf9280f4bc1cc80684846380def42687b8fc6d56e6671039;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h205b19c90520209661c40ca67f1da843615d5854a364919197e9545b3c23285b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a9ff250a5b704ba13d332e20ed381e97383ac06a9351a00ea9821113a337f6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d45572606c1d764d5b73d0818b5be1968cd6ac6ff66cf77fc5382bcf067bb24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h773301c24370c2b976deb430696b48f0392a92e05a72e13b1ca722f4c7155f46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23bf01d22910fa547f6f0fccf2fdb58681a852cb341ab85639903f4d2d92634a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha782087a63a2d08be237032add1c4c9c7b6f831a0305977b8130ebfe2f5e3214;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4845d721d8231f71126fb03b0b9fb105bf2078c8155f47344668f920a88047e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44038a1c1b577b59c4285653c0e440e73cd9a5719e689b4b6abdcd5bd8fd4bce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf619721dfa6bee722aaa0659978f3a50378a5dd37caa75663ef9e4f9cf177aac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf23d9c388cf9cd3adaf2a0d1a1f1411203e76e9cfafc7b10b7570b1bc06eda7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba2f90bcffb856e545baea704f2cfe2d534f889356f3b13b29629e5a3e992d82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a40a8ed0727bd7092e82635c0cdf6645b51d95527775c202bc93ac96f5fbf49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5c05f0805d33c41dec7dd61ebf4a7de2dab273e2b4044b9ff9ddf44eed55917;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf37847eceaadbd0894039790fd7c8f91a5fb296310252bb21c521e517ff2bc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5006c8dd2bb4239e509a29df95abf744887cb1671c7b0ef220f269b8393468f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h104d0bc6843279f3f007b7c78dc90169ef1ae1d82286cc985d43b069d0d1d33b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf95d9d245e6b45c4e8b8159a422b5090852f805dd5de8702b9b1246321c49d11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d9994c04eecc24afc8d5dbb1bc2c341514a2f260ef75b0ac4593da7c33c1a19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h220c27ca89901b79b7f5e4b930042dfdc0c429a65d16d3ee43c70519db09ed06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83d03d6d471f48a5c29f69c08fe202710c59d92f8883653af1c439bf9a8eaa4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74f91c25c751ed2a60d111071f4d8ba2b70850c34b3f058ca42ce013b513df15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86ab74abb64808a00b6424cc52f38cc45edb3c6d1f2ae33b39d28713c0afb6ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd8235cae8a42940cef635f5cef9900600d1401ec9c149bd1bd9163bad80fec1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5091681add43a94a454c04e280bd3173397023d180caed4e78c61c95cfbe762;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19214f8f4571664a1e06c0a81f62d5270948085e87d1002c0b03692e2d27a230;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf928245cdeef444ffd3d07ae3fa5ecc64f09d1fd69fcbfd50b6469ff54486842;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc839203e6272ae4a87938cd9307b1948841eb9a04119b6ac99ffd645861a97a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4df22b2c941cd17c9ee4fc5c183cc980831da994e4e1f355dbad4a736d2bbc88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6722beb0bc6850bde31f7cad0f58a0301c93bb31ef3b7b35d9bf870d61fd38e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a6dfc8ab037fb5d1f2061bf08fe0e256cae5fe0fedc8e2e3a4e97db03cac428;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h293afcd4d6e258529e2e5f141f88f7a99f6fe1b268417130bbb0ab810bd623a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce6296b355ddecc8b634d4f61c0c2d8710e1a7627f7d8998165d9bd4a3f8caac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0e9990c02b73f1464fb6eea4bd8e9d0487dd487ce8ffbd53875708005ed7550;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10b7d111fecce98b795e4ab94ed410a41cfddb970b8322c2058a1fef93e29c24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84dc023a29b9bd0f1893155c60d1afe72836c1df7866d789fdfb3d4ed6b78c4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6d054b6bf81e47bd9b109dd32133b47cc4bd8a460cd6591037f72b16a08bbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8a37d3a8c0101ae7f53b60d2a997eb72e686ac5b50e3248556904b8345e3eb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5bda184c3be167e1ac73807ebcd6704f1b7c2d110ce4d7bd015da246eff54a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea5babad8d51aff4c79b6b3399b22e1873fa4f927cabb43186ce8efabbb38a90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb16a0624ed2b42644c352d77a0c54a8e0edac4c633a8c881cfec6e36dc2a8a6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68d9e3ff45d4db5d33ca728c7effd62b27652b2432026f5c1522ace6e292e7c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80774c598a291b78975fc8c9469731c8010f481695a79532c085182832a08dad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfea4593e24dec2eb9cd1de1403939b5e378912e7e1ad3177a248621e54ea99ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f95c6a033a033034f864ef5b1847b34a56d01e30770851d2f667efcc0158dae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cdd7f8fc69ebfbb6111157bdaa97409226424aba71a241bb4cf7c6cee081625;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4280288aa8d4a8f766d909ca38b938e6591f8bc4cbb2db307f5685875bc20aa3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50dfac134e66feeffda328e15cd62e2cbefd00085de4bfa655112b2e9e3cc669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb93f861a916a18ff0afdfb89f93ef6e95be5be2c5647f99ac150759c9a39ac4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he39592804c6576773aee017bb27ed323308a55d93a3465129275131dff21b943;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66a180e338c635544a886a40a2915afec682906a4a5d83e37e2568954813bcf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40ed37f5854dd28b8e179e367822feb3b3edfd19d3404e8201a8b7eedea58394;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41a62bb058f2af53e9043eb7eabde63ca334d9a3e9cc155717a979846988db9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56d0ad298c09d916a2614da1cb49559a399cadccea8f8be64dbaa6fa8b720659;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b8f06985b29a0a3ec8d266130dd80af27e7b24ee38d8cb17b0c98990ec104ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he86fd05c8d121b677d1862bb6f19563c334505c642062d89d7edcb0b1d9da0ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e6d9ca37d4e7a04ec8593030e18ca2427a26e7aed9f1b844ef2768e8c43ea9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3390721af4b9c41ffa20557e3332ddbf6cf653a63e1849ba804199dbca609331;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17164d736f49ba579232112efe776e5386a57f68371a1fce2976706d578ae45b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd89b1a7901bf3f523bd441501c518bce1960056c0f582a19e64a7c28a549083c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf8f81556e9e2d32557e4fc1c40b1ebed52a08f0b949f30bc8fd44dfb61ad440;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65feda43fefe47876cd92a264516be8d04b957e6c1fecd19f642c75cef5db921;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb676c7251b5bd02ba8367562f66f613bece5693ed746da15ff9c1fd946b90dfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc371ae1e8aa0627bf724d635e26368d561c9ef607f51b1be2af140da2815a773;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f7dc162882f41a048ff77423844fa79b6bedc1bff8fbb84f24a535654df7bea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f86df210edfb2dd90ebf973d06c8a099110022619a7569ec68798b51753e310;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eb110854699d1c8474d6d0579c2517747d620edc60637dea4cb61582e5b55cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb48ca2c1e6ed163dd329d92d3af55382de2d573efc76dd530fa092367af3929;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf69837aa488c0084577d789cc02bb14962f05e1bae9ea1f3c0f4c530c3f84843;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb88fdddb346155d172c4f19104d0a0227466dc3fc782b0dcc9174f240c46d05c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d392988e398784f3593abaf99f3befee8008d17bd3dc11f7bc7b4e72a1549cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2866e406bb2c3891316951566c9402c4a5fd0693da1a3e6e154d1b50d842be12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4c7b32f16c4764382a6ac7bd7263a2f8bf759845770b6403a2d26a793f5525;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e8991bd5a5bc5615cb9d08cf546f993db12784c68ab6c570ad16741fff13dee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1aef5384793bc5a082d6bab2ca7e1b9c14c31c844fcafdd81b105e084259cca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56b5cbb4bddbbd8f458abeb51baf158e120e0e4dd2b0f66d9f51aa09e505e928;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3628d572d9631f32ee99adc6fcbecd0e9ac6f699119be94057e117e08c4011b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7b3094d0e3932a4e1045211055806e7878e302064fba8c4327996daaa43e2fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdca478cdb50b4db5f21181cef89d283d8c77693eb5e230d98ccd2880d2cc5be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fa386957504a31b99c8ddd26544b217035a08f08b112f606e72b98aeb594777;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h615fa2591fb0558ca6916cc9913e9cc70678131e810a4153c802347d9a9efc17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h867e842207139684bb9e5f3cddbde3b0155470c39bd8dd82fc8cbc16a3ec35e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1b273d0544a5db45582f0dd40330321de25ae337cce2c04bc00858d2a8c7eb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac1ddfec3da608b8105c63781c7e9b2449158e4e2d5459f6aec7ddb944a61ebe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5650a617c65e8790a957d1cb8d5e548c48bac47cda5530006eaf5dbd1817806;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82c6b074cce9d2ab0908eab9f659d11935f7c0aac399ef2069eb107aaf9545a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f0745b415ad2ee70905b66e554cfbc57a7651c346778d8f4b440d0ecf956cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7402803f934ad6e3aabbf82929280a5cda682478295eb4d225b21b6f9ada31d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfdf07da21521a13250d839316d7344c69fe488dcad8f4904ffbe10ab9a0604b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc584ec363bb35b72b275a558a734ee4e9d4a901559a9e84ed0222d0e1c223a96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he050da337431fdf196a348c60dca1347a19143ca342d9b61da68dee7a8800b4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h462a6caeccf0b780bc205806fd555a0385e1cea7930f5e31012bce69704d3c22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e01efb5046936911152b0d3f9ef95fe79692438b9fe4ddb564e4002ed49f60e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf692284103fe5c41db8ff940b0f339b6637cd0696a982cfffc040175d25d0b29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd935ea8b781e8473eac6c9779102b66ef3ec698e226a6b11ab55fffceba2836;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf15e4698dabc7e2f6af35290a579b165cdbb720e9dee097fdf922a0c6ede49d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe767b409b8f1faa003792eefc05138718e4ea95033c96d02e6ac327321dd98f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcff214f9d4dc6ec53db202284b30e3b09df2bed75445d978e4e279330e86ea66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0e3d2bd64c2e6b8476eab44c1b34e3f512879a9a68576b5311ecfcac00a7fa4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e5bdfe47562bfab8c0ef834599133e4d14c7a126053ed9a01fe967e7db04598;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f8cc81b349a1adc0be681a6cb4ea0f776d142d46f766aa6510fadd5090014f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7aa0d8221d1604c882ba619bcd3a377ad86ea65624122875e045bf85e711349;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dc4b2bddd00b0d367f240f336d82c0655eee01b2226e339cdd462ef25332c27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4405cf65d312e6e333ca38cd8f1cd5f4caf3343b90c4aff1fa45e86d4cbc033b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfae2ce58e1ea275866e363ffd9b1a030aca249d217c1050f8b06f66eb2d50265;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h169a715bcc6aaf0f061b5e7989c4692d17673dde39dcc8277346bc72047e2c8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b41c0329e88dcef6fa2063dfab232db8737a32defc7c4fd922695252aa89764;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h227bd79c44c0e1d23c83a2eb7653a4c7d46c503a12aabeb6751c5f8b15f3868b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87a15c6b6c9713cec29aebf88cc3c80c994fe679d9ce540d536290b9a696ab2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69508292f23f3418881e170de845ffd9dcf97fe55062b5c6c5d8873ceb5a2406;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21f283f5d0cd95802b59a0b4e9d122113c96c246c78c92a1816c7630d974d1e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1428f03940dae84bc751c4c62cf1245f898a9e0b5033c82c1e7aa5f6cb2c3dae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52a6a18a8ae3bf341c74a034b3c74780be054c3cbb14aa482dc092d708cd87f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f232f2e565771bb09602cd5795efedc19fed152a0d2c6b315afacf0f186d028;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c369b2ff1022d1be2e106efdfbffb34e200d2db6bcc804ce9ed03168f2876d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b49576749a00cbccd52e4e5cfb8efb17fa205aa048b69a8cd7f41a862b78f86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55245de7e1a97e63de0c3efd4f2e0f94d47deea10eff67e1035298eec84e326;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h611422c55e199df109ff2db8d2523ed5e94e079805755011ed3375b0b46c1e9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dd8011cbd3a46bd9f651a687b1a3e83e8ea17066ee28a6cc9724f241aef98ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5e01563ae74696e896e8ad55f755b5175d35397702c3bed990c8fd2d49cb43c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha076226480c213dd51da161e23e0de60739dd4a7a7a99132f5dc799ccc175ecc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ffb0018c052011e5ee41f7b2e7cde5290d4c3604d926b523b3a397353798ecd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h971432530caeecc998b258640b0b3fe32213dbef1afd67e118d34227b3f184d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca2e73e133e849f999d66357a38f4863a5b3a2cbaf3e9ca8ff01a06f7e91b9c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8bb242f601125628c472bf11bfa215e33603b2192be528f5b80454e814c03795;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b4ccfd4d65d51c0b45d357f87dd881ef3fdf08c9d677213c4d6b268c6aa7336;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42d06ee512ef3f61c8753bb01ae2895ea8dd3b4741466aef68facbe7ab5ecd05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2ce8164660f5e6162ab3e619488eb2b478a600ff74ad076c52f8727dead99b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25f40d548dcfcaf218ab3026bfba66e47869bb40fc2022253576eae2a0ccc03f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3de04e44ef0ace35885b2c7e702ed09f23b106c168f122153468d38367fed6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36384f437fffa6c004c519d50ad9c0a82444f370924ee02bec8c26c1150566e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47d51ae33e771fc13ebd6a05ca29d303c1ca389fa2ef36926007700161096961;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ca1b1b8339aeb417de870ee598e65df014ae2008fb647b245e0bb13347a20ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5aee5522f03a2ca688d9622dd81f01b23d672f0ea19631fa29ef45546a50e1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf72bc8adccfe3e3c81bec7eb900c1a2dfba382e925a810d965a68ed8033cd18f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78dcf778aa0cab44af84a1dc68d532faad5c0b9ef621a75b9e376259f18f0101;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha539607da06528d2f36994d6d34aba7f8bed897bc498e58eb6716d30974b2a2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0066b559a1b8cbd2b5a1d0f8df846d9e9e244704ddb6c705086f9118c7c464b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h210592684f30ab27e78ad239cc7753103e3710b8142102fd1c5d929985cc9c1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he796eea31f31d0ac6d9ae464dd39398f4421deddf1a1709f379121cb40107da9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ee052f62f2417f9096e208e2e5487dba9d65400b4ce38b4638c3f4f6bea8cf2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbebb92bd33c1df988cd9cf9132765d04aabc44045a8c209249f929a61fc1054d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd86c34f9ad0fd7c38542776cf249db8da983120daba20a3bbbae9ee091f839e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbaff64460b7c56d111288ae66aeab2083a733bc593be44af373d6d850c4e1adb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fc8929f624163703c33fd76100366be567bb47e6daae166b93a95bbc3387a86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d66cd90bc922410c363cba537c07b64cf2f3ab64a716232df91ad0f1260797d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45703b69c3686ecf9b0a84b2e50621d3ef58bf92a90410d639ed29b867e21171;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb28f93442404c6ffc58422fb422629baf8567661d8b60ef7584b9a54358e035;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc282c4890627d5205a326fb367934f7736fca1df1b1c98d14aef85ef05bc670;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb87ae74cc3164f9cdb706aa392f7b900a1fee7615477a18baaa8fc3af7f2103;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h509311b5dad6f232c64e009e25659be5c1d31a5f7e50d754b0846ad0d1b980e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23c9092dd518f52d43bc6c318061299d1d08af36e5151a7545c0c3e83108c13b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba6866b9ad19443b6cbcabaa94dc94b1e27f5177a2ddf30e196da46df16c96b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54050110ad8a4e4ef42e9d710fd282f24f73a8ff513698a6075a28cb726313c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h417a24edaceb3697c7144e2113abcd03256155d35aef2f80aa12035643606c0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28f2fa712fd7739027242c226f2233a565a35c7886b59886e3d9214a502b3b5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b1814e74a8453a352062d7069f1bf86aa2c0e0baf664cf61c7d1bf045d396c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f51a0e887389e3529444414efd50903806ef4259a3921317da237ce7e5d2794;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8366393443fcf948cd0be2771e9b5b5e2504a95db7795a299efdc586fa2db7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7392de946b38659beb00071fb54ba40de18055e6c63fb2a4ec960a9348fb27b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd04258b9409a554a7155e3b54b1185b6cf3d299c671259688ca1ef7728fa6366;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7c8097c84ab6164a5405e5af332345b92a69da7730f9e6c2f79cb577ead255;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86cc5c8f7d8be0a75c2afc52b3bba5f156e02bcbdbfd9bd5a25f48efd18c1a0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eaeebfae112a6a59de2ca7890949efacfdc7b7b0b1c0f72023704f72715817d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3ad4c295c460ef1b5b8894fd7b36f0306c2aa1428ac58c33febd854f06134ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9f3013b996a69b5c54b4e8d4843e2f7e94cb4c0b3f489f9eafabf814c98760f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h356894fe3e988c7b409685a57342182e739367cfd605ab8d91ba00993960aae0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2f95327e63c8950082080c11967a24906fb591c6174299ef4df74d58c0b5fed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccdc5a468bf873d73213ce9b9083c506a6b09fd85e6684cbc24c29dc676b68f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92f57e213b7ec77933e9674032b160687d9d57bec9da4c5f66777bbc98008421;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc254e0971e4cf4ec0e94cd9bb20ec2549b5954793753c3f37fc8b0dc5fd51851;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfef968c4d8b28cec6ccf02cc06f93d7876faa77b105d40aaa869726dae685660;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43405005439d80cd7672c021cd7b4852476a101f242b68c9bc47125da1e8226e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9daedc42d179d46999637e1dff553d08b7618dc345502c1e974f095741c4cd94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bbff19c7cbae26a7bfc4207dc24be8759938af61767079a5ec393725a1822c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f3d6918e703ab7163c9c6af9138beeb3a0287fbe87420a72582c8f30196f106;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h406febac4ca02b78d1d059b997172b16c66c6e7a9dbe5040a6d6ec698030faa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64b0ebc6ccba725f22777940eb61061c6b3f31e9a86399a59cdbfcd5f8715ee6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef9528e015f3594bf3438e4ed0b04457b6a7a14cbc6d43fddce84714058fcb1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf76fb21d0a069b2706ccd2e9b060f18a0190ed5c5337c2860e03d158f225363e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h220fc94d173cc647f847fcfa68ad029141a115b1910fe594dfcdcc568f098dfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5667174d1612915d126434be989b1047710b0d8510e993b7b16f95ca24a8c0a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfee31f866b17dccc5cd11a198c5b945a61d255124a4a50e5acf7741ccdcebfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61900c9cb2c2fa2713b5c4eec896849392eaacb979fce53b0390c79cd4ea1457;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2390c9865d067d3de0343b9b908375fc1d23e73f7cc9e3ca6e2700dd8c27a321;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4240516ffdba67f9cfff4dc879490927b8be1b4801e937ffc0ce855ee1117963;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h750ea855b1c33c968ad5bc8d59883c7e369ef9cb4b6cedf098a5df740b4d386a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56dd22cec9597473d0c2fc6a236573dca6c4c3faeef9e0375f8e951ba6bd487b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h155b9251b478a3cbd74af92c839c1d90c4d946ce4a1c4b8216cb3dfedbf2f7f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d811c8cdb9fcf66abb38e190b6b65df6abf1956406447d1f066e2196f393de9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5673747d719c72b32dd998659c90e6d5704bc39d86476608976fb4323fad1295;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6396985ca7636b9ee27658b2541e04046db36af1f1bc30ae1857502e4cb23db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf68593700d460b89fdb2cc4e26739e024e16fb852b3bcc5ab5e1971a4d2dd2e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha697a3c51a31119c9161d8cea4cbe1979f33711ce4d5add6cfcdc80e9b38691e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a1781bbc52e66d46366e085b4087eb2995b1d906f38be76f6dacd9b3826dca0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h538df7e310e4253d1057bd3cd2f2fa9ca8e94c70715c75316ccde3e170a8efca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39162e499c5ab7daa24a96e6b071df655371cad6abf6109ec20d42823d6b5a94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfccc92e223cb66516c960db6976c8426b39f860f713709669ed6e097cade9fb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9dd5823639ad78e76d200170361a4a9c2f9b9ad4ccfd80ab82e356d2a5cd3e88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba97395f7eb4f557b09898bc4437afb7f60ad5995a3bc6414164d80afb713a67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2faba412e2c886c9fc44c197adefde927988512837943d8b0b1b32bb28ecfe49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51b3e4b4528f0219407352ffb094134acc31bf5a0e70f32f938ef34dc659700c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha836ed8a8fcfc66e3ec3d762c1b7c6574702bc26e6a5d2916f3ddacabc4fe21c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bbbe1a8a6adf2cc1b5fdee39e26ae707a774c171c7515cec41cc03e542c9c15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he389457e2f6f1e4d3550aea6eff61f100c2d81ce653803ad3d6cfddf5789728f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c3f31af2a34d41b7b2ee4169623809c445f3127086df8ed3669e169fde69107;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cff0d05bc155480456d41b3a4fc26a3e43d047c817bc4ff92c3e0d3c59e1607;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33848a3ffb611e11395548f1d9baa29ff2604e5f1eec1f30bbf4cd48850dc6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77b516ae898da9a1a11efbe14c19eda055f397aefd73c6c039c3a2904c6fbd58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69c203c4b26c1c3d8660b30dbcecce842ec3e89b816a586515d3887f95b25d50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb6b1bd0fb52de3726d243136c1f12ae7350049e6c4d3f9bc6afbae3ccd6daef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h248fe217800bb3e95daefda428c761f5316f7b7509d27e07b765bd00649c6104;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab81a69d0823c69991c9c533db18a7deb0db5154d62dbdcd40b3cc208c7f0c5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7caf35cd8df645955eff9cb8c32308c35d3cbd206d81d8dce300908e77189e80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he142f8226d1bec03b85dad3f79661299dc4bf2efa9879bd09aeb25524fa2a9ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13d1da3b4ac555e304a12b93c778cb90fbae21a779157d71615c94b81efb208;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h181f6818d5bcaadd53cd4e092f224e50827343a00baab9af963f05b4e1ab57a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43abbd9c08024f55078ae7adf6471091b44b144576fbd916704edb3e0683e836;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3ceb282a64f5597e1b942f8f9f6efb362564389abd5efd492902099c71bd71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52c213abd9bb8039875410fb7d197a7667e72704acfc3174228986a4ff357ce1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f2f731cf416ce5f51aa0b28e5619268ad4e5124f1a9e1e0f92627191ba658b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e24b4585e4beeb1c94ad0f609ef4c743344bd1dff4e9a7b18fee2321842a981;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b74513e8831a6d9f36fbfdfd0a59c6e0fb4d7d53f597a685bccf8712e722d31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he677c23283baa84e4ede1ff97d6bec0610570740234a0af0dd96891a52bfdf7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h919857b7c6c17baa604136461fc8d7dda5cc59048f8deaa6c9d0ae5add9fa73e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b7983589e4d5fc8e029fe57c015bea8edf99cfc5d088a3f99751c1e6ee37c16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0d5992ef174d498c1aec773f63d0bff621f29393380e6e011b7f7f31687ba85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fab53d7ec1fd1ce56c76262b793b5bcdd89f02c3642e14c8fdae7a09cc44e93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cc509505f3227b414bd6ed5a687aad54543574547acad9a32dd3128cbc937ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fd520f1dc4ddc6106141aad1b83eff2b394a2492167e4be374770f4065cfc1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b1c6ea401e13354d143226889026e5cdc9d25983920090f57a26e6f1db096a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8e2c2f5f5b9fd7c89e9510c334ecf8362b77f3e2631b3f2730e76d564c5d90e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdf2197488d59e3ad87ba6f5a3ebcd190af459b23418ecdd6426def2eb4f8462;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h968b430fd7db6e2efc3888c738134b0bdff4c375bdb556bf62f077fdff5279e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19b079b998511115f35a5ec1cddf616534d06d67b40d9baf1e0ba18b4e25392c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb0f9e87a9ed6e4012cf2373e5fb184fb1c350be8b6e9b752f51454e6c0fccf0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d922f8527ba2506f8618d9d91f7d764519b609fd544d476ffe72d60d93b4d24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefb700ac02cf92d00582c3fdae41ec2fd41516c03dea8109b01fe6ea26f99c99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbca4e0c349db89cf9270c62cd9c7bacf2ea5ee974fcb93a606ee1cc4f0f78390;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7680b4f8a53d911587b197ce6c1a5c0ee00631046b948b10fa8e1b3c785dc838;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc976fc4c52f24066258b27a048dfbdfb7f649f768fd9a976264c7f995710f714;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd972f6b3e57c1d1f2fa5a885a640fdb0e84cd942a39ac659fc021d4603da8e22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2693188511ec699805c52778cb6d03a0499b7a8413fb9e74a462ab465c227b9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33704b459faf1eeba7f065a497ee25eccf645fc28931591af52eabc84479d9c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4379aee8c40f733a2b09af93ae1fbb660c8b108ec573c60375420a44b5f2aa7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha739d6a67696fa3861c3ac32a650caa4c4e9460002415be006ac15eedcdc4118;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e84e0d57e782fcf7968a3d3a91b920c5831f8fc505a5c089e7c91c449c80aa2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7caa847041214c9a3c1ee72a45a3dafed4921a88d068a7098a24e3febfb18ea2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20c1dbc91388475b382149050db562713722a2a4622126fc2687eb8362697b7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a636f79912274cbb30aab5e45e3e5d765d1a7dec0aa8025413521d68bdf30f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6186c1453d45191b7b9ef88b2dae4680ff2f05d02e1957e2beefb402d3ab910;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37e7df2412db36ec964e94efd31f2bbeb8d6bdbbdae1930d8366eb441cd790e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb419064d0afe89c9c37af604449819f9a422432013265b4408792e6d832f36e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbe04d101ed1dfe1d21539d260a14fa3c43e67cda82960b63dbab287460199b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbaad022f0f63a191b9053d2626f8598a435e5c8036a770e1b6320a461d63f4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d5f54e3146997da9a41b7f1562541a42ca8a286419b3d3b90e5f4f350282c22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0fe76fc2ad93391a44188eb885944c9dcafee0c6b7a676fdc8faf0e5456175d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e03e7ed7c3eb5399a1693723613c064edfd8f4f2ee552f2c0fde30dad570168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf5783dba3fac5a59b9020896f24d17b9399a4d5383edc62de18238ed0333a0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c3b080efca76751250941729afcdb4d59642d144c68b26cd42d3bf81a4167e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b4dd48e9513f5d8695cb5920826b136778c347d860673a41bac6e2ac40d360e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h313af5d6ffbf16feb83765d848612a224a2f53d617f2760fef90290eee3f87b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda9cdca0074aa7521f7b87027b602379b182525728f821c671ad514b7f1059fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h114ae5db0e79054d95073467e488b50d8b9fb42a3ed3b6c48e4f2acaa4219943;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d8abec0aad0676db0b45b87de28270529e350109ac0d97ec411cc622d6c524b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd3f3ae010d7bce35154c314dd7567dd5ce99abbff8fcc14d8ea6cc58cc6e651;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf876fcb842b5b49eb8626cc609215ae86f0bb366ef9a208bb33d3f7165af364;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed69834a7bf16d6b52bc8a13facf2ef5dbbc4e7212a05575231baf11e92442f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97b9dde85b2ad3715e4f5615f5d83e979e6974c3e7ad02ad8409c692347dd8b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7dcf2b3dec7863defb00ac8e3c5f1b96097d50f5e936bf13d1592e760df17b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1690b5f1fdbc2e03604d11f19f25fdb9eccd1a797b1165d344a05d5a2b9298a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13f4e7d4bb9ec7d906f516ac14bf07b0fddb5da157896e9f18e039e32104952e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dd248fb056bf16ffe0469bc051bac060d1b1fc288ebb9abda4dd4e0effaa1fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ba3ba674b1b991d0da1eeab1eab925001d55d31535129ea45f3b665a11f286e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25c68327cb95320f35f50b13bdff71fd3a2c5bb1c338c6349246164ff40a43e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hacca66b067b7bc3cb40582a6e5cf7cbc3b80615a0874e78e8de2c4caa39b39df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3516bb68201d0392730eec8db64e0e79350d927551ce9d5505205d071f5b02d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce517b7f966e40e35aad8a88eeaf44fac7608cd5c1b6b77f99e4c2d9901e2758;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49574d4b57c5550b520b5136e9726eb095ba11892991ff02c6fb7ed4a880d32f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h761fd8d20462337e1be581580d4e3680587e000db09ad786964f8f9da24a6ee9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12ad76888cc6cec709b3c7a946b4457042568ce210a2afd126e2716cc0e036af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e6383d25641f9c71976069b8a333d5c3f48a43036bfe3868d9ca2e0ad7a9c3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75e6e1e2f5bf936caf013fec7506aeb329de6364d373450afd176f361ba47069;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8720702ec0c5a077ab811656ab328a297af3bbc23682cb2e7db6a617c6e07f13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8f8336069e712638afe1e1f7a84e9d6a937a56f55efb93801a79a74431f2ab7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he025d1afd21271091554cec70638ef12737f3525bf22ddfc0c4753bdfe37a1ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fad83c695e134f583c87f92adb8f18659254b779b526c3fc613c9cfb852677e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6acd57bd6507b2582a0d413f9be1ad677ec6e754da52fa4e5228ac9d92cc40e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h863c9168fa239ec09af9a87978a823d5e60dd4ac9ea6bc6de6f8628ce9c048a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdefa7dd128c8fc4d2f1623f00722569a486dab12a56c41529ab46b33ea28183b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb98d540b3c5e7ca00babd4cfbf0466231f0be187f7c080bfcd762ba8711ef77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca1bb021c45f57aa2e767de8e94c9ccec0aebb664553ff2a706c9286ea2ffe5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e562d808fce08bee4a96f1d4da70f5e901c9c10880c02c30ef742a5f02e485a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10279e6df30afefceb96ef801c82ff1bdd706bccc54d483fdfd19ef95ad775;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he39a5e9f110749cfa0a96db856e3ae98cd4b1a0012c61f0147096323233ed9ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57f07ea7af8e4fe00ce74e1aa63d54ce544bd3d87f7126680fd180c1d5600ccc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbd15a0b9ef68dd89a0905d698f05fb2bbd3238650c39530b756f296bf769b5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h316357e301de8c0809a1af2122ffea16a304e9ab31aebd4d2a73d2dbad6ad05f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h552cf4bea3d0ddb57d5e1c0da43d803d10436b078d439ae4577b206e75a75b53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5209d345582f9b3d747f73de5ad70f677b2746a55438e1882f3b17a1c6b1a45b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h746a86ce12052a1e2712ec620678f1149e000bd52a9c746bbb7d95d71cfa80f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9a6cc30ee6a05d27ed3b44c3ee24d34af3cd90a7123ef9cac9399a691a4c070;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff9bb52f1b682cda413656bf0c130a8bc9406db0dc356904c2fd580d3969b342;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he72d341d3d5cc8982b68b37426fed1c6ca939b869088f5cdceee5d47750ee868;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3a2be21d350792ddbcf7c2b1e6f2a2ff4aca96797f953b5951f7a986ce94999;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bf0668dcdc724386cbe736d53b3838078f9661428eef924031414d128da4871;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h232b451d703d8878596228cf5216907e3e757e3a63628370477a076058997399;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2c79eeb0c593cb95dcc4fc30905d90fef1f020b5ac7f0a275325edab9cbe770;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h402abce370cfe4bcf3e18acfa9a12fab357fbd7098c3813433a376f6c02d4892;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6763eb41ad3ebdc72f9e8a59a17377ea34263742ad62db686165555783f4fd76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8bca9aefeb7ed7630f9a224f702363b9aa9777d8e9108047ad3b29faaf3b933a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1743d541caca18a2869af0737121b75b773dbd6d15be47a3e4be88db49b8193;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39fe228fe2ba17f988d935c84df9de40d4ed9d96a63d184abc4a37c6d32b238a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9e7243a96b2a41bc05d07af204cc3dad49cb2a5af168a059cfed55b84f71462;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ba206e9c5b387b871c852fe603e7b9405d38a2cf60070de90dadfa92659ee4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfeb8e7b25d67dbe38cbfa95be3e794c58a24126e4fc92892916eb9f6e95e420;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b4ab37ef0b7d4fbc96b161737ef7bc22e1aee97688f7d94575a592ce0655802;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h689aaaa8bf7ee439bf0c7b94b6a58e77cc435abfe7ceae7d02892bfaf72171bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58dfb35611b8fea49c753138b8816167dc79d3a9a05f7564d108bcc30f4ee36e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c813bea511274acb05fb789ea5f9bd3adc63ca4d3dc2a16b4c6d2719f722751;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa965c953c2355cefdca10fcdc0cbb98138d751a606f01baee2efa4625f0ebba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdedefd1cbd2292b76e0f5d017a5f882bbba4d70c70dd471b820e10818be20d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1495a37ac12f1338535423c41d8beb0f3d334ec48da8053ac9e7d32e18c2a3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac41ab525b90fb4060f31817dadff7b57c1821c5ad67a0f5737cf3e01f5121dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb014d94ee2b3b9208058e5c635db81b0a128857041fe65da0a9043ec3442feb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb205e7cebc0c796d1dff36c1141568d57113d173161810ba7b42c7295b51e40f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc613b4f1f0fff7065b2b210719cd78df42bf72a16ca9eadb52b3485819a94bf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16f559a8b78c99ceaf6d4ecb06547fa37353838c2018aa25fa31edbd5864bb87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5abebedc3850695ab1a47e6566454f6751d16563ee283d6201cd8409090443c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c580e7fe4e9efec4e2810a40d5db862754df185c6b8f08ecbf531944ba7e80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd76c302da869a3a50269f6287d5e5fe819006cb59dac55e29e39990bff4732c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4bc595ec352e76954e52116da1e4ea7593e3d71b25d8f967c99e68cb2d7fbdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6459fb87ec6aeabc9f9ae1d1a818ace639f9910ab08e90ee1befb18efe694345;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ceacd44af07eb5a747bf53ee1513b50d6c4bd4e04382fa1fde700a83d28ae1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3b3d82ef3703688df5ad02dbe47317216580bbd8f0b38be2fb034ed6ba6cb19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h739c051545ce5e33370e9d89ab190578ecc8be431bc6a08f4a8b471de6590065;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4146cf909288345b4b44e06d9ec686f9380d5b485746b89d036f2767142e3a61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d731b3802bb35020d3d04141d537c7cf6bfbdffc694cea0fd78f01b5a39d877;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d25ac6f6e02befada864023bee2853d9f96b530f484502365f52fef4465d98f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71fb9b63232b3752d7e5a9080cafd20ae7262cb1b21bc902d8c5eb5b6c9a1ba6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h692436db2f2ec5e03392aa502fbafdc577fefa8f22849700c24c13af643b70d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbba1952f6a36fc8ea93a3baa22d06241926e3181931e6e777f469b8891858f0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h208b05e72b7d718a37a316f6ce9e17d79441527fd36a2d5c33d01845a6e3de29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h849bc7d3bcb38834478b43119fdbce96ae13231368fb5c0b2d7c9a1c1a61c9e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ac14e8597ab318eaddc8dfca5af4b43a811b607bafa0c15b080a3563e1cdd4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba8fc605ede5d61b099007576791fc37160814a782b0ae7830db435f6a082b3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b684ba6b0736bbb77d659cc082f44dde8f112f6801a2342717b24a966083493;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h138835098724928d1a786fe26c025264ecbe392148c781810cd8cd1a406a9f5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9b73ff4e34d49d6e796cf3fe3609d80c0ce29ff8a66399958f994c3cef8502;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a41fbb5042e2519a31f2c7349fa5e376acf8bc21cf2040663c35968a1b3ce06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddaac0abb4e9cc65cb4b775ffb9ae091c59524eea0ccd218dd387e3f8e2a9c53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha371e9fd68a83f68c9d8565ae9b5cc032368e6ff0860b823a6d5441dc1df3944;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77c8eda0d06c6ba7ab7d62511d9568366304f275bd57e90b0ff0b7ae510ae22e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h495248bc3c8151b8f01a44600cf88f075556540fba4179106ba377c2ee25b599;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf5e70f58ac377dcb776148e717992fdefa52c3952cb18f58ccbc2ff18917315;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33f8884c27c5b5c8edbfc7a2325beb5b0b09cc78695c8b3cd7683fe58a2e008a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5682f45770b699e7e6f7a726d5d7c7c1e414cbcf1c15d3ca7043997b8f78dd02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h326c6d78ff131780db9311446465685806d11b93a1e310410cd53b29465ce926;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83b39206670fe4f27f94ee4301838e40a2c09d4f173cee41d0d7d102b91d689e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3616ce82f52b341b62a0f7f3249abdae40a732f58c8e9efea8f9479357e8180;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he897041b7c36b8ebfe7bd51d01d13bf470b99bf71f390ff0cfe7ea647358202;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3038b530d86a75fe9216355407b417daacda23b8beae124aeaab8c74797c32a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9da83d63fa4298064a131377193b28dcba681adce7fad5cb65fd7d9671983d90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9b136a11caddcb5d55c6c7a8a524967c54e9e22d7f18be36664ee6571cddf7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3ca66aa0f44ab241d1b14c9e8f2bbe447946e7850ff845665151da6f9c35dd6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ded549664c0ddc5a66f5c12aa833c03d37e09e63c2de03ed62d31703a5ecee2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha13fc6bbcf47b410caf320189874f746b939436695a44a5e2c21507e1bc3d37b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha04a4c5164405f1536bbbb77c2308f394eed203b3348d4bfbbed4aea393a157d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfdf9bbe39324ff42f9ea12cdb276a3ccc3a45fa384f1a096e8aff55cdfdd5ade;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40e87e123be93290a72712356f03145ed66475a0551e483c624b55d1c54acbab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32ebb37cf6ac108695b5d52350520fde143de0022f7a322347a15393d0528195;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6976cd446d0ceda702369067315a94260766ecff0de99fa736222792d710f2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6111790ba2df5fdaedc59c76fa6851213db9f579182b5099459ea71baa1d485c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h738625077cb21d954dd7cb1178ce3f3f7e7405978820d236ef77d505b936c178;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hebe0cfce23764ff20be783a35e727d074883be92be55e6d5a175c347988e206e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66d3bc89b0645221e36bce14731969073c313358cf74f579715e0a4ba5c8b8f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h352918fbbde3bdb5180fd78c17d866c679b19ceef92d515809ae8cf6a9314eb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7538a4f9aed67c729bedb1220e73be728d9df1c64d3907aadff10cc7eb55c0b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc69ab0a60f9eb5a18c48359b7188b0313eb7afeff1f5cc014bbf2aa4fd3cfc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc816bc400554a27bec1d2ffce3eeebda498d67411ec3b3fce1d76e06bc253c69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb12d751688dd3bb4c48b94d901beaf5850942cd27c1005952b9913e8030a01e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf4c48814070e639eae33dc6da52c3fb0e30bc96376b7b602d49840561a4669f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba4f14ec6f4e606475d0ec56f080279a2d1ecf9fe593d2019cfe08c926a9e42c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1729e2ba826c82836a7a35b89024a2aed321158fa1f3a07118fe5195ad3bba1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24ee154f96104adf38d6689351ba488fdb1b9302247ed99b9f62a156c7563861;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59dc460f07dc7943c15b9d8612a988bef03c45a046e1f465c033ef60a22a74ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dd1a278782a90c4da320337cae3c207b30145d3ce437a3cb0efc9a16a77f446;
        #1
        $finish();
    end
endmodule
