module testbench();
    reg [24:0] src0;
    reg [24:0] src1;
    reg [24:0] src2;
    reg [24:0] src3;
    reg [24:0] src4;
    reg [24:0] src5;
    reg [24:0] src6;
    reg [24:0] src7;
    reg [24:0] src8;
    reg [24:0] src9;
    reg [24:0] src10;
    reg [24:0] src11;
    reg [24:0] src12;
    reg [24:0] src13;
    reg [24:0] src14;
    reg [24:0] src15;
    reg [24:0] src16;
    reg [24:0] src17;
    reg [24:0] src18;
    reg [24:0] src19;
    reg [24:0] src20;
    reg [24:0] src21;
    reg [24:0] src22;
    reg [24:0] src23;
    reg [24:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b3473a104c09a8e16df9ee3674b3fc01ceb07a8703aa45532b3e55b8435afdcaddc9e6cc96b0f98d96bddf9c4338bea375d08c295d45dd6ec81a0d943939307da57b298445b90267488e60aa19e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e001340f1305eed769586ee3ac00e4a98f516632e1e4405ff31e925aa54c63d44ae9e6efd517d974fe603225f4520a264b6b6761bbe3b8a3f6ad2eaab4385eeeda0df967bcef718debec0d16e7f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb26d9d2a09218843d344eccabc757bd14aa9e036baabd14241cbd30cedc13d92b78ec562473f7e888047b54bdc2ab88cef3a4d707472fd451f15e5152918e9eede56f576f0a923bca2cb2549029d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3f884d554ce55399cccf90542aaac969ba1a0980d3be554f4c9cab38bdf07da56706dc48ca3dbe67e6567a58e87726cfcd71ba75be54fa2660383278b1b4158a3d8455d2d885772ca69a19f3e08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3b7c821b6580775d7beed926c47d0f9988e48f590d28dc463ffc6397dbfeed63d30ea1950f9f5963ede0887614eebb5741cab586dfe645e7e97dcf840b0610a424380dafc7d41c2f8be8a2dfa8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee9d20c39504b482c294ee88b15404ba4c773f460a33b223b8b41618ddfa7ee01a96f6119462b9fd7bea612f39dba03286e8061499a05c44145d783c93cc0feca3b26f57e4ea259a986cc9a2f96b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f3a9e1782dc710d83d46843e17583d449acb5921d4fd93d41672b617561edee3a3a60b908d8a4d4ae3467f0d08430a63cae6927f3c8083cba704f37d5c3d6b563c8fac2ec23e0f507b07360e929;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de864b286a869254be886c95fe59964b72c1df3c65d874b4e7789e6a1b6addebbca946ca3d76de11197dc2896b7ad46d5ee24469b008a26c1be2461a5840a857ae5c9d90198065d6ee17d9d47f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc3281a062f6d6f4bd2364b4dce13db49a8ce270edf8f20179fe0231865c8a835dc637f3a7d9f91c8b2484564b09482f0366840f45b64da85e7d890e14475dc772d9a209e3f4bcaf707e3ca5ca98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14492b165408e70781d3e1bcff3e8e73119c84361603822efbaaf7b1555f7abd0ffaba7b125954e9e62af224dd2cf6ebf2d4b6fb49b978ab7a857def8a5665551357861072745693195f53d3e119b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2fe48ff52abd8b4934e20f653cc3331543206bdd47aee71289c4d222e3a7c56c132813a45e06e0ead1ed97368d5f1687cf1631a422d4f9acf9c2603efd33079e886db8ed22e3420454932e34e8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbae40ec6bc8c52a5adb3f78d458a540758b79951f46d37f9eb63248cd98379e476e3e0f1bac44da2f86dce6fdecd47e4a720b9d249e5cc4a48e4a9e344ff6d7d70b120fd1f2d40ddb0599a36516e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92731e2dd7cc5cfca5dff6c7d9f79a822434c660c6171993dca216804dd4a93492a1ed8572a9229af4b0018f60e60a1709b592fe315defd7e56a840db1c340f2640a3de76feecec78e42a0d2805b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18603003c31ea75320b563fd6e8000b89e52a79f394c302b5210f1ae81586353bee7a13e4b4cabb756d5674a68c8def95996584b442beccb3a0e73996d5951a5e1a76ceb6b5ba59f3a18e1559c199;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d71f57c9e80dcab0505eb10189a91eaceea386ef02c24681d242fe1d5dc4d649797d03134158e8be7a130e8e2111a905052c75ce07a4af179aa8d658b55b4204f604742dab431764cfa9ada08e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b12b04b484537a90f03f361fd700f786955c8eb464d8bb504f5cc0a602fc664934ed24a33b89fda4bd634bd6a7c36b48fb6bd4ab0c72d36c076c49ab6df007f3c50339ec973c84e4a234c9af05c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63550fb43bc9d39df89eb1a8ab8a096cc45fcd0b3781ad849c7b9b7683f8d7da706d3b98ca8706a6c46d2140804c869b6e9d07e5afb3f7a5f96f3a4235443c3d0356f95dec6b9acaf29397b8f034;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c086c473e098819d60600d3f18d76f407819e0f6897d886deba7ac471ba28cae615f657c30221f7038e2f7a9fd5857b0462c0b2d2d792d5fffccafe4772081b283160e2d6b02083e321ce2cb460;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d77c614e38f6c31eabb454d5eebab4c26717b34e3c0c84c0142dbce8da89880a5c5fc78ba50d2390452c778868f8adf2d3a903dd94d3384f0d14ccc733ba8b59087000c0a57722c5fbbfc5fe98dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186f49a556cf8af7a42293ab5723fd8b3c1023682ba8b145d92b671a54f15717769e9c5375dd5d1202155d22b91081ae569355cb3ca55153b76aa829f11776da28516ec71b32462c4f6c4832c7033;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h384c5c7fd66168afa9073a2a449204989c0dd9cf9141ca2bfdf646d09b4c07b84db001f3b073ff2176b042f018599e58597f4b5d9d632388019b545f09a99e7551dde00f2c74faf687189cba5136;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a779a21e5d5bcb2ea192e186a894645cf9f79b0ea004ec8779b1def6b4880907458fe3d3c3dcdb457b5b74b3ce03d5c1fe5501bf6f6fcdf0b54710d427fdc62da83eeb3acebf578158f8ff67a1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27b56e501e7b8b893444901eeeccf33d445a54669845bf0c858fbc5e92b214e5f068578c6779404c3b44ebace70b89c8c2587728551f9bef1eb2523d21b26d3ffe714a44cdc99f45cc12582917aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfee970084b291c0e2599c6fb0b45c0d39a0948966e643938891f92c4170f77fe16258c240bef34e7601fc951a53e5ab6d975ed0daf5ce4c60e985148877fc38c0c6b999ead17c04b5e2b45c8b799;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1cf3e99e006a39c72dfe11df65eff8e4836e2bbff83ac1fa6315978ad040addf9fbf7441dc084e88efada73d2406bda272d63aeb97431956f8cf03d3a0596e6a3bed262a74d4c2d98f6e256ecb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146a134e0665cabf58b63b70359ff26e754e82ba3aae3b972f96182cccdd932a465bf48a2a46e8ae1bbc3010c5786e40983fc318ef1de65c433de2ed7e07b82b0e480fa8e019ab0c97c8e6af6c058;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfbf6f418ca05d8db400de9e2d6ba66115cdd2c684d17db22d6c787a46eaddd1b90fa785a62231c1c628d31df88a3d0d4b9f4b1f3d87a7f62b1185855656ff4ca6c9d840588bc4eaccae432d4f40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d4a6b495167913bcdddf5a065427f64ef86285eda2d07a9aef6282b5bbca182429c60dca7e5460ef4619eed3b0fb1bc8c2b94cffd419b416747b212aeb9c95933ce3d4d13ff8ed59456002d85fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c2d57bb2c50089d3d60ee89f911c44d09deb649b5a221860ab37e5108cc31fa086f7fbb59d60e5715a2ce9502f52aa717196db46c26313c7c36c280dd1b6fa0d634aaaf71c64e476685a1d2b939;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd424857206a64b336d375be8c2d25e95e6e7eed89b3fe32cdf3022f718f740089cdae82d5ef77f143ba15662457e2e070090d33736920d0ef328e250e4d116b4c77f2ccc29d8255c369f3b3444a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123efc79e78bdb23988f8a5def1588e8257a16e12d656921a21bfcfb98b6c20b3446645e4373e3315626d169eafa736b7ff32885d636078283013b48ab78a2429ce7794b735a81802f66f83909df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf47f742ac5e128f253f255b7a656582afe0076aa6a34b9f264422c53f004df48d2e7c79f33f029ba843e5c76b54588419e47b95cedd93a4d732704758d38aac154ae262512412772db4685370e24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha78df75090d291052f16a6bb95a038f120e32d91e2276297fc86b927bf5ee87b47b4d983310ba64e2752c41b8dc6ba84d6e6ef52350c928c5a133e5e3d68eb297ccb20e90e1294e0bc3de3e3fedf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196053b155a8d229083b672a11bc2d4d6a4d716fb35ce9fa4e291bb921ff78da5455cf38639ca17999db7c8f53dd5a168f75140ef26bd54fd104fcfaec97e62e4ca9017a4480fc841d9532f436a30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138d7e6ed315faac4df6f82645ac12e9453041dfc17563dd3887b909b488f51f229dfc68eeba553d320bb39c78fc074a737157fb7b3ceef60668d5f21381f8abec6debd1bc581c4b8cf50a4cc4bda;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e922e0c2652abf91faa71d869c5909eb862f1fe1de8e9550cbc02d47dfe6955759e9a34e947b092796583258a4dc296671883c73942ca0873c454b1ff295d36667a7c5ef291f303faaac0403cec9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd3a911584f3b3d2c285d521f4ba007baf4271e55c24de25703d3152f4113e14ca5497ab4a02b26ea362d618ecafbd4a9fcef7e9bb6a4f3820ba5b3f5fcf857f91c69398c89c33b54ae4d34fc91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d45fde08d2249b2514293f3bdfcce56584caadd27816517f3490e56aeaa6f20da8a3041ac74f5566ecc5b38dc16ae0a803c123107739623df9e963ea63fc7647a49ef7d4d9c31e861779fed8ac0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36560edfb166a496725daa58da1dd46f2eff726cde8fb1c813b051340dcb2d383b7c0247bedb27bd84dcd60eb0df7d76cd2d34678716fd42a50acbff7278f33a22798c9a172fd5173395746a53df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ea9a334eb1ac7061fa8867a474ad44d3b84ce14564aa0741a5febe2afc8d2beb9dc121d1dabf96ee311713a94c5bfbb4052c111363a79160144f07411918a3488926f32a3c2e8f2a1bb24719bb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38042f2b2b0269a27b64b4811856e55d312b36aa67b6c33819148121b35d7940769269d5a7bedb4830225919c128cd0650888abc9d8b5e8c7812bfe041e53e72d97e9bcad52d0bb051aa6e5e7191;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122eb1e6b111ac1f344f4521d89b4acff139ff6c13f62b90206c30d70e0aecd2f6ac0edde01e9471b7d657b6b4fcaca6b55f5b85f79666aa9e19aa0f39e9e5cc521690376c285d4f0d1a4ab7a42e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ed034165b1a5c4e64240efd166f3b0c341d854cd17549e4fe6869be5afbcfe7aa9e9dc45c27fdbc2e463286f4ead7a4f53784ab780f2b5168023d7386b7125d9696dfc3f195cbf81e10e92b7b7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4800f52579f5e1e235632bba43f5883c45611745935c3fdddb4a0a370b8ebbcf1719a5adaeb500fb03c912746626aa199c08f15db7c91b04025d0a12ac9dad68b6961c768924cdfca84b67e539fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1438b54c060bffe269f87cf49136bd0e8bee2d427629186fb027a18b4f6b7ca0d1936df3b7df5dda0c2b9efbcec8ecfe89b29d61b629e852ca79cb40b041523977516f8ae4bab9455b1beb321c162;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b246b2ee3e724d45543620881957e66867d7218355a01ba44d2615cf6be062cb71ad227a6845f7f9120343c759198e248a64ab9ae9e791a424bcb5e36db433939b9104a07e5086930ffbc5ef9b3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cc0c3f7b857167451854ba218ad88fa7f97a97f23074f9ebf83038f26d091187c8e778ba10d4fbb03e204f3795361b22583f534e4771a2f32ec52c59a5a00984457a87050b111ccd063da168eff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78c0ce005aac523704bf5ebcd6698771a391d3cd2819020c9e54a906c7b124523790a9880066465fbf729af48b18eff8156a4a9a0a1a4153e33b727c55963bc02fd2ebe9fc329f4d62533f855304;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e70a04e2ebb8af9e88a726295bd7550b0c988ba833af9494a016b876cf1bc0ddff7e723e1d9f8a4df5baeebcc385331fb8d9702637514c87ba72e76921a8799de43c435a10e78f2d5dc1335a539;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc69c0df4d5124d319a0afd7d615a0496e218fc3beb70df9c87894b24ba7399740d5e3fed36fa0f5b2ff31c83c0e36fe3d83816917cee7107ddebd4f7526bd8e386628f0af4dc2dd5c967a3ec6a09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfeba485cbb013ca2250f8a520d01b9047f0a32ec8776e127de70afa3b15648acb17d58145e0872456037a0150f1afaf4d2c9b5d1ce2a505fd60c57c25a90642818298d1f8459fed6442c6195d383;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b9afe7aac29c8bb0252303cb38921c29372bbd7bd80e2fab5a547e3cdb328e4fce9ee18ad52ac533e95dfdcf62bc56e1b69a3faedfc0ce746419ba09d9451839476890833e286de6bb501553804;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9928145bc41074e10e0ada4917e66c86cca1b80e8ac3e75c3ec3cc765af42f9e58febf0c6395ea447f0b8573002e3aca29a4c8bedac1b97cc5790eff6502f6901720dbb1297751fd2bdc23d4245e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a75d5b78894729adf74e71273ca26d52d120dc1ace45c4007254fd21fd87991afe39d1f87e7ad1898f7dd3b1e14096620dc556034da8e9aa45d48928ed2f48c4ebbc8b5b6d2f2f101b62534c3ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6b84bf7237369e0678e33f3b0a83101c8ed39fb406cd90eb24c647734c21a676e33740f52a4fdb3f1d1f9e2cf9d3a2afd5f9ffe9c17bc21f999eb7dc5568a54234ac8a9b04a066f79a22979bb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12238f610515daab618017c9a5e49d4e4e01bbb48c6f000c8431da14ca1ac13e3dc49ed222b22c420975fc2b9d39fdd73730e41e1e3d7405c13d3d1caf770102a0e43cff30c4a39169fa943917e9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bb07b7e4c9f55089715f1683cf0a39edf70a229b4a5162da922b2c874d8d3e75d75c3fc7edfc78c05aa1bf080dfe3fcc0f740f82c2e925a11a12128c79b3433a754b4053cc7a740d78245fc94ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f8bbb1ceb8236b5dc91262ac9fd9b28177808fdb82ab9c6c234a8b2505f828760006cdcad12c56f43611dea4c6bb3e9e2c545424c9ac760ee9a8607db48d63a2c82a86cdf19e9e8ebd91ea532ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195b3ad330fb06598b56e77bb965b2f84827c15dbb5d9f019725aeeeefd6c83490774019521ba17253d93b665b95343d00877969a822a87ce7b79e1d5f5c4b65ae336b52b2fc1112c02eb0582541e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1280f5c34ae859408c2ea3285352395c6dc5b7ee1c6650ee18377899bdbccba32cefd8a3206f3a1d3970a05a92ed38ec7bdcb7e2ada8de2503050dce4c0a13421a6718426dc185000304f0d239a14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92797f92086314315f55b71d99a9833e2c516be35efddde42be3f4f481dab05874e6a99bd9acee136083dc7474d8b78a160dfbb39a3200706095d1b515acd2cf24d3405ceda58ee7354a558bf488;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113a3dd618ab7281bda297d320f52efde916f1874090da4885a39794c8ac5ea4cd6650b6f6f377e5cca683462fd7456ad5be081e83976ce86682fe3ca4f8b14e28be89eb205cf78b2c2ec7b8ec714;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb124730fffda675fffd7e82664d4ea9ffbd8daf9be08fe1adfd67672948834c5e43bd237008f2ae074c71f847c272b37ab048e8c329cf6cd891ddbcd693e8b8e7a0d0a351a518629759fb8d3abc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he84d9a45c281757b7eb9235fdb810f4917e1fb77fe193ed8ccac9c8fa231611dda603fcdac2d1e6d99dc4a704989e6e8905cc7e019b15848b4aafebe6a955d521503f1c49a59bdb435e0182d2236;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0e79e4033a62fac6e742e3d73733f68e7a8db1d515ef3f74f758d2880ea7be2aeb8c85d77b090d3a262ccd42189d937d4ddf22b03401872c2f741fc2511b09ffebb081ca1c623f51f2c3a920979;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd88fd445c595521847b7c31fe632ebde023e79b760737fcd19aa545a4bae7cc3eaea2a4d7f1894ba98a80cc10c0db99e3e4a4be5a63108b3f18c814c3984b624c2086008d338e19a872d7f9d244a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64e19861f8e4287cd7edc6b0a0bb033b642c7da9b9e6d95419a12a6d6a481850f56d1d4c7d04cfa6f34e97190f282f6fde26768667c0b4a383ad5f4bf3f841deaad4c0dfa0e522dea0159015fba7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41c57bb6f721ffd6a5148fd2bf0b016006b12cc29483bec6f7b5e05604537bda4e34225c3f8f2b300f765d318de0e9a0b5a28f9937741f9cb845c494c844b0ea2d56d1354a66dfd834d9de1e9e1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96701480305faf13f48bff40e9c0b5916f4ef88f77dd3cb137d0c6b220b6db512b7fc7a8505dd2faf7c836ab67c56cafcb5e13b5c53316927f82b103707e7e82f8c66e29b3f01997f218ea6ee122;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd28c8e1036aa2c69afaec0114a631ce9e0f65f94be65fd537cea91ef7ab23b4282d1250ae124cc2cc9050e9388bbfbf1a8c0da36d9be9aafd2bcc11b03c9e3be49a32d9cfd0e60203b09d4105d46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f44dad5be276510da55f77f8fde362c56d59d2f6ecb1b4ee51f50f9578f2bc220f00b98b47675a129340ecdbc245a6ea8fb4b67e319ec742b3514b843ab4520db94de57e2d667bd5425511e2014f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16df2f7ca05175394345ad038824e3a60f73d39b7a4c344122a960c0992687af83885cce6007f4aa3f63e5cc41eec090cfc5f689e9f501db8548aaaacd776d6f255704aba2c723f96e5366809e2f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a2f697839c2a774a1cd25f414e36030843d23f9188277ae3c0d52d5e9d0504a3a37aec13fc5a56d749c2f47af97ef6d0a94f0ebc8ecf63201aadf78f0380961c7ad068b7836c84a87f0a0b7791e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193ff6b166a83599086c2b7243f82cf873ba417ce31903829bbc2017778aa80fb8082028b712a2cf0a093da198989d9a64682b9aeb1d9bc5684e04c704497e2d319d1e667260a9cc40cbf9825897d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15bbb559c314184d431d2a63aebf946b4037f7e7248d7e79b599a9e80331c437b851f5251ff043cfc55577099681460877a531e2ed9586ca87b1d8d54d7c9f2d36fb357d5132b8d7a0525125fc2ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd30538cc8a3e03bf2a628d8d2ea3d328a272fb1406797cfd1981bea64f5eaa9bb68c661123af51814ddfff752f3a858b63a98fdbb8453906e7d75bb2ec38ab9eb4f2e0bd69c8a9882176d6409dce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8908ebc681b60f43458687caca3cde36f88d43a67c111c0f4d66a69c7a40446a6c9e74035381aa69aa77c80e6989d0742225272adc7ba5cbb439fe0e873477ead97749c61532dc05683a49957a35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1370edace903aaaa6e0aac47da9785a5f98f771a60f81fa7d211d26023fc0827fee2bf02a59f7ef11b369a1e47dea366963df64bfa24770c84fec0f9bca83c8afcc93bfea65d142b9ce73d2368828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1484247b299100afbc7a9a5e284fb44ec3374f41511d0cb58626fdbe8217625d05311e1d905b90ffe8b46ef7af3602b3c3de12b08b0a8ab9f9c5f20faf1ce28acd67cc7aa4bdb00b29c51b5c89fa9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7378c2008f0055b3dd78424777dabcfc8ce4723867dc2c33d18374a6e8b8fed372bebf7b915226970fb33996e8f890d09f869dface4a37c211103e901c9334bc17de8bf272badf7804e3877d3d43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h571190e0e35c336fa6bf614afbd956b9f3b5319d87667206e8dab99869d88575d43c24ac80f6780a47032ecedf6b723f1e0a80a2c32d1c1076e29fd9bdb1d1c87097359b4f822888bcae3ab73f6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heac8604cee8809fcc9791db39e3fa631a5a8d2599468bca16128b5ec1064d7440840827b93b3e4e0be10dfc409594a83641e2e90278baecb2eabb3c632aae32b67940601ae1f0a17bdf43a9e29e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107c5a1303c0c567e8b23e13020b7dfd96381d50e4c8f8c9aa2374dc69b6737550e2bbbe5d05213482bf2cfbb03ad37e47f07df793548a971f22e94e31aba1848c5ba642d15f8803c16e72238374b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb35dd0b19656d132dfaceee7ce994c128a709a47da9e5b9d089419cbad9661b5032e381786c995cd9487079397f6fe79b28095c280eb08a19d47b3ea61c782ac79b2f5cc00d7266e9c096e477e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf77f5a4a7c52b29f461ddbe4328136d80f09bc65dac4c630caf212dc1ff3bb66c8ed0f1b889673d90e18078355bfab2632d3901aba3541a9f2624c2f8cf8880958e877efa1e037634e26f8e9e068;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf765b03a9ae4041416285fb38416fcc1f07ebafc9a546ad7e447a72f360ea355bfaede9e182a19ad84c4719ce30792b4d4c8264dca628babcee96c60313072645c59a01c066fea65cf4b5047078e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e9c05fae099b8d24513b31bb5c0e009cd8289af49bd14041d44f0598e2fd64a10f24c564e13e0b6b06ff6220e7be74bbf3d1bb672d2c32e47369c43d34ffb6f6290307c33cb936183a31277051b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b8e6848e9e2b279c82ec7991821a9efaec822f6f98622a9cfdbd2806b6aab6c5fdcfdc9e3161aa23cbf28b7778ac509f54faea638b94c1c514e949354ed8d515cf1c484ad64303ab3add20751ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129eea3985f911a38385eba4719e8a89a32e7c0fdab49779b10beb3996191270ba88b76161d193fc9039a23a9d7d63fae7ba94822f81aa997bff95f02b91a0873a42269c716441fe973bc5e823f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1cafd6adcdcfdca38bbb9217b1e376a683e403262d4d0dfaa672f2c0ac08c55d3c58449b2d259aec2341c2057c1952f89f0a4e78c3b426fc05cdaabaeb5a59fdf6fc59e470a7010ffede4888878;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2189861075cb260531990fbd65d57fb068c60e38f77942855ca708bbeee345e156a26906ba0479ecd43fad7456bdff0983f9ac93e404ac85a100327a52db91b4c7fcc50460cd7546862dcdf9a86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea5406dd27dfd34d7aceaf5102d350db1a48e3250fdecc077f53960e80e6b5c5b56c27c2efbe8d6ea17bc09fbb98bade42d3ef0630c4af31bc6d826401b89e73dfe8edc9975d77adff6003496a0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c4dc37e92369996f53fc652ca7258f8796bb49ce29f89687cc15aa0f829a92551cf9742ca578139e414b0075c685c91fa5cc70fddd52da84bc45515cb1f90601413eb1a9b65591bae94df9180f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e10f0dd30c099605a05547fe4c307a2aab676a775c86e9b68011bb0a3afb15959276bd2eca5b768d842cf32a1a37e9953b1fbeb159e5cd8781642e125e442b39246d37dbc9106b2b0755f70f4b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77ad9d25604a35412f258621a2b9af659b02cf00202a74790db37d4bf1fc883c76073e6b3642f25e30db816e28d62fe8be83b42a36bd92bad2321e8acd5e02d44f0e5a8c1ea22bf548881602a95f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ffff8b9073a489f280e918f71b7f215b62e4a609c2edc4f078a0364b6e94f4a5b5979f91852cc6438a8547584acbe722df2225c75e136e25323cf439cb18f310333c16075a5026aba7e57e5b22b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166fd713cd6bc710e37ce32c5691336f0bb2e95434f26089f79f2c63b72dcbfed2dee2542a8a3e51d76a3aee38216dd2c83b4b174c8a9ea140b67317a8042003199f28b7f8f5527f59e1638e52954;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcc95168feee82ed48c351125492c2e03b55fef11af45fed7d40ac6a6fc782cac813f9b28e007b514d5407dc376cc1801903a2810e36a059b8f12086ccb531622c6fb02ed6a30e651207b43cf210;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f6e1569ce4988249fa3539c70818216f746981122142751cfa9f61525c6366440f5e797172c741de6f3b11d4bc46fcf5664f5e05a5ce3bd9f4c199e9cad4f3f9052b7046f50fa5d8fcd89b62bfe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113245b2ad2946e5f4d3ba353c161f8288b107106d73d6ae64f30a8eb44df4598cfa4666fa88247458c7be89def23f317f3801decddb200c09897b34d0b661b186e1d0be74650b9e38f47da68dd4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h920e457e44c9f9689e68f9673a9407fff9561bed8bd7ab6cce985ca130145904bf8bfd6cefa6fa0c263171768f91441427d9412a1f44fd258cf85370b4f8616d7b5941a50b6d635735f3c0b822ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32a4409346a804979d3da12ebfa30058938d887a1597a1ecf72b5f3dad939761b148e86af5a3d8ebfbb03f03d98ffe0abaf7554ea5bd91e1f94123a3d810a710e20190d4ca12b2b168dd4e3d5e7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h594a5c4482ff2e6ee78ef97b803b9eefcf9eaaf3623cf1dc2f16deba59dcece0ca8c4dae8e6aa4b6206c7833795ee3f13599a23ece7f96561f3b6d04f208e4f6126d3a30028823832bde044968c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c2e245c3860290ac0c994a983dc72b976972b1188f4323d6ef8d6c415a1c01dbe359ba0db1bfdd5a6043589edf8507a8d7191b6567350dc797640a86ecbd6a7b4800d96960e1b490766485e6156;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e25fba7b242f0fda9bafa9d926f50505490e2598e9cfce8899c52d6534719fad9dfca0547c99fb465b323edf29da7da789668e98e2d442df354c046f04f2217f73e0ec5e373ff8ca71ebbc74bbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112c3dfc60e0282d8ecc4275d799efad7747ffd582c2a0913068856527e32772d9a7fd6672e222bb2322d4709e476fdbefdc62fad65b12d30a428255652a63c2d442fede2b27d2a91f94486ab368b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40be454ee097c22617ef5415c16ded7869231adeefe5ed67edabf31a413a1f17f3aaee4c17e204b568996d12e1e2c8dc255bcc2ff712d36ebf205d23ca1b0446537132ca2b4f39a440adf8500a51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf09264717b7d76533d2fab030fc5c2e231bf729495d5d02c2a264cc381be05867956ac4f7cef3ad7a8196c43e8d6668aadb0ded450298c449c61dbe82b6aa8a034e20bcf1066ac55777ed3d65814;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1768cc1b1f09e46a0a7a30e8f1c7a53afa059d0219b0bea0c4d3fd7de5a4c12f571a74a5dd48e64e270aa66f2d9375e9ba1b8f70eb44a8174d4c84b17db8d8e373c1e4cd52da9318d62f4cf97e34b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1806338269593ca38e3bf70f01eefbd37cdd8f94fee17fc46ccb255ffb965f003adf224ced8440508806605f2bd7d22198c6b9a0e7b31cc57861e1ea0eaa0600d2e2ddaa3e9b30e441baca0537fe5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1626001e07d99199546b3d529d758c816afb7554b36235fbffd77956c7366632a7546f61d26a055ee6a147443c50ab95681e5c6d11caf5dc47031d0df8dd0f67203fef194e395507c716ea2aafd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111fabb6d0caf304ae2c95af5abce06d42a6c868c2bc45dd888bdabd009a1f4faae88044c445e26a513bb11161db32ca509e1bfe893e23d695dc969564429ada19fe383d0c0bf3507b2cdb0a0a92b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf86144cadca1aa33d34b43dfd26180d1ec2d4235e74b157a97a18ee4400aa363d1a03dc3ee6436854a51d564d6bd1099204ca23ae9d95fd3d2058d043389e329f5faeaaf7f2299000bdce9fd218;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0821bc43b49a7f2ba7b4c788b2f0f0a4a7b8e99b78d2cd1198e2cdb7eaff3ad4709960d7cd6fba9bf2878201fc651febc246b52540248b962b81004f85cabafeadb489ed46257fa71bf6f07650f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd05bc26613284516105ba6f9977d3a24882aabae306abf8f11a5b7d62b0b8e11471c927ced1a6abb8ed3913fbc21a8aabe9ab3e0f09f8cf795a038e793ce7a189ad3c5acc7711b9c7c813432744;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c9527ffa4de7801d592060a39d8d205b34cefa9b98979e815db91767e27d72ebc2baca3703ee960903d7d9fee0a6d6b62e16ec6c2e2ac6594b667ac12bf52a42bda1266d9840564fa5a574c543a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcc5ae2a535070b19e02450b20ba1e040f638def5d137b5117f207df3dbda08571ba20ccea5513b07cde4fdc2e02c398ceb8926617c32e091e76416cefc441d616afa963503bcaf2c79175184973;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf9b9769038813a42447e6765828a470511f87f7bfb2b507c3f8679a1c16a0b8077b5ddba0410e65dc70cab423781b61414c8b1dc90f6ae583064275e5aad0e8345446006452c7a8f9c55f3b4af7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188111f203c3ebcba72bce7ab8e655668adb282c46144e3a3fe45519c8f207b1d2a17a48245a592fd15d1a91f92fc290abff31b5f8159dab768d556e0a89f91eb8976b9fdfa9214855f0a5cf9bf40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habe9d54420bdeffa03ca2da85c91785676bc82ec7c2f7729d49472bd901a04addd6d1d1c4dec35f94f33f5b80442687566d2b77d8d00d5baed1423ffb193ed7d1e0c99129151335002d3dd9f0284;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b30d1e039b41b0f0dc2a9257f007da0462b81819cd42fbe086eefabea9a354b70cfd03215e25eea3a97343f60543dc6877a41577f8f83bb41cae9d3a616af60682e509c0b13c0d460ba5d5c5f50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197f933b96a13df2edd7781b34401446b14db42c0de5157f80a05146d232a2eaafa6ae64941c3521004e9406a255e3459f8f2e2f27c47ee1bd4550b9e1376e431ebdf9ce9b2604f47fc9ec18c0ab2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ac1c5ee4f319f9d42f82f8ec818e8233713bfe7fab4a33a2bb23a5593d34d9e140162c8cac9290941cc42ff5a53f3cb9f83f7325163800b63bece73d607861ec060c23e49fafba00e84930e6ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103fcfa9078ce660f94255d5e73e2e19c7b8839bcf575fc5a26653e291935a2fc341ce352b89c1e0e2e036b144e75ad61b687d1fd470394299c37b81b2505a092a431d3d9a8d079336f357b4d3636;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b721bf5358ccb309c36ed9105504c972d0314cdf2bb5d20037c11cc1477887e59734fffa15e2ce29ee420ca800309c5b391fba1840dd1c72d69ac0203272a0ecad23fbf3e2c619ac9175778ef4fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f8bf2a5f6e28a6218e8c9ee0eae7ddae2b6d3eda83064e51bcff7ae9fc3a47c3419b4eaa1b894b657ca9e35c5fc2c1f63a2f5e0f11aaf55452e31e226534a25649d94f955a4b7d353f70352eba5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16401c3c3ef4e284b4a83728ee9e60cd2b6d5c6fc99225733b0c40cc9bd65ffa06d29fb53e40f8ab9cd74a1c158248d6a214feeb71c286ac60c51339d4b198e5da91057373139ab0dcd6f7857d07f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163be19f6f82911c13ea6d563ac0592645970a9b161b5992f82e95aee1126a2b392ac5f6c3bc04afb2f7cc14c30c6bc54e8e5a5c5ac1ac1dd97f2246e47d7cbea5a8a77aa6d80c3dfd3d435168d34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9dbfc071752dce2515415e490be1a75fa93a28ae6c0fd70581d61941bbfc8cff6f4f0b5ba1ab230262d00d434fba2f295eb5659e3c2f81024118c44e32085ec5740e87a1f921182c0affab4b1d76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9016770123e4122197599063527672e65e54d7601400f1c16542eada6234473ed27e62d93da007713e1833250c78eb642d873d289da2df9a2828c4c6dcc42cdf1dd15a7d17fe4941959071e0c2d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5fcf2a0667c49db94c01717243b8fc6e524957f04a67c8d81b9277b53861f3becb825f8610c2cf559a89e891b69191dc3b63dfdf67b9d49bda186ba080819f0e8bab101e99f11216986f50a02fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc640cc8d3156670a543a07da3d4f9e43dd78dc43d2afa839bfe3f2c68f9c296ab59e1c81cda3ee143f8faebf8b21b23cc1fddbc4a4c70f2825fbb7a24eb74ba9a92c053b4a1432150443096fc5cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1577bfab9b58a11482e36adf981b96c7ebd3d8fecb1d64ee9600542141bd9843b8863b27dc88481c015f06ce6085fc4847b2012a288407a305a125ffc1ab9e9950dfcc66c3a27e2704081ad427a6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6309b533f086cff154a496cef9cfc12db1567b27643d4b3aa04e80a0cdce4f52047019db74e58df9fa29e8337c5906db999011225cb957e185550ba701dd3ee2bf3b01758a1fd81d73b48d3298c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a81b4bc3d7617db479065727ae5be5fcc115ae71187bbff4eab924878143943adb656da09a51e815ea11b465bc26ef04f43460cbd667e1bc1455ff21acda6fef7d3a940cd353ab2a12e5335db96f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4cc4a6600572cd20b3384e894246cc70a646d255c03eb720cf1a14a3b2a3cc12730f2ffd79cae73d62e59ba734e05f4142d172ad290c5a64fa460f52042873de5ebaecf3d0b641e43658b4565428;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17debd526feb59b00b48320d3e1ae30feda965004e603461084f53e5840f346213806c8ec8593121d2f37313a8ae0fc54fd716b0a651c5a5a7d49759541600668be71e9648d241e1a7265c5814d68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc60f5724250ce4455cb467de242457e257546606631f267978b3c53a4976d813b1db6ee0c25ef43415df389079f693efab252f41f1f62454f254464411eb0f0deec8caa7778035d7f68e67085ce3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e25401ffa1b9640202b893a1430704e9358b576a473c5ae81fdf91b2769bde428c04b43395ae4a393d71012970c392d5d980507712ce39fb55db8114ea835ecc91318b079fb5f310bda47ef5e45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fcf1cf037cbf3ffb896cce249f45c39bfcdd26a359d59364fc33e865e1fa9b46443b1588bd368c06b2af55a81c018e50c638278e2a0718da2081fbb125733329f80237b0556bf13421f1eb23bb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e39420b098b7f22b6be49dfae1314a9cd70c1c26d2721b2cdae5e851db7e967aae5c95899b89a8256d8c8e4726c55bad2b9618d347a7eaca85fe72f7ae0c11fa7d5aaa31debede0785435c6c104;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fd01a6e8128390eca7e05050fc79b1fc0ba563c00c963eb976daaff04ccd6102155360d25a5c70f72607236c000ede6c0774b251a60ed7e256bd16343e48a580a5cd3309aa75032a09d2b5fced4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h277cb9aaa5cae326db3dac542945e6bc2ce29b0613279d51718c90dc3b37a09063e21f43e8ed9ee82037c6caaee5b5fb0d12075ba8a4dd529db359a2e2823869ece3ede6409db1276f289f6529d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65831666e1c0fb1832302e1422a2e77c223b53238d9b2d25feb253a1491dbbd8e4cb3846bfb54805ac26c1d63d6cfaf10bd0930fd6f44c3d74139a8efa20d663fec69e90b9d7e6328dcaefc43cf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2aec723f095d6fee3adc8d6a24461d767abbecd2a9118cbc11d37509d77ce874853dc1fe51be252024809ab35d157e5acd665f3099e161f976a21e7908215211a7b32ccc666c565f2f432e7eccc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h811d2bda25f4926ca66b7e081b0a5cae5eb792e89838d4e02bc0fd7e46b1c3aafab17cfdf38b7d128ec4a3aa27041742e97bdc71f8ccab034432d4a161019840887250a39a1b6ec6b9ccb54bab1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163b68ab644d87f2cbc4aa474b24aba73fe8521f376fbd65020cc8e9dc141fde5ccbb9e3e42fc367eb440d0b594f821878da96b1d00d1ef0864b580bb867a28baf778b5aca5bc26624c3b96872da8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa3127510fab4d908720fe1adcb1fe7a0d6cb0114898eb9ce7523e9f9a2658a2d139e8bc1a9a39d9dd93bb30b7e5ca99d4b202392847914a1546041d1462d6463d27e294b36355f0c6db541825d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1486899f41e2a71c14198632944629384750e79ce1e4c7c8ce72aeff2a5e595397995f16c99c53d1442c3fef05b1fd4d47387ae4ce2137aa026327562b4d13851347784c6911079d6631f1e52f41e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141d0d9979d45885f40f964023539f6bddcfaab92fa6cbcee1d8e3bfa6d9667b8e0374674c9034ef259c3e25c1c8009ea893a1a986e1150d7c277dbaf38c34070d8dc72f455e4c68c951177fde07a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h218a0a5b7d0218e5bd585a502ea4599b63c3a5c764e6d3e30af2cdf93932e2b75db85084593935f786eb8322c1803465244986f6b6a8256e81167c853d648a78ac79360636f17f9640dadd07dabd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heddc569f0ffc65df4b80832eac3c279b47bba0dbff2a222906445d639420ce747126cc19c081846656f850ae5efc340690ea3674348675bea433234ad45df137f75c25acdb299d1d22bfed852148;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0b5bea4944712c2f7949789ae8e794a7bbfd1845ad7e5a555d3edda9e1b826bd8b2c1ed12b6c2509f3ac42c979da20b9d5a4e24777c031a7c78f8920233724ebbe604c1d11ebdd174aecd091fee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc0294e3f61c50b563c012b72d2cdbdaceace266741232058632e03ae64b8e2cefc9217bc840d6bef73ef66451f6ef03ff46f0e032ec4ef3bb39cccc0594f70838fec53c2216306ef7b9d633e3d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee3978a2e327ef6fc8312e271e6134907e7a6043352dab2730ff4b03f015c3ffa8e6facb858f4cd53717a84db38853db327d134d80c548b37ba63d05c50d68553be32633d91c8b7e4f813d8178e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf903876fea619669deb8e27b2c647f46b119cd4e4e605b6fce5973a4036bde88fac57b9bcc7e0245b3d852fc07330a8978e2a1c32f6e655823cd95d34b237ebab493a0eba8744de3d7f8f0b1e885;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc90e028aad5ea0c11018b7333460a51838ecf548566c9b2bad2ba2e5ef2b6e973324e503f10f6e19021ed22fc85c2d51ea6cdc7a2f9f6741dadf23672f33c08bcfef5811c05c678a625703da801;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cd5084f7a2db036cb1dce9613443fb7ad5863477c7aebe5a466a0489c843fa8b3a946e869b44da32c1f22071c365efcfc1387a44e59da0127be87d3f348389337683dffa49fd8312ad4a60f7fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7a3eb0b598ecbeb25d78d683d624f55a811d2a05a206f6393e6b9a060540cb6cc627c93fddb38fc2f462d543d4db55289d7f40d6ac16f0da383e910cbcf30071a9eddc60e1f64c842c4df162b04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3dfad45f77aeaea69722709634cb65440165b35c03c490b7fdcf347874a44e87266c88558b95d90e2fac74620f442cacc4636ecf0a31d3339701430cf2d0657380af011d27b1e459fe8aaad72d3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae2c742447b0e3299dde5d2895b0e864066a5dd55de6f9bcff74ed6d7b2a4653e190c055efa1f8d1dc15650263156c33b3db4e2dcbc42abd6f5e563cee94969b905f76ac2fd55b4a4f6afbdc3b4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1792b743dfd8d43bd57cdb6295469ab9d0e19908e7367db91ebdedc1e28af274249a4bf727b892488167df6b9475ed60d8c1b28f9fee0470adac9485ee3e6ddfa7eb6a529b1af67920fae20421c71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1477f5338e21592760f63ff429fdcd3c1f2c9772c291414a56ba2d8f77466f80341a9134f8adb1b728c7b2cd0fd2e6a5e5df10e37477ed3511f3844d5be3819038b5d890eef76c953bf44cd20d6b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h540907c856c2806e7858fb80f6db22c422cd2e559b34d8306f5c8cca7291c352a8cb6d0d0fb941266070cf3f44f225f3e1cb1267ec62a9318cf08e3afd564dd4fbcea4976acf8b812497a320c616;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166e82649e361ba54a0ca63b6675eeff0c8b21b92bfba2c997692e7414b8033e2e60b788f026edc643c2e58ad032bd85bc7f43364b81b30438a315d584efe42c6bb79fb9484e9aba318437ed47302;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7462c08d918f23d131debe79341db3b04cb9bd467b9a2a46474ce164e77d669218900a48a9dbdd21a95c075fab0613463abe5be8e163b8a2dfae90cb4e22ef82c10e7dc3fcdd88dff4941edb558;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61c8b80e3b673ea8829e0c6284beb8ce70f65d1aa06527f0503e2b5f85fc1093ccd450de7fb6b21f8c78431bfc338b6d01781bf5a84a5ad8f03d6371f32edbdb9e6d04db1c3ba6814faaef83595;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e91e849caa0cdcc010c72f57054228921fdc2087bddf9b0e65187f2e24888dc26518403df312947ae982573da2934b8242a8d5e9229a12d7635ca1cd9610def5c5b6bef27661d2517e10fea88aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb269a0359ca5b0a15c0f1fdc2510de8f48260b9df0b2ed50f35c035f20d7d40734d76b7028534d325141b1ce9d7543634263c4559a29aac26481e006036d0a7031232ca2cf4afe02dafa905b9ff0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38035dbb1773027ddc46e1b1d467a84d4f7c830a07255771effc7f27283150c62c4c989c2cfb7bbd439d4e4984b05f77195dac1c2b24ab83f09c1b944093ebfb1bf2a7e37a7a6e786adeba01df3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a952b003b9085655522979d61b4a29d691e2545eda864b37a6aebc207aa80a10364ec215a9e2f92ccac7e1a0d37095549c7f194eaf6b966cbbbec96bb8dd1a4649e2c0fe7c1f9ed9c0d7c8f76828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ce050defdeff8d1fc994068719cb6e470bbb8d382622c7df8e3e166b2eac5a31e4352b895ec17bf4ce0ecbe1cd7944f762d2c5f6bfa0e46ed300ad2ff729b9054dbb55124d11294ae673038f635;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c9cefa765a9f2b10da813a76f680a81c53910e10b0e32ade926909bb76dbed6aa7601b52ea9d3bedd6506e212f1ed75dfc77f2cbd163f8d4c277d3b0479ac6824652fb72d143bd1eeb0eb024307;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59021b7c4a259d49e2c65ca8d35740de2fef0649c13d6cf19b821b3ac1c2cf468e526bdc820ae9243e69453eaae78b8c43e688e9101de537ed8d031786f99910c84470b03f7dd8a6176a1e6ccc89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1425cb06b157d07fbad229b2cefc8d28426970e95c6833ebb6e0402785a9c86b7aebcbc00ece1f174879eb668dc7cb8745f22f5ede29c295185cef388ca0bea47fb3326b4daf0cd812193fb3c1411;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14153925bee9254395928c734fa77af26886d1f137ce4be6734b47f115d96853a9496f3b82a32d1cf3f7cf8dc24d6e4755566909d10a18f18b271b1c1fe592604626252a2df0a3fa5c8c969887157;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a824dd1dac7aa5f553fbc7331ab6e4636eabe9e73276bed7246b3da7f529ea938f36797cd962c30db86036c9441c46ed3bcc781d07f448361c145b0d482f8881ce6d50baaa8be87b626e0f80ba1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d26b2fd22909e4ba1bea46edeaa33f14f341e16485d69b1c0eb8879e22cab068db151464273598dd551750c09cd95abaca432b4249537f3a784b42c9867c32e08d23506b2890a16d7145f4fd82fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb54ba94b33bb23c6e55c57368973be94b11c6b7fb0f5be9d5db8a49f8850857f3b254e5af5d886a87477fbcd30efd63b9bca38bcc9efcf85832a3eb429e54f59c370b3b986f8a01b56ab7aacc9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa01615858bb3c654b829247f36b0c1dc0cec7a339543d3d820ec1c559a38e416f2c03f56e8c2a5a4326d637ff9efc7d6590b949c60b63d9cff9fa889e33f0b26c36fa2e98d4794b03236fc6836f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf42a489142880f2c760fe918362fb1f5a73ca0bbb58ae217ea46a0336e08da066a38957a55ecca4aee8eb29c88caaf80224e7d86071ea5c629f0cab5300e499609d3f791d185d2f693deff1a6e75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5480c132421eb8f35ea048c224dd8289f641bd0e632d17cc8c36845dc60ff691145c68717cab79f77322cacefeb8bae3877eae59a72c4d6e038bfb9a1bbc5eb266472beb11dc5ef44161124aae15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163c6515a364065044def0f9cec5cb6605c5dcbaf17489f84ac5526008b20efd113a8ff1a24f97ce123c0593a6e8f3598a86a357eccff08fc3ee003595523886352cb9155404afbee0ff62e859055;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d61216c164128c0f86f757fb1145572126607a1ed74ff6b5dfdeb86ff5e5f61de602c802f126829db1a15dc95fa63ac064af7615a552fab526ee9769de4bdba66414f9f3a906e3ac92b05615a7bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5debe2ea840769939e4c8d08e94e18fc0c5791eb0ff2838d239dcc6c74e555be39fa5240b5a13ef5f3c08a23a2ebf5989f3dd23d1673e4490ea0b3f5268c8b8665e345d40c043b86ba301c4e56e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4b2a8f9b37689be8660fe2169d2423ffad7a0322225de7459759adbd4d6596da258e427c397a75c899b608fcfcfa3a5dedf93adcb8af40e9b5d9deccf90d8efb330579ef776080dd62360a1150e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152379d15aa719335c940b78559e82ec75df3c63d79cef93cad4ef2092014991e657acc09d55eaa861da1c77003aa5a70a238bb5f4a396bda8565f7e09ee3b5c89589ee4e73f40098729175da4d71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a7582d031c199d367a52e0717b17f0fdc7778fa4e933fea892d3a00668bf513119620520857438a4393de41804a989967ef45aa60c4af50974cd5bbb0d5be6b165abb56b413a8d1da32ce628573;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdee10a8181e0309d935b4de661eb1b618053f2026038e175800f00a531c0c67bffba90039ae0e65cd783c25a7b77bed2cda3ff29fe45114ff406b4f615205f7c6c2458353dba0a58a38530c9cf8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ceb7f54ed87551f9c47dbc5602a8cc436b65eb41240a93bf5d120bc9a75264258443ec70e9e30f8f7da0bd10fbd7f1899ed336f1927c32998cff4ab0d673f122b901949343d5b815e566450b942;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc15210f03743fc2fb2e8d953a378fc3b4ce86e72c63851dcd965bc92d209a06a0a719962eb41f03505eeef44fadd7a7f6f1e063fb24970d23bf1e956d34ad598946c73bb9b0d979a8283dcc0788;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h959a93cc64a400e5dad682cbcd1dc8af081fb7d343e9edc917aeac5ac37daecbf4533f4c0fb24650efaf59a1f4d83042ab01718f415f36a1ff6c3e5742956415c07e88e036edf38c9ed38e6e4fee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha90b070d6d82ed9810eb675aa7063bac211f9d15f7bb0506a19d9e529fe93eb307ce01e042f1e8369d54ef62eea0e5bcc55aafd8e3325cd04cf71494ba948080cbe43cf8bfe7fe024f06f739ca29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1905589f159c0c545fb9ac8583b450a2e6195a3029bf0a82b7cf4c43fea07f15a18b3a955e411181e9b85d325cf3dade7f9944981fd3e7c34120d104961bb6a27b56a451b4f2928cd9d9181682fed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8aa258b51eb6aa2f38700c2fbcfcfdd84c8610c95b4bc876bce98c7a06bdea57865e8deec8652259e4ca6a2c7f2c383a05ba48a94d2bb8265fb01c029cf34ef55f3420c217043a0f869ecbb262a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2051ee86cfbbde883baef51fa08c0dc394a8af1016c29f08a2ecc00a44f862a79e0b9168c63447b2b52ce3850a78b6d81791f34e47c83efc19d60d0830a4e77b6831334e7e8e5008987d7acfe7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3d9db8addf40eea138198338ac99975911a3afd165a01e06ad9d0d4a23eb3f2cd2115e3762a05cf93aae2b8dffa8bb863aa9f5349030439f98aea753e1a5b1544f38544c4843e6d30db644df226;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1125bd11a41d16455db3a7aee5c87fe79294b5cd93cd272b9b440b6ae3df14687e8bcaf64f9e368d6addf3072ae02e1cd76a5834ce9e5846b60df309caf1a63d2cf1f9c55e12b816c9e956f3b5a5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e97479557d5fe773e3ac398dd882262e572211ad2254aad517d6347088ed6de7af1055f0df8163d704f0b49d84b8cd607dde2d57024e63e88402fea4b2b1e0c8919a0a4da6f536a22ddb84c150af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6ced791c841f1ed43ac4e421180c76c09754c895bee621e71697cfa423d7af1dbabb2c85e99c18e92ea0dabfd161fafda72184b138356577794c7c45d406fc434c304adb6e24e94123fcfd1b7a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0ec18499ffc302e48f543e1d19276d1cc27741275d6145a4b7d1840643af8e42922ad7f40c8dd70a030fba029b5aeb7062c86a52fc2da4e72e60e374760a7af31f407d7c53c372344721217080d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127cd60ab8fdf127042c6cbef79989a012f552158df17b07d03073ea815efbff65d3282f384059513688d5747a016ebbf4e32765412179af10510c6d31514e21f9d813e2b8eedec24b7e8be56e8b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1939d3a337e2d2112416082d024f45ea81a8fa1196b58583f59d3011dc791155bb1872f1bf1fba8b51fc2ad057121c079b237bd4e539b539f197f1eea2470e69dea95dc00abf745845cd84a8c0b86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169a9cab5b28e4312c52e42ad7e92ec1178e764482c06f7e2c3c4b0dd26dd8988394b6499687d60143fac6fad612467dcbe6fe37be954fd7bcfa94cbd58b19bad5c2ee9a0d2062b7b85d01350195d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddf060a00145c5cc35739f39c70aeb696d9a7fa6767f735275ff2f0421ca3c9d7297e2cb2e963d8459b08b6650b3422098e0c7f848a31d9d3fc6f3c44ad028226e065ff65d13350f020a7fb18793;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d13f734852939282cc6d9d81bfb3e56d1b9495860a455446850255a75d2d55c7fdaf11f1d78b489e463462ac0b268887ef14d94c98ea5678df308421ffb7f5e0691a58be286e9b91ffa1639e3ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d888d6bdbd217333c06971ece6092a6e6f34e3c517576cb8cdba1e2556a121d9fb285e0196205dd799b656a9a3b001c4c9215fbc8fae83782dc6c42857b8c63168f5274867424290195a761719;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc03210171c30f8a39a273b9af308344e0ce345b32c49dd0bcc8d32c1ddb9e041ff458ceed5678c532258b93edf8fb4852cd7481afe50076d078af2fa0bdec316304990102bdfa4b94202bd6b7a87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ff4bda5c8fdd5f513f10f958a166be4144534be94e2a8a4ed44c6638ca9eed4f26f131be467049ec5bf699f914cffa58537a4dabe60cba7d1091e3931d30e297d326963ba5d70d44d1486058f56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1256a1b93f7cd35eef1f3fe8ea57f3d4fda6b7698512a964e6954c684df17c6856978c93f89a709565162f72b04ef41d4cd2091dcd422c4111cd5e82aa49ec81addafbf5cba28682be152dbf9acea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0678192846d96920aff7871cea3063c69eb26de27c5a4524e20db15fdfb33dc87c32365f584321e7666626ae00520e03e4ea7788b1e319bb1c98a53dcd5dd28f5748bdd65f024ba1ff411ccde12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a57275d8d473feb4fb2fab8a0f9f111e1ca1747e0e952bf8545016551cdf7ed20b12c6b49e5383c75f1415ee8d2e5972882b92b176a42915d1ce7d3a5bd0d346d3f9d2d12e2d1cb0bef662901e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h705dd1d03be866876abad41ddf4df0401a76f6676e481de2ba644887cf4863a1fdf684f00011b682dc95867728da548e8bc9b8b140dae47809bc4fa353baf7839a152c0c740c17b8b82bfcd851a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a2424525caba1151e21dfa06dda67ab538a3981d23790365dae11e8c26663c0d1648e1dc20f44f6bf12a1e77327a64f81ccf4b3395ce3d108d71d85571893252997d704e85f392257690cd3a421;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1095dae97cb4ba2429c9dab43de81fc3085f13c7b9b2a592ef4c0d79b9929c9230909449b79c2f9dd573866a6e17f18fdb6b5f6938666e7e41ca483f6d2ec0da4406c58a39bc0117f5f2b1d5b6403;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f02c140d49f8f00a7e881c37099a333e3e5b318ddc12f59b863da4c68a21959bc1276528502f56a2d19e8f250549926845765e2249643fc93cd825ab9b430763011337d4de563f58f4d43ed4927;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b703cb13312a90424407bffac348baf5617a924a2e2f93b8e8087764345fdf5a6a76358ac1b1aecd6b99c13717f1f895e8646ab29c7b58af4c9c5a77a39ea0f5a0769ce2a61a622d009216141658;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2924be7fe9429a57a961d15ccd3078f1af7cf78c1379bdf147a8e0de2d913e8ebeef4d54e10329727e2fe060fd30bf6abb93a94320f61ed46a649039c8f49542eb02a251ea6ede86dbc26b6346f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1256538862765ff7c4a18d472bcf38cbf330c20b835bb32f68a3e35e0bf9c72c41d9b18f70740bd7d949b167fc5feb9d9bab93ba0f195e249ab03930a31c9834f2a530849610eb131e4f17a714df8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122ec0fd492293c074045c71976b6630f54855020c8025e3cc697b231e0bf564d513834be8afbd46f445fb230c7720cd42ed758d80e38e09435665e23a39619aebade2bf0d1db48f2e92ae62514cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3e6ca1f2b1fae3d41d190b55d5af369d522896231ac0f9e83bcde73bb6fa683c5031698eeefacbdbaf64c3bd1fb5968105d7b075b2d039d1b0412475d2d731bc12240c94e93cd8e8d88aa2d7f61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1a2ba793a396cf4d345b3fbbcba69d10ec3b12f89fec5e341a66f4760c23fd4a275d7c9ed5176bbd432e34954c4e7225e7ea3676785d33fb6423e399712f9e655e9a6be999538e8d525c7bfb73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heba83d7007237d3d3a967c12296c9ee69324df08aa8896dfd399201f74298c00e3f56a59bd1cc722ff5211640a4c7c04d29ff83037d4c0a82f4c3d6ee016c2081aed6c8ea71450f766179bdcd3dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197de166bb54e33f2ed9df8865ab25800a1822a69cd889af3d2c70edff46b33dff729c2433e07db0454aa5b8050bb05791d7d8c17c5eab43c05fe1df8bc380ca44f2749c7fd87ca91e065c5bbc1e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7b995e19bdf8ad6a1c31052c7dbbabd78a5aab3755c53882259df50970b70afdb63071492e7d2bac79c45bc7e09aa34c9015cb9eac2e3e4b42df0cd03479389dae0eb048c2f750a5ea500a667d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbc58669d891efb6271c48db48944a49e0efd1fd9a1d498d728ab0e2743f7cd0926a63c60c05a99bc79e7359bde536d5864678bc638003528a1299902a1bf6291621247c366178e1760a29d12b1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb01fed595f5023f24707becf8f7b624e02ed5ee8eaff0571660ebbc365e5a88fe4e4e32a843b59a3e72f93ed7b4f6c8a03a87b29a6f3e5ca4f8e7ba7c5cd572d399ede9130f4c9df2b52ce21d1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6895f6e5b45c58ca528c8e774558589c6ecc2c4e70f5b6fa97878483c0db5497bfbe873e25e9589bb4fc2b864d0c3443972e131a60b8490f1029b20bb72e512b1cc2af9ce01c37228fc4032315d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18269f2984499fdaff53da40b16b2e8127bf86df147da05dcd71aad7e03520e665dab1d7e584fc4200439bd479bb6d14cbb6a8dd20487370a2db0d8ccfa5740f7127860c16cdddcd38bae60b9affc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b60929082471e91a5d7f91d7b5460fddc218191c9fc54fd34f1e5c6b2f72fc7c0207630114ab98132ab48949adaf31f9fd98062fc7e54e1108024b9432a021b4ea2c53ea6a11b35f6c9d7916871;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7431121f64c1aa1cbdabd9e59822989d84971ed27bbc35d3ebff390c30383a6ac349647a73bf486c9deb7907bd2e4c865b4cff1a018c3836941b3f8497c44562fd9d9d4ffab089d41aafe538d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61a5706c1aaf89cf4ceea1da4231c153ee3328468c481019c3fdcf4efae99481db0669b76f3b86852ec8c70c0ac7a53c033966d4dce0f9e9719f97bce6497b80cacde79224dce027c6a31cbf171a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19aa8a7812f474f2cf759e807b593c645413b421f4fe31f76256452c110c47332d93f205b5a00076b37d1d69b1ef102d0494780f1a0888b1519b8978a45f632089e2a762197792842859e5e7a26bd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed313b833b6b87fda13f2baef25a7a6fa8290ed5e626b02166b4c59850a573c896bd4752054d9a31107b2d80c4bb936f00aa6ff602ef5a24ba320a180d50c49ed834a717cbd4c591fb574d68b774;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1667d444b76b953b2c4f6588a600a48a9361bb0746fb030e5de4cc325dbd99f8e1f539e501062a46900b60dfb28303b2e33c2a03a8191ba8341ae0442d689596fa1f0153ea068d9e4d9420ad060f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d30d394750f7023f1e1a5fce7abd8f05b9d0741453fbe38c69f775d308e2d32d37244235a66cc9a508e69ed2b05e9bce262e2dd6d384e453ffdfd9870c8d8a2bd9d02317dbba72b2f25c105f5048;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71aa1ab275f7bf6d7bfe19b366817ccfebd62f4d8b651311a6e1bd80117f8f757c662df10004516f1257afe00a5e67f0fd5fb1420b66331cc2bf37a28973dcfea4ff27c613885c78564cbc9599d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a05038abfd6a891cfd9932170e7fc3ea8d38e2adb2bd94ddea721f7054030bd49231b19e2763b4fb5d4874e25988f7890a2e9d47e522132d337cfee89d7f083c32ebd70f652d9940d0fd7843881;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea1a2992deb1e8aa97789b4abcf142bf4079b2f484d813415c43bbb899ecf3c56101ad82bb3692056fd51750c1b2c6360e0759a29e3c2bc36d7320235d193ba7ec67f26126238b7c555c9926ce6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8acd2fe908f76f797898810a08048183859a5f8d560b2ed5aa90f6bf50a48c3b1c1f4a84ec875d1637c0238d4051e0affc163de5b20f04d5a0fb3b374d88925f8395004e5171994e7cd6ea1487;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103d42647e13e8ae4c3efdaa9a7a69c817423d24298eebc8664784821958a94a183a295deeb02a930ea2f2ff3ee2c0dcfe530c3818f16a0c1aa4220c4bff79ac20e13ce40b980e09c8ef7e51a53c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98cfdd7f2fecf19499da41a54400d8cd25c1e8a63fd23a606617a5801cad7d4feffabb8d61dd64bd912ad33275417d9c29a5d17fb509be3751188c542ce2b5bca6526ab9fa98b078bb674e8f6f6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3bd54bc945de78d12e21fb914dd226bd45bcb77928ed38a47bf5371455b083e047a43a776de54ca6e62eb71a01c971b1359218b80f179cb2f168e43cf2c008d7cb0db7edb437c2b8cc78600b09a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4a28d931e755baa6e064822c60de7b1872345b20099aa34be6c2ce6f2f0e1c3bb7aa6edae993ce93dabb9ecafadaa920179487f7a10b4b3139ba017ad0eb2a9e2ab6bbd20c97f79c478bf65f8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b584d7a825c486df611e9d0cd750705d90698a4cba3139ddd2df7fe999fc43422a6b0e399d8484b883203e6ee68593d1d0e57a69dded5a584506d71324806a2d92c1efb4d95fac2a88795a5369fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e38c4d9073b8af75aecbc1eaf48cbd9cad90ddb64f9240a3f84a7b8b13d64579152f0e75cb69482b4bb8c0fc77ce257a858f2a2f144fdc3c99969e8e0173c9f289a50393258c225ee2c6008b01a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3759c2df9537929e4bafe3ef236856f67b2cc128991fcbcebacd7da1a23feece2692d668daa1ce2da714b0de6db2298f1a5854685976e89fb6861719cf21e9190283cdaa4f672718877b69af6b55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130e76e92e8b7b51a1514c7ed06c3d76b5c4ad430201450717a61d66fb4fa794e986f9bf27033b2f6db61f5b754a69e878675f34c62d9cf0aa0fe4115130b74f5a010364586cbc549a41e360d3644;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14310e975cbe6461135e8d8f0291dd354b2bdc7402b53912307fd2dd19fc6cfcecc7e504151abaa0365fa05a628e843ede01e6a817e313a4daa42d60ce6cc8964ede1ca05cd8b966c6305fde0bce3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d38e1210368e5a8e338cf10d48ead66348a611be6ba300d1c74c989ddff1e70766425ac502b05d60b962da7172b8cc96742baa8e36192142fc4b3a28ef43ae85e902d141c6e67fe21796f972b8e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f9f94d3d3b22070467eca13ba28ab2555db43c0e34dad776c20b354c97e8a66da9b6117f177be01585ec967ad9991f3015404ce45f3b15b618d5c6a02703abd41a046ff17a61fb4e73698144d35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13eabffe749fe3edaca6c7d9e2967e6000fa58be97b45cc50c5f61fd8bfe03a3ab37cf062efa0512869c925ffecc8f5dd23234377f44e14e53ed0f98f8f62648eda2c8abcc07e57dd7b71be930824;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b610091a357c7687a0b76cddaf2491c227c2b80ea652086e0b568992fcc04894a518cb59ae6e4a2f2c7af1ef5ee9d745e7bbde1b7dd6b50762c1893c7646aa2998ef2dbb82720a12bdee1a75f7a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5999817cad47e95a7985f0afc1050634c01453a7147763e3ef15472471a03239fa12c49604ceb480afc4ae71063920c5f06fd8a1b0686ffda7df0348a333eab4a0fa7f27ad80424ccf515b0fb004;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b0e352cab580a1e03dd469a08b33d1d8da3f803fae77cecefc2a3f59ab6ebba6a1bebaf6381245ad20ae9023fafb0611129b55b3b7aa1a7a0dbd33651e80a8dac4a467e1170bb63cecfb600b595;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd769d52b4d16b2beb3e6a47a859547fd79e43bac87ce136d74222270e13ae35f1e507b778d709f7d27d69e8ff2a35bd9b35047e1adce98fb864d6d8992830c1861f99b5e3c76c53265e4f84823ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11843de274ca4ed3114749f0bf9b46c46f24f9f11d84f23a8bf67f1682593692c1517192f43675c586a2aa650c3db1f03c58ba84c80e45c732b663095eb4202faed44314eec6d86aa41b903406dc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c9456f3750ba6c31128ec51bd6ed579bda85623be92860da64e852ba4e06df7d32251faece35b559c5db3a837aa854c898d342e07c5522949713d9d53d04169cd1de02e7c9743a623f4380defd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d251c0e852df932dc3d24582df021b5ebe9e1bbd1f1176d33fb40db000c0abbe669365a5580b473a92de721ce65c20820d8e97a036a06ac489d5e9b1d1b2b7c81b86fe9837a46fafe3a30a3be95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h528f3f967209d2e35e22782f3e0f22d3e2846c6233604845195d5a876c39c228355222e78cdcf33425a7d88bf4ff76874a79edc6e3cf635e82a8e826f478b648b45b230c3a4294f16bb5a1e28e7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f8ff6a50b436823af66bfd05a38961fd5f6035c060373f2d7d22206db731dc44664dd3cdf53b7e3ce366233c27fa2e399204e34421c1433f70dc5a66a7330802484eea7489d59e6655bbdc170d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee3c17d0591ca83a6065715fcf149c3eb96a44454533f5a391e58bdb9b3a0d9384d142f024a0e3312ab3a0612a71b4914fdbec19b8519e72e7a10a1774b30f6955f5b34f8067bd7a29a08f979a51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d61e8a769cece9c827d5564519d0285f43de3ab44d90de6a5bd9d80db43514859c419c1b9a27cea41668b25c49f672486fef5a55aad3762bf305da81c0256df793d389e755857399d7cbe2d222f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1085a84936f70b06eabec2cd6e8c45eeecac7aa763eb71548bdb90cceb48e8a634d80109fd9df4b8f37f7660c9df359ba7aaef3543db6b7dc3747d9678139ab917af7af7d14dcd42eef8a4f0793;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110fc4465c5c0e86d93bc96bf9f420951be110d5e4b14ad62406baa0007ca1cc56069cf8bc555605d48ab5c74793df33a22788a0a3d5363e955a2791d5ca2703e3ffb377a1ce62704a392d95cc85b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cd94d9ea5e79f6fbe0c3df0fa3f687018bfc9fb03969ff70ba0373dca9c540eb83f8f822e1d1dbf14abb5b4e951031968bb1cdadbc938dd8014f7f8d49e395645b09976934ab33fc271f8593d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bcd914a6bba0b2b5d5992b293e632524667408c2a74f8fdfee73c1b4d9184c1e6634c0453e9cb82f77a94e74c5e244293c0a591f9ff076f3345fa7a6166b932b58821387d246298b5718ffcc52bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53817f87d9ddcb8f7fe77c37ba590091c73ccb8486486bcadc6a6083676d269bd3601aef220f5b94ced5e030e58d96824713e145b8245b4ce2784712c4b39be7ceecda83c5f465e37cceb6e72563;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h406760109f9bec3f7326194b52fbf26cef870062b705e147e82c8d12a45919ac6fd5da1f8e4a1ffbdbc06bd3e24b3d4bc33ab65ef86f088cb9d5644ef09597a70c37ca1a481afecc4fb41d472184;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4ca4ff60d9d2cf595107cdb0aa9b026f246a02530420203e4b2a1203f69209a875d0037f82c5be923266dac901222a2014980826df4dbdcfc8fa4501b9497d4491f113b9d3fd5ea18e4403c2ee7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8e8b5f3fbb08d905c93a27410b390b34d76f33c79326594f95403a608dce652f57536da4006d22a55a27e3e25027a0f9a951f7d5e9a77b9999abd339086f1267937b4f9ab2af4a56a244e4b972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee622a01ada6601c7ad68c9fe2f72e0e362aacfa31d4d93a416843fb1cf43c7f5a584f566bde9998c0ad3c7ef8e432a05876440229ef00ef4c8ac415810b24006a8d4c493b333fd70cac634dfbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4377f140829af3e18ec8a275238486ab079b70ec45a0012708fc72cee0fd2792fbca66abffa53a7c3de39321ba781a7bc589e33236e08cc3c90c337aa249db7282cf4a0e3a0b8e926f26067de405;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2fdb492e029f95cd92ab960ec8e2aa058aac4b496a8bcb7b5db6b7bf7275099c86537e963ceb1d23ce0f4770a88e2f1adc80f1ec35af4d8516dbb9e2eacf432bbd0e2bdd38c942af44e1fe0e9528;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17174dd08288e83faefeb4336cebc30328c1c8f076133b0bc3390c8d6e8752f665b2b48929745aefc30017058214f479181aa3534d901a26db96b4733c15600007a9ab8921b84e79618e255ddb013;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5699f687b676ce1b6833e92ab52274cad33195ca1c2d8a233cc73d90e7b87c50ac6da0111301f947fb8ded89543446720b41ef6fb9753405304d4f44d693c572962e7c82277a6a418d415825d00c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42378a9eeaa2145122b33b9cb18b5cf41ae10892f3d6882adabd2cc06452d35aa551b718bb0e0e32a5e5d7708bf2b3ca715af68438b0f20ebf24f7fd823b0954984e29709d40c5435ed0bbbaa11f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha071ed16be759793d980fcf243a35d25c80a9b239e9e1ab4eb45e35e88280f8b2d86aa64e20addc53255500daff942f8eb99499fd47105337a5b49b1cd01615b983179ac258d345d7fe9995ab3f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d77cf78d8549b2ded5d98645f28960e94c3c27120c47542a9f03e5d5ce7011b825b08623644055fc6630292882b2b7282454f783c1ecfad29e5901b23a1438848d3f65c50e5b595a19e5d493179;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4474f8da91f903cf6c55f5fe83c0a3283fe2cd99b13ef8959160d5122510d666d521e77a82b7c8bb41a151a89b2bc52f005d35712baf804d6b997f01fa51b15df271e69e3c77651cff387bd7bc95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1585b6a80c4bb6c10e6fb1b85ee64c5a77dc7e10d1ab855cf7ac05a39d9191e87f52e25a30b6fbe04e91dddbdf430c7d9416950490270817368f3bde9630b6ba612c9f5adaf357aaa9e36b1f63232;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2889b0c4aac615d885f66e7867646b739ed270107d118424816bad54f461c6af38327528c0b033d85ea937c13ae9e3f8e4dbe7bf67b2126610b2748d05d6b66698c75543970e3359cbf33237322;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb2523af1b42b683fee15a86a335a296812ddde1d2754267c04214e60946c9f3e8d6f314d787a1a3ace389e1427c94e9a60d41111dfeee810f980bde350a28842cdc6f90dc5fb6f8496edcfa0112;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h151d1f7a416c2d4cca449ccb10a28f291a210b8c39d98bf061f41d1a92f984e4e912ecf9dc842df68f2c0e7314f232616898151e57a8f5142147b4ff4c5bc8f7b77e00e381e731fbb36a7a7ce6cad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161f62c33bb1b9b0c8f3c6539d3c1eae85a9ffcabba4783df03f714fdf2aabfd343dd9a394cd4c19e58537daa094f8f73957c6eb34b30f2ebdac42e815fefa9a2cc3439d67e718c1150ca9bc480d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e1a0e734910bcafbd195fef5a90db544bf3bf2fc314ea9b0f8c024eb7c2619fce25622d70aebc0058c3c5ad473bdb24fcff9565265c38da845eb99f2cf52e22238d150d475156bc936a7127ff25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1070c977a920913cb5b258b501d45fb438f2e96daf3ff3c8f7b90d141f1191591d50c34ea4f9393a5971a1b2c6e0e5837295316493badc21b3a1b073286f3dc7ee3bc09991e4ff449df88f50a91bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1192258a0344ae18e3aea6de3ad5dd45a12611eb42e823d7368f65fecf28353a46f9173d460d0053890d8f3d889c523cb2b5082cbd1a3bfa4ced3997dc7ba74e4246311bdf8678cd4fcb4601c50e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105c1bdcef7f57a67c663821a4a176f4de7efd9dcd0af25f190be125cf8b6b196fdc3001249721f0a8744cf14aca34590d45cfdb5c9a1b1f218475241dc23d00c4461ed5f8d78541ff023fecb66f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1098adf0a8daf4916798f36a804ec3976592adff6787f0317e919a84c6cc1d9a75b99c354c320e7aa8948ba708d0d5989a07d22af77b6fdc98b42960e52c8bbd6c59a710e9df6c6e308b00cf9af4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h748ccc00ccdb3a3f077ef862da21db0eb58c86a8e2c814721f9bfb497fe6c9bae242e3350d7afa24a00f4b2fc8cff62a9e9ca4d3556b3dd58477eb86439b85843ff6f8c3283f17a635a763728c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6deb868f4a30f04432f6a8f7d2a43a6e20152ef9807eff23ab0573c2ed54c01f5daabf9416b3a1de6cadad36ff70206b0de28b212403dea798392421720145ff401fb5eeeae83b8e0e1bbfa382d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d9649efde42b490571b1d635b6a59b9366a86650d93b27993c32661b87e1c2bad58f6295d439d0f815e52ad365a51c41bc76997dbe05dd7c4d1d980ed486524058b4d2b386c41368346e659427f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d36b39a571a673bcfd2fdd11bf78621da6664bfff89329fa4c61dce58a1c2ef1d6d4905533d79f7a9c8178abd8b91f186479bc70ceb04e5de2dcf4de8057e2f4d1f251b487d3dd5e65610a2e3c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1420f554eb808c1505918e5d0dcf8ecf240e2db03e3d2d0f697a6497e4a2d87e4517979ab9905a4bd06c227a66c16ec2a6efc56f9ebdff3da78f5cecbab6934ff4c76f8b1b320a4be008cdcb472;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122135e07e11741db9e01f3d3fbfed6bee925c8ddf85a75d5ea0dfa71b22bb9566222b1029ca20fcf706378a1512067a39a2a18b740d0ef6e2217976ad5a6a27c3da0a54bf17cb72fe56aaf084ae7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d485473d94b4e7ff5045e255ba6db156ef87656762414a03d65a7b8d2ef4b715d96cd99f8a8b590570f410e973b4fe3059bbf908097168940884387b2d00c81aa4ccf5a9c39601dc664c053675f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb44c565ca62e6bffa2e14f585a300241b88fafa9a4def6c383807efacc4a52295981ce9bf99ad85b5f51fe82599c5ae6785410d4a1fcff07e6158064b219d8bf7364a1af465e6816c4ba8ef53eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129a1deb172432402e39028d46d7079ed7682925cb6ff4b530012d992bca0f9ec249ee411bbc21aaa62abdf6884ed59c64423170a90251f7be4fabbc852a552008fedc98ffcff1aa025552c60a908;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0956f85b3a640141b94a7665644eb5f58e13cad17e9acc31a49478bfe6174e0e6f23c384d3fe4e399a7a2c311d6fac98785bf3cf201e2b89988573f5a880f37ae7c01e5e03436534b947a451dc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba44092745d22706ee50bfba4fc211d898fd403d3e87334c5e616bab1772245ff9b966e148040171b15df048b4556d6d52e65975cad1f345a2f82b0342b96d727bd005127162e1d0a316ea6e087a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d5c6cd0565086d8a458d873f78545a4e8b43362f510294c3ce530cee79579a0e1e2a232ad327ae2d534d746cf2d27dfa260c979b5ee2384dc6904f82c5e342718a8fd57c5948d19b46670d2989e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127e0938905d3e9908cfd90c9850cb25b501b2fb8a978f4e6505158d7ab1d461785ed35945d58a09b1b01c3b3d292c7631a6896b047086fcac503392bee19cef4c188165432851ae483bfc9a49f74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b7fb73f0089ae3b3a6f40b26a8bf073ca348c608722aadb3a05f8126c86c669b7efc6486adfd2e5fcdda344f8b137c6f4024effbaeb91b36c1979f12868c30869b419b1ab376447e982dfa0204d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4a3ae5fd1ab464ce60b12e11fd30871e429fea3698cf46d08bb7cd07f8291af1243d579d4e3865722bf4f54b8df7eb46ac43c1a62b6be1ac6cf62b9df21fd5ef6aad40078d5aab72a920a0ef588;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16dc6bd1b50bca226a95577a0ecd049ea864fbadb3bf27cf94f12a7d825391990855bdfb468f86aa102b044584ceafd92d79a09952aace014de8aee74abe4d54543101f65c25eb005e0699f80e00d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc0d402602744ff85cb27a6f6cb582d1e36e6a21f6c8f2476acc6688ef838dbd0628405107bc64c6117dd6b3db7c5592821c51bb4cfff4b3a5d50c48d1c167c4953b6163be6d3d4caece39c81320;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1cd19db8218a7c47e9431f22022a69351252149a46bf03bc3c878ee64f1f40f53295827090191a7e31fa6a4575b5b655fe282eeae4c006beddb86fe786d55e7d827183c99f1fb51fcdee66421b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e42434b3f2a4a9b947c706892127c8b99f2228fcc9a4806950baa78df08ce9809416f426bc07883d4f5caddb7cc87847125e7655f48ba07cc482a2ec8a5c84bb14557bbc2da0556e9e1eff5245d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179583b32762186abc928e41648dab3234c595447aeca4adccabfc2510415506ce15948c8bfe714eef6d0ca249a197a9159d8c3bc968fe761f1094ba13a50d5a8c35682e3635e337a282563a01058;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habf1b95e0ef2cdd465b8c6b579acaadd6a6d52a37e4c474ec7c2df0fab0c459e6a4b07707b0488bf4cb30773e03ab10aa2329d35375863c2522d0775111fd433ce4462b34169c93fa05351e83ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a55c75ae35514c0faf14e0fea861a505094301613c9207ed65aaa61f687d0f40625a6c1bf4868555b820ba8d10500668da1c5512fba6047314b1a2f99f7892031729c51d8e9132a49e9905fc86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4fc8b734f71d493d1ede18f108e8b406342bea8202fce461aeebf502343f89440c0f74bbfdecbe91f6b5ba0caa7228aa91a2d843ac506735cd854e87b08efc56a98a63d841b78022d336cef43c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3bb8f4e0ba8d9cc9f57f67f3f2a671691634a49fa0d7a23209734b535c32ec7f9ca2ad7bd1b7ffaa3f7f6925e53abb74e8660d8336f9e7ec19a811c1a823c39b4d18119994115362497e4bd2ae4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e11626cc502ecd03cbf34e99bc46caab543a9524aa7878e159717033eb2f504bef2100549bf9201ea07bf4fd5284bce7ad5731460bed65625026cb21cf7b2c16aea3af1d1d1af20896a2cf84fca2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f66fb21155f87fa79952699b3faf64cc4085e90fb8e2a9e5b638c54d96f4d3a7446711a73963be15b9d0c06429b1476f805f1392c6dc4edf8b52506837e84c3d53f0e249c94b697e69a52ea2dbb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d220dacdeafa88d433ff22beca1dc48a02df3757e358e45052f7658a3073f4edb57fae9d7b2437e2c7f58a1228b41dcb4f5039f89b167d49622334cd4886088755f785a2e44a34208f2adcbe290;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d794b5ce24206686b8f57a4c47dffa106691689bf1e40859fd184903289695ec28ce88900e3e4cda8f45f6b5fba4762088e8c09ec3db8f45bdd75a95c1d60277c1bfd9215554453132774456278d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1684a79b3d7196ec92a76b31c50499103dc6bd889b237987f1dbf1e3f7eab13f232a17f41d967c031e1e7acaf32fcf23beeb43d002ef59a06ebe3da03dfbe703e3fd839493dbba92d8046a326e350;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h618bc3820efa797c2968d5667d74e19f73919a3ee53912cb632e54390502840b6b1744137b2f1c0f24245971b46518fd49d00666c01ca418db62d49ca109326d77dd00df326c9589f8cd3e71c9d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72a0ccd721dfdd6d7d673b5a7ddcd62901f09bfb512a4ae000e7da83333c8ad58e25fd6d068a4085a8504af1fdf0827ff0bbd7c4bc381178a6200d97ba9994c87d2f31d60bd34074f88478ba3baa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd6f4fe9415528d32c2bbaf6bbed2b1d0c248dd7630bd2381ff7c79e8c614f7a8e51be41a34474508e8c70ed8ee5ef44835fea392950be2a6c43f35c22087bb580f50f2bd39ff05f070bcc64b0a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3dfbf62298b279d38125f8caeae20c3fe18d514ab18e277c46b4765d53a0ecd99bbe189f4876af86df0c99f58aeb4180b3b5d545cb4e993c5279366cb1545b1530abd52efd2ba4ee4c0db324961;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f08ccbf5ff1733f0851a476b002efac65c8169591a904c69439a9a0baf0a76fff28112613258278855840de89416654f7ef9a0dc1831e36504517db751841454271e432e41900dbbb64a166c1d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d8bec9a944f415f3931a7050c42ec0a9eee8e723468bd3e0cb8b4a1c453fe27896a47aab6131785f130a9de3fad8ab6301207f59ab4039a3d8a55a683fee9285b8d6337a5d738a7a592cb9a89aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b081b8302cdabecf5f13cbac0b7a4a8505f1b088272bd4fba402baece8d2592f6cce5124eb392432b6e909c75be9ee0f34e5e8a68ea1c88e5b8a7d7ae35685f6d05845615bc23133619e01b27873;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h263a39d55dc4f025bdfe908392e9ce6aa061d6d07bd25e6aaa7eb1c1a008838669f8ef5ce0e1a46cb1ac190ebdafbe7cc57d88bce0021ca646389f5ce077686a9633a422ec7a27d5f1d1d1bf4e1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e0b6ce074ad412ec7aa42fe5576d9b1db5d0a343e7494acddd4fdd0559b2382b337b554c308d6c673f4957d5e078f308fb3a811b40e76a9ef9c7bf6c0ea07054827d01d1330515e1772cbfd5b92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebd0a63d053d7d73e9f51b3dc5be878e827efcde664f7fd8894852d177cebb48f287d7975615995e17ebee73474ec71e0cf9e95847eafb97eb1943bf12020ff5f8677eb372506cdf9fb5bd2ac6e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8027326035a1a51f0c7f826c0e4c2af0ff8ae980a22ec0aa1b3d6ffedd484f00be985629b75efb37a3d6af574a4a39c2c56551e1bd55d2fb46818f233047a429c03e60600bc52a346b394fda8f42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5acf299f0a7535ee4a3a58c9018db2fcb66c8a2373dca3a3fc13749dd0756e256034145990dc452eb1542c97f092a974427e9c9d4867a95abd734891eeb61d23f5bd103626e6669b478cbb563821;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha56f3d0194311bbc73f21f48ef38806b3f123fbf3bbab1ff759feefc5ba17c77b052cce56c1ce0d918d801c7e326cc370b3ef31bdcb3b6040a8348a05325e0480dcea28ac037018ba3e2a257f179;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hadcca4ca70ddfa8c0ffc5740258c2c2f4155bc5a7bb59ad466391ca48cafca9c16a0a7b67f6d2ec24e95f26300fd56039e145d0074dafdefa08479d36359abc083903fb4b1851bfa25fd1221e8e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda743fba4f493bfd2cc6acb2d27fc04031352bdc970e71a49ac9cfc1446512d7caa342130016a1acd79f7a4f10a1a51e183aef4d485ec12df5c58c102409d98c6bc72dd71bbcbe257b2324bb8be5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1868e9cdf487108c640732b3b2ca6692cfaafb4528cb45ff26155093ca0472f645ee8c7d4cf1df795bcf5fe78d591fde8c8aea1a3d172307fab0e1b40f1a5d2a71c51f284403fc98dcddb5f7ae072;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19217116b8c7bca6344f70dae31761b0fd8f73df8b62f8c5b36a0e6834becffa8ef9a16b801cad3f14eb249f6863aa1718c1f1e54695336bfadf4f800dad8b476f264d0b2988abc0d7e870da49a4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ef54a44a2640f774d195003689207b86e271ee657ba1910efad983d944d8530a4fc9706f57b4dead86869ee8acfedd2217dbbd6a8bdfb6da5c0f475c2e82c61719df6e133224275bd340b2d28fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5eba2d7940edfa7971ab04895e8ce57725f86a4f89b850992a4ef24033e014fad5f9e7a8f0a74bc21f95475f6dc376d7a1aaf38f3135aae85f95c14ba96e3e908c5972cf4aa6aff6568ce18264c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff8ec6660c5169007f415893187018c6824fde78a852b094e2ae7a77d86ce9b0631e885d4ebae230f6a66ad05db96941fc143558e40158ad4081d9d056de51a40da3e94c4d0b59093dad51c732bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197122c599cad2701b1b5d70e9fbe55e2c105c65d9ef64077ed716ead80f65a7641590bdfcad9a01216287a2630c46f35d35666f67cbd652c02be70a213d130576f7304221d574cde8de111ae5f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d20ae8d0701fd7a4a99de0d222629a7b7afecd756d6125e69af04ba55138610249bbd617e3a15376e666ea6a407a66213fa9bea3b593288dcf9b510fb9bc9a4333ee88e4912fc95b19deeb0eba0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e75b3eb85aefa5d319d51889c099b662c75c4ee6e92f460fcb0451fe97a90e71538c2e6590e32188c7cbf66010e0d7b160565e10cfc99738cb0e375b221f2560b65c99753bea4a60724e90694ec1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce638d20d6007ba5b00ceadd17616045bf40da1cac82cd0ac035192a5d4ac0ef857213e3064568ffa3ece2f377c153b2a40ca5fb0441ac8b28d376d18da75e4d6db62d2bef46f5d5d4c8e4f336e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcec9b059cbb27c1e10f0eb9f89f32f31659f186a97f1817dc928f4b0daf1caa2c3fbd0e22df158bf212617ec048d96995b908bbfcd245e50260b10cb14ae8e7cba834d65e3da8b2512f44b2500a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e6433afc99f8a48bb1753ddfd22d11fcafdfbe2b80564e4cd00aa009d18ea3413cc65d870db653578c924bb5b11619fad7e92bf3ddf7522dd6858a4bb7507d4aa4715befce91522b9342b005ea6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150a11ea087938c0967d03a93b96dcd85d5f0e717fd6a29d23392b2a577f2bfd8b6b464591af7c2eb7fd8b0787d706942e47c8f7446874fbeaad5b42cc96482bc274c5bf8f4c76cdec010102e89d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109942d05cd4107bfe587fe6fefc9f33c959f717116524ce2e7c175f38044efc1508f4ab469502cb328056a191b1f4abe93ebb8923ded7aa294333a15bcebcc753a9a690f08e032a0708ebe2e3814;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c78f3f97eb18ff7a8fd252f7c9ea3304e4fe97217be7ea954332678b11746963eb77d83527079e7d9158dfd86d896e69300088fcf2519c41d725f40713cbe7110c6bf1ed445675a0f58c163a74a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4eb63c6e898ec98563937b64f6422e73572939da209d8c93ae5598a03aa06a47d8021d748faae5c88955927c1727c5495940ecdf8e74c6c55b902806db5b8555a97bd93b3688a53849a1cf852b77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176492c20e2cccac32c4fd946a77a979f42e3399a7c84028758024fc01c001995979006f239666a213dc4e29454af51dd4049abd078050961bb0339a209681006e0c7929a52c751187ed9d7b28046;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b29a85e5457ca2b8ffbdb1fd4ab6c8d543ffebfc88831f2257db2df7cfff7421f565f436b5d55185f119c99f2691d1450c3b2c3d0eb7c75817b88b27d2acaba3a480348c84729f55a77f725054c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba2707ec3afa19693ad0c8ef517ec54f607d013efc267a7513ce0497a3bb8d4d24798ada91927c90d0b085a6f672739690a8a64ff6e29ec37a36ddc7475476bdd8127e3d4aaf834aa1294c5a5977;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150568e500dbd4165aec7660c15b40404e242225d1b80b8b8eb190846a581d38e25f62b578714fdd89df7fdc3001d1f319eeb14b9da018b0fb20bb0a6cbe8d66b5d997821c15eb90dd019402fd097;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b838cfce54965da9aae4ccdb36414c3a016139ef4aa136c6ee93c6917dd138a6a91dd86bccee976f8b4b074d2085b25839b97375b2251a594007e8eb350e9e0e9ed76e7220d093af7cb377a583dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126707f0b2a327de2a5f401983d4bcbe21fc008cd5cabee19a41751306a79eb5d66354f46079b421bf26fa8dbad798522b094b1531a5aa4aea1f84ac820a6d1e611114030fbd126b0f9f515b433e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c66e8d1cb6760b73c0c75c2dc82c9c0ba7a729aa5abb9808c406eb2fbfade444e38a262a4b496a941772989f3e7c241c74d700151ed02f52a62bd9e3473c10c00c54fcba6113429782425751cd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199ff62ae14772805a6000f698ca4469e80cac8d64071cf9e5836ac6a376bc59dabb4fb167387c69cd9a34df0bf0b6ecefb0d0f316ef744f2f95415387d49e82549330defd00c1de8b3aebc4996a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h568e2b371c11bf54afad9b2229a4eb5c2f1d9cd03c96b86658449f40b47c709b29462095ad379c17924e332ed69632b4d74de5fca40f7557164cf0fbf00fdde8459dd60ad886cdb80af5d221d0c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2d7f3949d8a0629b87b0956143081d4d394f63eb3297418bdf9c22d80604296c7d1a63646b95bdaac0f9127fc05b8fdbbf4bf9f4dbee24fd0e01f0de3a024a8f4106f4acb199b2b152fc65bc40d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7598a80cfef44031285fc8c6bbf913253957e29ed00a6c90b9c3bfef76f620c0298392598aaee17b688f6b63f333b9b8b2e81fe18bf9ca4a5191bc8a042416c6d46e9f5594acde925a514b85b492;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16169cf2a0bc02d1d46b06efc56261c6c9ec602b73fc70e4e7201845cd6982ca6b0eedfaf7733440f4fb363e0da8c626379a1a4f14bcdf8bd4f34280238d13e66df97f0a640e156eebf38cc47b586;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131c625b10bf90ac5e902d4a03ca49d787d8e11cd8c8e0765d677a519eda8df2d1724ee5ed70fccabba450e23a4a9df3802e208712aaee685bf13ae874f030a13968615815e9fa0da781cee91a43f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ac22c2813d787a86e876ff0ffb4bd82c350fe0b6e7b620423cb502814c2c908754f159c65e0f731eb650511e3de64b8a394734efd70b2a3ae1f8de06c9941e0ab08af6d05968b023721c773678a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd0343d073baf20cd82f6c9d8ffc53173d664696d5dcc6fe2a8fcbe9c1929b66012062ccdfc08b655e0c3d49e1033da5f7446b0fc0e5ee78d5ad3379a4ef0262aa1d06a5702a2392a4cdfb7f4e7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11072010826724f328eec710d221fe34673174f1246657f8dc3adc55b40f28dd21f59c451d6aeeb08bf8077409731ad2f8cd204dd6fb6e537314585564a5f293f648a6fee798887a55530bf4fc5b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fce075982f0a39a0b056b1b5d6cc2157405cb128a92087d26d4b0797c858e49b392f79ed08cac56c814b3f592b7f93a624cf199ed48ec1f5d1c1311409e71627e6f1516dedad17b51e7c5a2f7702;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74dfdb7e70806c97bcbdbfa46d8230754e06d6608878002045c4da94fd804499b081394e720a0b9af904d2daca25b0c52fe7c63d27f172a48f25bc7562ee1d22e011896500adc81a3d205e15b336;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8d0807e99637e773e88e28d76cef6c59f36f4af8673bbb8debd384b9a023bdf79d571415b5c5b5de4052e37dab10e6312d35ec49bb687131bc713f6b807ff65a7033d3b7c88b5d7bbd8f92808eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1412352d0e073882d22d81805557c219c988eeff5b652b558934428fe08c4de62608520f8396f6db6c6c547526cd3975a99ed48a956150d47bb6d07f3f703916ccfe10787ac4a032d08c8b141cf11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194d30e2b15791b9227d00dfed3925821ee4b9fbde69aec6b660969feab12bc329dc17dd2221d2321ceeb1643c1087f329cc04a2f02114c4558a83c3f15d24759f0263f4d5bb5b27bc74d6b8a23f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d8ca6598d5eb6d304aeb3039cd9fa04c93d816628c9413082f500492977339e0004d24463a56a35b197dee12a3f215306477f5c6d8e71108f6b645cec22ced0c0c179a0dea77568d263ecc3be71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10df9b95056fc11afde17fde8e32896eccaf17f37ccc0434f31446f5eb4f182162344079514c78342685c85b0d51a3d9078cc74281e0478622a2e9741326b269882b0e917bb2eb4ef3a790e15f4b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15186a5bd8127683b1a4bf650a103268579ea5439011e1708adc58dc9474e5b65b5af6792913d3bf1a9c89df63622030ea4378f0e1c3a70822f4be0f15cb3143cfb17fc2017cc1b16df0dfed98ce1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157535fd4a5299ed8666ffb21db78690dfd286ba2ec02155b2d6b4d33103353335aed8342300b789cb5e6cf6c7b358ba0a82df8f4cdea572397932548f73a1ec803f4dcfa7efd0699efebbec3ea7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4e16c4c22b2be3eb1f78f36ad43f9c5870549a430070ab5a767e6c9b9aecc5f8807f7796c97e8edb9af80bf3ab6b3f18ed62315ffe23de013f8ca16ad633ca47bf46add6ed1558b5204b73d886d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac8d23aa79bedbce84a1a1f53cf7bc2fecf9a71e2caa54192e3a55b997cbb372d36dcddd7f5c5d513c559b25fdedafe10f38fecd2f63433c1652b7d48e2a28d8fdd173cf60fc84c062c3a2a22012;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a9c362dd7212a6dbe8f295d217a8d2dbd7374f2c5606b45b5a00aab0a9f024ba42e6f09f2d1cc899eaa8985ab56d1701e810f0d2cbf5106af65d4402d8ca79c0f1092fd0e9331e9722cb7929d16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11cf46d1254eb1a247e7d6004578383e0dcde8b66c29558ecf89cac94084f99299955089ea26044097ef2dff3f6602c2e03b5cf93ab749be82589527e839451c628eff12969fbadeb72ae1687d5f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca52b8e94137e8b15a32f98015ce5e44b4485f77e97e7cda9ec4ebdb8cb7df14ea496db20f20cd927d2a35113d11cebd42907f8f580861d7561638e0fc60dcfb0d76e739d05cbc68313ade64fd58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc06c11445ce5722d12033b1caf7399dba3d526aea9051dbcb56e05325788849d289419577cec713ddc151ecceb9247b9c486923d3c2445f486d7b3fa98fb02b8bb5a389ff31e0c004bc5bf77472d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2bf5dca1b7dc6749da642c176b6b835eae1eb9a84ce5b2aa4ed253a90d5d1acb53642d763a3f1e23346a926833e0d2c153b978f54daa5990141f66e7f95b340e726b73097e902b1d3a35016955f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103461595bfb02ff0f75e352efb1b6fe5c124208e26c52cbda470250ac7d8b7d81f63692fdeb0f0afdb10e1b0dc79223d6f6ef9984ebf15542412eab8d570ad85fa0166546eaa67015c2d1a7a2a5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126898e5b7a118de6d6d7f4f7a6ee7ac03a65490d89e5b05d585412a595d7050f3f4c6f7407bdb5198ae911049d9a55c44e77fbfb410bbe7f0bce2b75ce02c5009b0e955b3549bd06ff624a775f70;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ea39786ddf64a8ff54f253611094c3553ab45436731cb4e5f7e024aff718ed8501acb5db524705fe5a8fd59f31e74b82ae33a66eb2ce898bc5bc9e70d286f54f6febb0b15af83e6c06b2472fbfe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0356df273427dfef4d0b741b9f191cc2cb3744a4d1e7a63866c02c3b81f04de8a7158a7239e529bf55a69b400cad8f753f1050486c9ba07a13075047cc38f34b169103cba71111a51634ab78e28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182502118ca99a8e5168443abc7710353a87e24dbe95b23df00cb4379b6e7d176d3adf95f4a8843a2d50317c5fd3f53f35b6f8b4ecc55f87abf8e4b9a27a67d360b3fa09bec67638be3046befe98b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dae282b5aa1343f66bbbc4b0e4568142c52dc2f50f6314ec9c47430108974f3037f66d7a3dc91b59b60e6510708885e7a96a2fe871a366b42897802de1e2943c4d60407704aee4dcd9f34c9e191;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d6a74677d0186214ed44149da927ca37dd8e81e6f53c57bae4a1d35c843bc83aed8ce1da7f8c70206262d6ba6e9c4aa76217bf83adf4f2344b6ad664e4ee864f99f90e3b526a1170f994ebb8960;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3ae8fcf79b472c9936a84556fe839ee5919d70a138176a3482e1a224d7996e2df77a5ae7441a9dc4eec2296a88775ca1728c9b744e775786066858735efce5fc90c2e4edf18dd65be136c8685f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e8d16f5af0076cc31da6e861f36579eaea83103ca4c33631c97dd20c3aa442d59d979262fdac8114e49b04b0b3f9160aaddd02d890e4a41761622bae51ddb09b6986756e88f6094e662c01d00f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55a3b3ff4906bd9bd1bb8f54a4db7f9b7af43e08c711f48c48df34c63d8829529c5ec5c3dc75a5150ddf79593f1f70f212d959c41a7a880fd6055a442077ca6a06b5e36aecea312a54b2cda81c7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23a62668c0807e6b5c261986bb65c9215777cbe81788ddd52c373aaae5ee2797bd04096e3b10cd8e5684e1429f9afcc374a0d0bb5f381496fc9105e0f62276c54d73c1652259e726356a92b8d94a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3aafede76d0b572a7b2df7ca5ee04752bd3fbd6b91fbb121419b71d56ecf6ed7fd1292b1708339744ec314612e95072304e53259d8fe79bea70d490f64bc5dea457d7ae77809871b091b52124a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f957e973173f39d6a19e2081118ccaff1893bc0f5acd39a01f44051fa077ebe1b68db83e025651591231d2a82d9a4fef53b8dc931f14012c29435ebec51ae3f0df5a441a60d0dd646ed6688330c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb89f09c1cc77710229e13e6e66dedd09d1296292da79585cd8fa5f71fc1d4f36cb2603a59cb8cf79136a98f14fa92a88fe22eef3af534bc7bc459a65f9b8c08d2abedaea5e9e297da11d481c02a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd818879d3d854a688712154af10bb0f947af3c2e7188cb33ca71d8561694a802a986024d9a68d2a5b51fa0c662fa8aa2f0c9a64008e25e8c43ea94ae69e06e592a865a9aa4b0b3955ecabecb1c86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1921e63c6c70f430a6fefca7dee3eab02396d03ce8d94f9a7bd987e33ff4e8495bc5853079fed99467ad7dcbf8824aea8f84cd1385edd8d70efea298d87c2ac9315f445f9d962da4ef4734800a2ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0d3076621e03eddc9b42b6ebfd4c8b0f988ee490f401dd10cbe7f386de3a22946747aceb6be32cee905591c557f52cc638f4c9b0aa12ccbde370a98f3a5db2ac8ce02bdcacb41a0a801063d3d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd74cdcd89a53024736cd0eebb32649d39a7d40aa0eaf63d5d7c44e45ed25ac78880fecd9463d3d1324f1b1bb4b0d6d0987ffec50b2aa18f5e109aca905b5d3f42d9dc7760ad19c4f81d832fe7369;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f244ee0f9b6ca39dd8cb730694662558d51cea452654dfb9796fd84deba30d0b6812e72883fa38d703295770b97db7a63b746826eeefc2e3473513ae8031feb2c13f1a1e41932336f8c8582cac8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d67c676aca1de86e76b18acded8d1724e914e45f08fe008f42638a3cb891aab9aab24a6e48681b1def13437b44145fe6197f87c6f5f4f5f2966b861f2d9bb330a236dacc36d1bb4b98a007095c31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habece57eec037c3752c82b960c3e71ce15c411fd57da551759c539a040f90321c99dda028e162b4e8756e1b3355b2d4969a99d179080357c8f265290994088fb67bb66484a7c1fcbbaddc1dae8e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f48225134cb4315b2ea8723401cc48142c6cfbde271c4957732a8405b31d1263580ccf2fb9deb3d0e5c1ac4c2236966f28833103addd5d4a44ec903fd2510919063c0f376886f0afc8acac7939d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1554165c01c19ff1bb4659e3c12306f8bd070b0abdc3033ca36102ef80f4ef20a4a8c31d704b817d270744aedc6ec1853074cda0e46db85fba08a9cc441964906da0845bbfd7d50de564233941e47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99133bd6a3605991ff1166a628e47ed91ee074b877135633a570508ff3ca130816a8e7555fde627d763ed73c80bd53ae7c87d53be17031185847206670a6c146f1fc1d2c506671194b69cc309a98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12651a1bc5187b1f20361b3d2957a6e6fdc98a0f6532c944b54866190a6f2c5d8f151c96034102d44a23ff7b016dc875614c563abc97a9af9e587e2b169502b6bb1eae6fc9e5594913e071cce25d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb1b74aaa9956ce97afb9d390a913d55a9d360a54468231e1d893c7ae789c491125deefac9a0df2710474b7d2cb93a7b071990506306948a6d97d83f3774029683b13a0de18885fe5dfb8693f319;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0aba5aaa3a65d94612d52ee14467e016a03955f8f0ca3c7a75947f51dce8218021b75a9dc675afab9e1f7c566e6010130ead58d6c59cd6ce516c8c09c0e64346ec7e13314c71c23c2eb3fd26279;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98d52be4f5a0a8d5dba1eb08738ed31218e664d9919874e9e09d25affb442095a00f7facf5946bf7c7a67e8156aed5c5a4d477ba252075851911080990b36276187c0b468f785d04df971d0ff409;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac1eb90dcbc9aa9dd85e9d30177a5f17abd5265d471e17c447c786a606ae7e4e27812b44adc76baae1dc6ebff2c7adc8d439efa2f308b57dce52c3860b02ba1f2cc7a014a3ee630a386db92e40ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f0f0de27d7236d5cdeceb143dbf42419b606b1bf887046ed316273ba564d498ab3591d8a52f461ab6381948fa0d44d8d1f365cd9fa9c16fdb59bd926fc5ef5fa3aa3f3d45615764d6986ae24ade;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b3c8e56763acfa93bfd8c6af647c2096971b29941503eb9e7725c353e03cc3cae408c2c5b6ad0dd6194c688e47ec6baf05327f643a5b3e28f7483c518f177c471c2a471b7f68ec3bd796cdaf848;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192de4c5c9d624154a2bef07d7609d651413afdb9052b926bddc398fc44d83fd3aef26b88eb28e45ef9be9893e38941392888fbf16b3b94133c35e3521395c59ab364e228a1ce9c26c27cee05c209;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14aff7c85d9063e6adcda922f770da65495036104cca3f45b10d628a19fe9dfdf7d8f63b92abdf639dedaa918f0c770d2b24635caa82b54898af251499a2ea4263aca4581d3653aeb708c886ab8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf262ec26b0202ad4d3ea8d8ad75e6160b4d7d0e3a459902ecec1ab955f6ea3b42e854972ea09d13e94e44bfaf5e2b1c0e2e42ac7c62b927955e32ed25414c7843b6663b0c81c1fec8e9af15b7d31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h705a4c3fa3c383925466c59da3428d5e71cc36e75149fba2ffa79cbf05f7d263d465a6c5f803894070dca5fdd271abb719b92e9260d191fc22cf510797ea5a13c1704cad8b497c81940f1c6b84bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea007d1992686c97ac7a32ba761d595713eac2c610089a1fdcd3722a1c5570894a02caf958b3b92b9783d4a7692d5f3e323978fe228e695b8f3d9424868ec158cfa8dfa31e2137285fabc154143c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he05738693bc73251acb8a063772068358015d24f8c07577a28a7546b281cd0f93457057c767c287fc6a680edddd9778ab2cb74d31f5849da3dbb4697f9efe31e8bb3126ddaa2d58023b18196ab50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1395d5bb1c10824dc0912ce49d9f339b4fcf21f6628a14d47350f693895d240936cea2ee8022539026f2ee701510c698e48262556d837fa9d1fa4668a861b9e56d30df6672f19bee521db13dcb6b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119632cc66be6466e524aa63cdbeda22a8654db1eceaea8842e9f167075dc4d711a335d28531335deb3ace467ed261fdd983db8e95cc60bc86a4df216fe075b67e95bed7278ab9a84349b1aaecc78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154971b5c11d29a0bf6834f0d65d4cc645b8ae25d3debadaef50b15afe72365078be6e98ef58be558591382fee79f3b048b32d8126f69ee1e85df27572cbc7fea24fa84b1d1650a9965af0dc33964;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b89b241f7d9a9ac9e22d10ae58fe16e7158ef8759c3233b5ed1f1b21b0159c1b0977060ecca45a8f8d4ae17c0cf2ebaebf359bdf436d8d3fbd890194a33ce15fdb5849e161e8a9f45120b4d1dbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h811e63a0cc81151e4e84a715c80bb4dd15079cf5543309db4d03bf468c47d095b1dbc8ae87de4321bb22714a5f4a29871b96f5be4f7a72e1e25665ca2516834a56ba69afcd1225dd4f807526a810;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7a7d0aa09a8a0d8a87e727f187d3fd29473c05219d2855476feb129dce8d6468de74422621edfbc9d389b94b9476627c1351f6f20086c123d393459e329a793ba4262c735c31b0a080875f181ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc252db2bf0020137dd52dd4203bf9442d54134887bf93e0288c5f0b648a7ba2524677fc43c8be527220cfeaa8f2ce7069ca403dcca6f95c84863429be8ed55bbfc281825290992a8bc1226c6fc35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1722ab579fb837436662cce80c01b44d4e3138e13593dbf9e70d8c593b5993b46d2f46f525c6bde86eb85256eadec640b50ca3a1b4567a00db14c18d8cac04521eddaa9a771e19df06e6a3fcac91d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b40b47c958b1563194796582cff936d7b3514d8ac7e50b135e4fd44ad5ed04de009f66f2553fe60d62d04fa9a6a8c08e7ef861496c885f8089d8d6faf186dc92536aebd8963dfc59ad5af6db56b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90fbac66f9607c6f5a9e88fccc304ef8aaa3765d17546e3ff5b9c2be96d4971dfa64763afce51595c5984de49070297a2d9e97dc8f9ab30a76baa4ff74cf816e28e52d759b02eaa4a57393f2b030;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33d4036f4b6251b3cba8e7d886d9e30405dd10ea4d00f198f311c9add509614731ec218742a2d2d4b612855d53b0b0ee7ff379893e88aeda7f19b14be91ef86a2b3cdac5f66e6687206559ff6df2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c687894a9171941ccdd54eb3cc0c3baf868c2427a95e0421b568b5bc52ed3aa459b1b2e770ec0ab02b86844660a19c4508d5fdea09794e3fb2915a820cdd2e6011a5d2278b4d5427ec3e135eb252;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8eb86236c2d3c0719b34db915566b4bc339e621b3f424afe6086aa41bfcb2c72c933201d3b585c04fff365d7ee1967f27dd4f1dca94a5aa2c5f1fd626a0c896cbc3cd8de65f9ce73e1e0a5966d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b225b3eea0bbc747bf4f0951bdb5599f7eded4aac74bc1dc912680d2814e48e23c38f804f11ae50dc048b136353278736f6eae176fa8f3fc7168d158a4b6b95428398719588ae44e0587dfd2cea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7091328bcfdbdd5f687d154e97091eb76756a9602fe06a7c0d9a097d475729a6d8c0c92a2bcbd731ec07f4d83aab04b6ee52eb62e82731a5de8b9f283e52e9348dc5e0752715abf6b31472bee46d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41c84d661f2d9951c94f2917893986f9cb77ea27cad0622a2d694cfa714b72a664df728a5d994cc72522bb0681ff1accf82f0a81cd09edffc432e0cb0c1029a52db3b4b41659f7d32dd0d6a9d7c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7687f662a2e8cca3b13f410eeb8b7f99127fa393974f4edc81d5316fe76ea5ce735b2435c811b7e3d650bb4c245d10a164f61135a92f3bcde24dab5ecf41cce1cfc08bd89036bac146a36e7eb9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h638eaef91df63c93c7d780b512f077222be73a484e526ac141b406c05d02ad72b55f227a1afd0f6ee976f6afe93aae878998eda127797f0ef0c4805d42d1c4e676584162adf45830085c210dc7ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbee09e25b6a31a1a6022790f2b4a5382d82902411d2867618c622931162687b070d5f4f954ff4be0d7e1b09a7fbe1952f84c0d7ed36623cb7fb2d1137b73872a58ff2215bebb52182714086c373e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc20d7076bfc80d17b758ebd962cf5ad6f93ed56cd71613cece01116a8e13c4649ea17811134635af600bbe9ae0fa12e37d835cb7f34074b6e74518620f3d0429eff8636352147f2d0fd0e6ff7fc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a25db1c64111fc8b370a63264de60445b415fbf04597714a387006fce1175cae181526f92b1f6fe2a011665bf444098198539e0ce379c817ca36256d70714cbb6f6c0a070dbfd955855f87bc5889;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79b162df7ab512ed06f9320cb25633f5e793ff8da92feff5cd45ee839589d2a7f1bf54048ad0c1dd08a48569849d1e3a89fe395b5d333a1edc556ba1e07ef6df9075e1b9de58ed269b313bff880c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24adc8a47d121db84465e6a786d4d524fb299748d29445c8d3ed3a8a1c0cf1cab92358ee5225768c65b87796c105ef1afaca50db4101cd2a07889067ab0260755557d365de081598053b482a6f39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171a6c86614c897f7d5791467224e466bd272f1511fd3ad07df24fb79b0f8067e1722311fee0713f87bfd831c6a5b55dc733504e0d72ab9d6ad468cef7ac4fe9d9b1830db7f1ec41e811ea183570d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h377604859cef5c2e8a0e8230049c0c4d47f81f304070e30891299f74e61d2e3ea7384f1ee4381e840071465dc87bc9c0e478d48278318148338f0630c5bef98a3fe4704be29a195588235e05e4ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6252a818ccd9f828795bed7d233e299932f0eec3050faed0d65fb380d7bacc3cfb925f271a798660838f74de8701f003cce02da2c34ec7ec97903e86f20e0501a7738ea6cbbbb511ba7a8f8427e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fdd9daa85ef0f4f35672a5da4d3eb0c2511a068f28f47cd444114aefb436dfa21dd96508e81369519e8f215cfa58bd142bf7176491897f5f07c8b8324e0542fcce1e075ae8498481b93afa28db7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d2c4bd3e66cf27fbb3fa8d3d6dfc1d08edbff7fa8dc6ceeef3467faf8a7860ba45a09cd35ddd650530a5d258e1df888840ea0ceb82fbf36d8fc6c6b9cec6f735495a5c08aff097f79e78436e01d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f037a29330e1cb8b1558e121bbbd67120302030203bb085e05961b125bbeb7d9500f2fbf77cc24884a60d76e385fc7a7505663e7a16f8966e85f9d91f0f0f8d1e3a78d5d9040ed66ab8b41772d33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c70f88599694390ac4326bef9bf2cc8eca49b1b9354fc23385806c29eac4ad07ec3913ea5f9f6fc0ae2800c46b86b11c8eaa0eec1f5b70b20d1ade99f6bc0f8f9567380e47527fbd787e688280f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9260ac785e83c67dcab1711676536ec441fa090b7ce0cdf410f295b7ae5a9456e8088bc06f4ea083a4785345e698101ceff14ec4550ba56256e40875a594206c7096a9bc5ad0ddbff216dd8c92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd343e2152e6c45c561aff4042bb0f9670e09096399c6c19e2b33483b4a2eb05f4a8e34f9fe64f401b9e4d61486211ecf1b90feb182923006b8a9828ec1e8579e4b658bc0c86b2974e621199182ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had3e641c1a10e6fe5104ca1df0241ddc0544e4dcb8b10d371e3e325a82e6ff23be1a01300a3acb24fa00be3d0cbf3fb7e74e402efd84363872df03af538f09725d12f0410fb0718817199eb3035f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9f6b4c9336e5908a3a192859a1b80ec369129ee2bda4a003487d545f6122c6cde4b6dc310addd2afb1d92f79b80a46e61bb237f17bf07ae1269293422ddcd238773f1186c3ab2074107d7e52bd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8153241ce52ac9b0c52a4b73066d76852f588eb73130f69d48c2b51bc779196f6d9e4882538c38c2f04df12807f4abd632940805619c5fe0259190af46de55db6e2e4dad8c8f104c51c8929e11d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha37b08c130ac234b2d32ad38c32e9832489f28b483878972bb7d989ebfc6ff6b8d9358ada6d0fc353ce1a1462c2aaef73954f55965fad4b4172adf981846d3fcbbc6965113da4f492663946376ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138db5ace48e7edfcdca45cfcdc4f2ab30e41f7e63d53fd7fa7514d5d5a4fa931b275fe46820a3467fc11d60d1a417005ebc0fd5f24d1b11e752d8cd67d0b98d33bbfdebab234a3748793c6b55b33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96d8c1fe59a89670d1826dd23a29d250d3f12a6dc5096d44e45c809211118c99ab91dd45d516d2c7a87f5e2c9828767be8bd532bcc657046c92f80c12ecfa32d0553abf882a242d5ac2890105f96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9eb5a55406cd379ea432aeab8e416620b3c84429fa3cd01f6c5a3f52d52cb7d927480f3ebe6f34f55956fb6adebe4c3389b91032d7fe21a4a80840540d4a2aaa9487713e802cd31b39f9aec8767f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e7bf8e9d8173426340b5dc561d28b1a415d5d3ec0a4d56bde1e47da2203e41e9d1bc2ccb04e0c1dda514d17d39d54716ece621c327bc84c513cf73428c665f401e2f08f33b1b20f5fdc8a499b4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166c7e70e0b83ef04793039414e9ee22ee2d7745cdc3eaf6ac29a111645e23b9f06a958e72a34521256456f864b0707ef1d6165ce66fd85e67246b969a5c70e68cb7d40e9e8b06a1a0cba46de7ff8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1205a67abc2dfa6172aa5773adf3de7c73dc195c02f344b5d096f8302f0c88874f5728787accf2a8ce18fb369cb675f6436907232cc5abdd70c1633a0317fa8627833a917e153096285b1df716ac2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb3a898387285817f8d2624c684b83afd7ee5e4898cc2553acbbee4599bbaf579ae7c2ceb8654f5bbad5e2700f55a7e4a8077f0b524641b4ab252e58e3fc7a7134b38dea712e886cf3e439b58f73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b9ef9194d61beb0b3e8c55f8618fda0b9d1b0fffd2d869de974965068d8613857bb0c7c594b771cd2d9c8a6fd6d5bbe967308819542f8ffc0cd2f245cf07abecfb0b23c913c9a6499632af46ea6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1410686a1c4ae2bdfa50d8714de6655fccd7855d28bad44807aa91ce5688017b6598cdec12b9d7ce65b592a745d7677606dd4073adc1496768ed3d6cf83d1357c490f33963e0cb566655d288e267e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5be3c0a60489e6034ae8c762002cd00e3c37548c1cc961ec65b1a78d2e7fc8a8d756a3f1240bd3e13f3f16c70a9a291b29c7e54603670baab0d7642980ebd5aea04d62a4b4e9283c16b1eeb4616f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1579344e455ba6a0114bb1c895e7bf7bec84cc83beabb80b55a8ce197225c8039afa3e89d223c34bd882627bda24ccb36a65832295d5999523162ee160ad1f211d4965f0e584b12c9db9acd599ed7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc62507fa7d53e3b8a2ed4cd203e8b574052e7de4a262caa427a8d2277fa5754be90db9c48f9a324afb698f6cad7f34ce5fdb29cc8807cb85ce3fe81166fa2c5aef25fcd5bee6d90027ef3d042a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h535bb02995d4a4fb7c63d0939715e88404ff431615d0df2cc563c7317518351769c77f48daa75e8d604cf54ec7d95a576e33c4711230ad4796d366da51734b622d99c555200fcd66f7bda48b82bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a732ab8f6d3d64c12f106d7396ce9ac1c54d9e1f8d4ee2a9e48fa5bb3373c70c6d26850f5be06a98e8ff86d35c93ff568df94f5cdf811e488c7ca8c05ddcf74004c00df716ad91d5681ade57cb59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa0c4a819f98607a55e47dd29f3a541ef462efbd8bb138af0139dce59720a3e502735eca4993a2c439b2eecb39017682c520d4764a50ee4ee9998c4ac20b5cf14911f6a9155da90dde2e7258d1d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15df0522f4379a5ce8df004cf59a9ea22ccb889e94ae0031989ff3b0098372627df1edf3d599ddbfa34b595f8110b6b43e41eac417dd3415d948c130804333160fefb8798d1ed10a8df8ffb9debe5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had7ab3a7d818a95205e0f20bbfe9f7b5904b86a1412788a1124a2ffdc6bf1535af59673f9f1a9858093e13c757fb36eaf359f3e64321ba765cc2b531601edd63a1d35b339f7ad31507d5d4467a0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172b51d4ec004a3c21c0817b28c0b29c4bd1621c6982191d7e3a2dc62f19b8bbb73edee66d469d7553e36e8a4d351ed3a358c0c644a329907a6621e619dfbad6a0cdaeeaa644f112fa9922d6c1ad5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196b339bafa8558bcbe08690df4c24af66c02fd533a64397c1ba37f7530aa2141fceec46b1b08d917e72f641b60db0361056724f6d206221acdbd756973a57b9a744d23472a8cfd3cda0b52d9fa2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2aa259d1ee8e7d00be73152a76ba7430b916d33e542f9c2177b663277589a46c503899ebe458b05a817b45eec759486da98a74bd2cebc9075b3f1a67012093fddd9b5c50f224415b295cafb14f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdee5adad89577ece667180f6d14a18a70f5805c11467c1ee924dc71e67be131aae6d546aaf8236caaa2b983f144589e042aa68e646a69076c7a929b306442a16bf63086576e3af3e0d9fdde160a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8db5f11a7e866541d5732eae738695b56dcf07c766135d3ac460696240dd6cb4a1141a3ced90edc64ed534592996bf4e4a3caf6ec2abb19ff21b4327b29e19e86c68610a8c49235d500ab8fb531b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76addf8ccb87b460ca3ca35a0795c3d6b09e81a96e4601132360fcb68e2e1ad4586c97f47df9df39e3257519f4c091dfb5777139cc6e750ee03ed9da1fdc28305ac9ef0934bebee7b81838419109;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2eff6498634ee8d6e6317c8f0bf33d91039761a9d30fa04a99c96f7e13b95ece5aa55b2a297f1f35a08c6c5d57a943a14ea3b0051d43b3bb36242944469238ce8155e257038157c18c806b61e037;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4af41f3dc8aa92f8aa827b57b2f387b1b5d057c52945067fb04d4afe0cc84d6e7744a0978d7e4031626c138ccbdb98db55f1376b9f2b48e0fb8468ffdb5208aa246b6443cfbad53db702e7bb75c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaba0cda85ff257847d4a620b921780f4ca837c9a4c688878980f25ed038f2f786447c80e8d8f157f5f12959b321a901d7a8f62e1c456e59220c6e7771fe071153bb379487a307191d0f229cfcb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d8c0ad5ce2fdef6763f35c60103590915c3532303fc0fc1b793e2d9c9196a2042ee3fa2bcbb9b90dbaa41fe2590be8eff50a1538cfef97e5c92367ef171febd7f9fce6e6bb8aefc12028feee34b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fdef67d8c4d742059d076c93e723aa56f96d8a4671ccb1a9c501cfcf24c03a1484aa790e58626ca087a5c794076d2a804f6812626aa98348a923f00ab887945576a46a1399b909f61edae45285eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f0a46182b6cd69537d62b27fd163a947f513655195ea9e8cfe8e79cdd61a65bdbfdcda8ed91ba91c617fe19d5173433bcea365e65fa85152836a317256d43316d16af0f3fe1e5358ab86c5ddad6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4077c0b37dee1e6bf2d0e610138d2bfab81a2af874bf803e084f0cbcdce886af5652213a2f598e793b786a4c87f9addcc3615b9a1eb8ffa899d58716c7c5fa5128094cf1688cc3c8aeb344d85ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14850b8257423d678f2ec9b36cba0e815a3fe2e5eefc09560de6b673fc4105652cfe3ed955e2454ad816e927c0b38309c77b4ef8d91182ab438b31011ee59a582418d4da9d2e62eded5bec292988e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haedda8ff56b41474a2728f23404cf8c739dd8abc27a6ed03fd6df1bb9a142e5128fea85bccb3cdba391b82d6f29a89ec2ce6926ccd67d4d9b807317aeb04c9ebaf57ecae727ec185a23b1122ea5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd398b11a6190e197d7a1d9eec6935b0cccf9891965bb32b5a795f441d5dfd609b66c2763cedfd41fcdc63b49d9c646fcd67fe42ec1c9a7efca4dd486fe73177abd3bd49c29e6020a31beca9d29a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137fa27d244cc83894f9efa8956a083d57cc44e19a723584ca85435335bab36b33c48cf9e298cd9c5bcf63ccbb0283304ea60e895f9e2bf965b9f828370ae1be06df981215f90f0226d6552197a25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd19bb5610b00a006273d81f0cd785df3fd4e31697a8fe05159c7ad22f1285bb2b3094fecf05ac034497f34bdee860c6905f527cff31de461a009551340d29de0b9e087f54200ac12d9f7ea617099;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197df9a016ffad96619e5a7131907227de69ac1dac689b5a84620305a3d03cd95bfd447f7860090e92e0b3a93758474b14183dd5d9b751e9b08b8f186c2eb20ed9dadc6d4b0a08f5546213cd7b226;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e714a5a0010201806a4c3ea72d2d8f0b08b4c61a57b3fed512d0d66fa78f080b3273db6c3a01cd63c1d58ae669b1ca4f75786a05d21413c806f96a9aca645e72b8cbdf675f4d4433f42ce24577df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf322c2e04ca163029d7b27444d605f988de7d8bc8011d5c1edaa44641695f3eed968728d0d9299bd8d3b8b5ae7214d06871b6b0a3edb5c69d8ee1a23d3903a106bc561caba830f252b3021c9a61b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd3a4f3bbea84a06d2e2bc5e92cf48faccabbdb52f346c16cc70bfa7e24b3ced443e2ee79eaf053afea7f1f6b957c35ab5f835943cb2ff45cd4042095ae3b0dad8554e187d028cbb256d51c95f9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2e78944f34056417665b8c41d193e2498143cef045b6bc90cd083bb5a380216b9ec26e2a173026429225d2920ca239d53c41823aaf4c866d73dcdca5c998861da3fd099194e4b879d46ec85247;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6e6e65b16b8b9a3ad0645b0dcae38893d634a96c33e996db048a1a43aad1f3205d5a8b9322355d2913bd3355b5ba77c232a3ae44a7100fb3b6f4088d7f010ffedaad1c22e5b38d3d170c745bd6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b92597033a32b6d490e8a4b6c5fe0ad4747106cdc6895f01b3b37b3cda61057e63b77d662fcfeb1d7a28cd8e0e17e4e6b192d2bca1e7bc558203a10f663452df0d9bf7f44779df111912297f6d29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6de861acb164e241f05456ca66bd10acefff9a77a7b124fe7f10ffaa9f41d4d3900005072837961c4f2ef7e1098daa725fe0506d4b1858292574af2357c17c345862a4c9de154e7b37edb23ba52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1285a9e85adb78972fe4a27b6a587d570ca7a34ed1073c038e2e14da29754a0552c958a156dbee6706d9f3021b99d9cabfc61df0416da905958e8345f9ceaec2dca8b486188044ecf95875657106c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e7b38a751864d3c6ab16f8cb7f3457d552635d998ba572ca5da00448c0b364458efb0a683a78eb11c8af2785b76f15cd929c4858d7d13b359d51af6084aa56bc05e254f1103fce2d6a008144b2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0093710701af44bd9108a6c92a330d19a60fcdd1f170fb2314a3fb8ea0cc12865659f352ef6ac99b63c1436ada19673012e5a7e816d8726aa9151088b76afda40c602f73c76b69a9b54724576f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ebb9e73d4defeb29a2f021c87f1c3926d0b1ddf9aba845d2f239e67620c11d59a9a3367f06ab96ae5d8da934ab247e53ac10a9f45523cb5d26971b1a160fb144719cc8850b4756d73b5f58ebc2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fa8eb5c368dfca4d3ba09d5999c85dacdc450b8eb6f70bc52d40ea2ccb4f78367d8162fb21097be4bb72ae921f7ac78e424dbdae1887920a9cbafa4c4af6a41be645df83d7455bb8ba40631e99e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169768f9fe742dd81f27a22decd029447c1eb80582f3d7325e662a8c0a17dcf7854c9121246fceae2717d3322d51e5cf569c3e0ec111614ea4d9550029650e9d3520972470b4c2f110e02f8a2d16b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h73addb389853dc681145e8346a9169cd7e1663db02417291b6ba08ce091f4767ff14ecc1bb572e418085c14477217593596284dee3da6f2b5a6744a1f10e5e2753886b5faf11ae68e1fc07135155;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173178b3720a249a36ef4087386906410cc5fe423e8cda890a38dbf12b67e7a758b67b3f1bee8bc5c876471fdd35ada84d60da49c9620e98670f0090bba311c930b3100719f1075ca6345b53006e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49cf222fa43d2b2b7892105aa86c258a01b7892b0d4a7a0f65a86bfd24d763463e715a1832483c4422640b0bc9b102b670ca3fef547cf1f75a259de93b3d6121e4511ac3ff5dc6aecefb5a68997c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e866180fb3e6344d76088d98433963b57f90c02426ef7da9677061cbfb2cb8932aea9e375fd5f9c3cfc7783cc54b0cb93e211f21fdfa274f51c706cc2a4b126edba3f39a7e84cbf640b800a9ad5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189bafb23cd675354bef93153ca729c9839f67959d62e685a6c722adb8211b45e7a69d573122dca0eb210dec116ed092b2d880c0189d4e8fda73f206f66900aa8cb05dee395146ce8eda2def4e414;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118d54ac61be9364f895281d87baa4b97e13d5a9640177fdc5d68a79885ad808403a485392a84943002f17e776b8e70401bf9fdaa7e5bf82fe1241a367b7f195bf4462ed85cc1ce3e61474410112d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e490ee99418fcbfc49b621d4b3e97d25bc21058827b5a7263ad908af571333311f9262ff5767586a587631c42353a2912c003b1fafed9e9305ad94e2d887089e18b987255be0a33df3ade39ec0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5b387335d353aff3119dd49dd98c57626fc655ac95230489734b6c90615ef42eb18a07c40c83fbc4ace24a7139773bd469b5cacf07ad544cfe89e3d9196b58f8748e28017a630e9f2acfc71c671;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e5435020dbfaaa4035b25ebb9c447188599253921be3ee34f2337f14007decb5c6d81c1661710dc2b4ca78e7f4ea81fce966aa3ebb1e78ba62e5b65ee4291babdba123cb4fe81623cdac8f9808e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157f59b81a5a915d2426f2fb31a0bb450356b75c1a34ca239e4dbcd6d36219152747bd0cd33ec45887ca7b56c32319fa5e6d6b42c4cf21f8f0c722eb131111236ec29f0b60f93cb046e885bd8282c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffbf0f6d175c39d7e7b2d2ec0b2c59584870a2e4a8f4cc660eb0d3aee415077503d94c6fa1f9970ff7880828382059e2566329c9800df385c11aabb54ef5cd6fc8b6a1264c16e354c360b013d35d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacb32d86d820322350c168c15b9a840799550c635db1ba04832cac936bf150afe4c986bd1e3e721216e2c99a04d0f253f3fff956871c1ef18b93adf2f980e406ccc56a53dfd4178af0b582d95119;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35ef2faafe06a9b2de8c0849832732a8ff7815dac1302f0313ad50d1abbe3d93702db91dc0e05e1d8d99e09a3ee1308fbc634c0893a4d3aa4dba0e7b853aeb69f41f9a1028ec7ea732b3d3a0dba5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1669832ab34f1aa9f5407aad6f09fa0440ca08a083f7cb0eee919ecbb590fc98abee0fea77985f0fc4ff6e180553d396e2200e9b531a42f8ca5661dc2e3d6f2a37731d137c01cb43634dba61914b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3337e4a9a221cc458d6cd955824ddc33083b8ccb547043666863ed408d718cfb42188be24643ce8b3e5fc7ee99f3daa3e88b01dc90e802375efe5c291b4e4d4b3296e1224f71a3a443e21b65913b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h547c578f717acfc16d4f37a18d76aaab8501b8af919e61e5a89b1c883a17da74d93b6e7f08add7cfa2c7e0817f57bab7e8574769c367f04c7eefecf71ed74d6bd1d0926bc19736a43df3bae74f06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45fcb3c5c219160cf6fc194d61560d1a72254e0e7e9e275c4bfcd5952c47497508082b85167d97d754d6279613afdc1f09c2d15e15f4e27e2c2acb33064ba6226e15db36b085219b74b1736babb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f626c9b48c74afb217b6774138c1adb68f100368cf5b01aa3dd4059cca11e422cc571962062df30ee452b2556b1a65507d4b65b28ae6df7b9363cf644462025e0d60d14244360a8dc379e95191a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0adf85a671d5b87023ba4e6cfc6804d15d6c7e7575a5475d3a74b6f5cabc0a2861ae31647f8d5a9463d1dd4c5fad26677ba8902d6c256c4e7937577902a1a5c5222b690b81303130dc3d210d910;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1825f960f64131989de43e42f31a0955a111a3fb030127630af8c6a9c0bcafb8a3e2bca21ef3f7f5e11acbb5db215b9ecbbe4298569e53d8248f8cabfe5919f8bd7bad5592380666c4850a3e08bd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bc7016b86d167edb854d8beb1161df0cf7cff58aadb9fdfa7f35003f22537a96dff5c6a08e435d0cf50377fb8579ece60708a3a38e7ba352f09d4f4022360b5bcf57126d0da4909cfe8ca83c5bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38c51d68d9c35f430f1cbc7763102ed943162ae65cbb8ecaa7c685b59ed161f6a48630242fac62341660a71a502b00b3e4d160ea9cd4744335c0ae56e1cbab0880e8d8c57392ae0320aea8a1be44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24e23f9d471221a98ab88a4226b2ee1c690d32b2c5275e88b8b8204e90366c10df00bcfcbf1eb5fa024ab287b3b5676de8dfa0e4bfa00bdf435d56806c71ac5915dbc83cbeb67bf47e8939f87897;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e3269c69f8ff4a78d33f6c363bec23981356b62a000634a9ded27433304ddd31c5e7040f1a5f59570d7c471db1c6e392d266e418bf7aee443d61e0e8120a212b9f186e7171b8ce9bbcddc95c0ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h595ad3a0f22b656b092376bdd13b83ebf1f1524c12122e9952bcfccc940736d9bae6499d2d2d5f21e21ddfce9f3d1af3b1acbb94756967621b88779a74e5161c74b0d4a215dafbaf06827c4d7c8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c2ccf9a4f900ae1ba52694e12a86b831a42cbce60884ddd07dfb268e4e4965bf11a0de1ed9c04a834142a9ded9383ff839dc10c3782b7db918173cb31cedbed38dfc591f51ba5be33630ef70efc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hceb064797dc54aa797e6b92695d29bbf350e28f821278ea88c9ee2b50dbb04fad9c336ef6fb1d407cc384ed7a57aaf0555ffcc5e209bfcf673cb4de7b5924145918e27827b1ea8a4738d18441871;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161c8db7868f76a0477c5ff11076d873e77c17503280da3328860f11931a1551e760f69837e34587fe8f0c5c9632d481c59241b20a039260b0d8311a8c970343b5d46fbb75ef180e700440123c04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb828ab56f8005b5c7d5e6da2c22661e3be338a82e05c187f94625cf8e7ce4a9504d46d665dec84dfe8082e52bd0c315074c2ba94cdd94688729344089cf750980466bad7f0d2126ca69b566e459e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45634985e9f3f8ae1a40a2d93b33783e0eeafc90d81ecd61007b111ace9b2dc5d936a560109219906a02ecea5c9eb87ccd404fa9efb282d5570d991cc420fab1bb6854c0e9fdd95e9d9bc7251836;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b5a65d9e47a53da6c6f6e830e84bc95f431371571cf03f04b20c7b7606ec5085373391475c6189c17821dac237c28c683dd7d03cafe8dc92015714b1ea485212cdd94d6d99e6e511d03b66b7d4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe995c6e371e93c2806a932850f1aadfe971f5533e8cfb654a7a1f4e7f2a6e6b4d73414f4cc1111f7d007a8a9448875590cc1c644e44f29eac865d3ad325ac88190199f26e693b246e1891115471;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154911ee01a934151e28cc077a27bce1af02844e986f9d15d6b6fa98f39e7f2bca48c808c44e6854ab726f9dc030136d46180fc3127588db73c7632844d95c9648179374e0d651d745537eed029d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15614d01c74cdcdddfdba4b50c135912904ead818095a24c35d0c23b32d5cfd6e90be0afcbd06c32602d1911650a81782f24dd42406c03e4623e66c17543ce639797528b69621a267bb9459d2b2a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31c20c7e0f374cc74884e8a00f4e4922d153de19c4fd337986d49c3bbe027277d5523e9d502513b4fdab5aac2fe29287ab41f78eae5c19687125c20e2d68aac96724082f323c6cc22d15e55a0f30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf2e8ac22481f7896da73e4d0a7d519b3f6ad588fc8d415662ddaf8795ddc26c88a98f218835df59fe09bced1d271acbdd21c57fa26c03bfcd189552aec6a47c89da83b83bd8e9d50190cc68e4b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12db3ac0f3caac7fb3739e7007c3396cec1431e434b74566cd2ccf6512ecfe801ea821db7b9eb829d8097f21205a3b2282d0888392a8a993da19689348fb603343d8fe25cf08cde8c3d5bddecadcf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18495129ebdba28ecc1045e8acadac64a25d315f750ea7af0f018b0cf53b6df6f7dfd0c9fefd71bbeba6efa8580b3a67445d28234c3c93acad89a72b088bb218894e706f0addab37ef756865f52ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddb1c882d303e87979c0fba60a7dcfaa288fa585a31d20ccd76fe8927ca53b5e90b8e413d47d7b18124eec667f704bc1301cb7404591bb2f39996c7df65aff063f0a9396db416f099de70540714f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1098c7132ccde4c8a874c2d4e75e8b4218a22bbf25521487e4470a98caf4f683d75948b2e82a996890f97f5bd9409aca20bf9472bc9c8576797a787212b63b5244952997f60f4f77d5ed672fbdc3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17826653622b5814423cd85763c1afd9f36a987a10b50911b2c15a0eace14031dbafe708a3ac443e77d064cc95881871dce8be4e5c1408f91e2520929f08dceae987e8d4ffdce73d5da34d216c7a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f33a3ea647b8754d74ba14d3742c0b89c00ff865982b44947a0b3dad9e990b9c75ae56df750bef70a931f303cc5ef565c0f4c994664b3a8ede302f21189083065e8ea21a98ce002e0028967cad2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d89566a5410aa0ca3484839d60cdeed16684158c5578c9daaf4d2edec6ed4ad986ea5832e3772ce6042bf68d99ea1554a725f54a684aa8353d0695c749494908e04b1924c4ad9f31b9c80ea6df1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1998e94305ac9df438c307a968d9b4e7431530c96592b48f6e930ab6c9ec7e0c8117526b94104884333291d655dee1ead4cf3500cc3ede4bd868ebc67bdf70c8de0d4e0777de8bf99af3cd8500862;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1433a5bc2d35aa60297803f87646aabae6148406700cc2e1b838e6ca681c13f213ac06efce702581e5e915d581a01cf0a3ff257adb45526fa1aecb52c893ca919475a12b5fcc4002d36bccb3e8e51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9e2da6acfa5a2ee6e63cbac41da3b6dc98544a424299eb92d7e17002c8a79d0db1103050113ae8d3fd46efd26ee5dfbf6889a6675da4556a78e26f00626036009bfaeddb8fbb67d067492ad398c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119cabe66865a7acc7b744b345a32c0f5ca5732bd02d1dfa52ffea1d5a24bec05d05a1ad056b36f879b3990a1773061c3a5f82f28fdd2431004d7af7aa95009be4ede1a7cfd1f91d717a92013d739;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1424d13acd4d58a243485024f9cc0d5e17926a0bd50962ee0a8e105ed1a0399a14ecfa0bfe400a66b31fd82f6aba0b3b28bde830cf69fcdc4380ceb784aa494f370329972ae6356e421a86cb13b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcc320a3a323f3be2514190f9aedb244c2455a9e21082ab84bfb6a9521e9c7fd99ea76f5b207423af176089b133bf16e52c639bd64ce0949bde6b9214b89c12c52863920526b2429f31d60c74294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb4d0aa51ea96d852a82b48d34ffcfd17c5b9a66103626ec5173c799c093afab9c9df6347fa3dcc6a7c97654d5f4e8553253dfd38c5110f6581f881e72ca15ba28a765cfccb01f876d66fbc68f2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha542eea0c6380615ba010b710e41de080206dc1f946cf4b901320f248e776b0724ffae2432bf5504b67cda7a3a2bf1bfabb2aaed11c3678f6c9e7c1ec1eda04d119e7c6521ad709914601dcd196e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1473e820c6efde04eb3840c878c2c5c2fe55aa82b14a4810c71064de800d4aab05a57c811bd09951ba683adc093083209d0bf6df671d026a2ec48fe0d161a410149d9ade3fa5aba595fc2efdb08f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa11ee1f43961202fb0e8dec0706dcba7efc358ed6d94691b444cc7f74c1356d047e72f5c180f62265b409d8be1e44bdc8f6c2e353f259c8a9e3ea359769fc7649fa5cfa1e23239beacb4347cbbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8859f320b4c76512e4c3c3440da07fbd8a3e38e813f6f6baef5e7812b9ed184a97e7d389779b5f6b86f9825db28810cb95289a33ccb86c3591594dbc7d097f3bd150c64cf6874d2b2af17a6cbf54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145fe42dc6eb653225b21f404f03de829a2af8ec1d87968fb7a675458e1ee6d1f151542b530711bd503012c07c0e5d6786562e6b3902b4fca06dc50c72900e49aa3313b41809ef2bfb9c14e6946a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4343b3e45cbf04395203935f91811c0ef6db3d60850d7ae5db02ede5921ca8cc818ab5bea1eaaf42b0268403beea1686c4c859a4115c6d0ad9f88cd7e4dd04db2b3421b41fc7a63a902e6ff88cfa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h151faf8da7639bd6fa0b2e99ba69692c144c0b423130058d5f68b72837e44bfedee6e5684a0e950fc342588ad40ccda5b12a892082edc7ebbad8d2e389d8e6c92d2c4f48073b8bcb84fd16332633a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193ef801c8b0dc0fa8d8e41d01a958917cd1db8580e0ad63c367dce707ac578a1ea270eaf7fe7a12b2211425682aee2a791ffa131e79c62a835417cbabc502c1bd4364c7db87782ff47eaf955a70f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14228a66da156d3d0b129f69d173c30d5d57dbd506dc49c3cd0fca684493ef4de1c2842a0fea7dd78c5ebe4ca24ef514ffafad4620a5dbd0fabd64464ff6aa6fd78e8a6036381fba2cb01506c581f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf86e41e8083ff671ea6132b511f13ab94bec08d87c0d80686072f019a1afcf2721466395f6d1826c056ebbdbf92ae593c5ab8a3a5a87851c56ae559aa5487208e5aa76480060a1f6169bce908e55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f79d7f3ea742d8986fd2be5091555df57d76b2b5d62aae1779421efdd1e760bbac041ebdb5291b1d6d34c45e9351163cb28fffc4085d508aa7b2e6a5ab54b3100635ccd43bed1c39f8c18da589f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a266df5301a43b9e5703ed1552097d6a6de74e253db44385bd3dc13960cb61da5916c3b10de9ab597afec5b4f55ceff29329ed37f4a8873e30dbf93cd06f440e787a25a8a1da23ec42df7d3abe69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2670a76c2a8e492999cd89b22320f305efe601f41ee43fe798653b0d9b5c46309023db0a60fb3e41db52b995ddd61d3e49eb6344ee57726a7777e5918f3b3dbf5a8597b3aab31c7dddd8dfdaad50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16144f9ee8d40034bfbb2b97ea80febaea0d238be962600d0d8cc2e151122cc71842c74afc2e48b70d738588bd636a43f1411825ce68049cebfa80d8966196108b6b15923c6fd9d7088010c9a77c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebe640ea30d088a10f8d0e57ca92969e0e76a1390a44f2d4c06639f928e0659a4e755ae2a5dda6bac84d21f2b5125ef44a17bcf3198eb4485a3fcbd684c21504c07bd6708cbd3d32b8b4b2f85e5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3e88ce157431ad9516f0df29eccb083b1c5afff85861b27fabe39c83be0882a532fcaf10017ac77b0bd5259259eaf285187280a2f7a65246a9d2f3e408d9999129d954a0ab83575503d93f0c512;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16110cf412a3d1a750ab7c7582a24a11af9d68473ae0c395bf2190cfa46718ef25726fbc6ba907983b961746ad105bcde5602a55ac9ef0e16f028f4935ce1aa10b3ee5f5b53344ec42af6bf5ef63b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d2b9965bcf4c05575acfb46f474a2828c2a31e281b64d2fb3cd956c2086008f895aa15e2449e4f20a5203fc17599cc7a26c668b8bb5e2a1e4eb1023371d83d30b31496c3d2d8eb2823884c4568a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebd80fc2e4a98baefc7960b79270c65127efb0052984e69ea9275adf4f3bdf4f149cd2dff7a1e71ddd1e5e92a371cb93e9f65cc9c9160319b7143bda886e05e2b403587e2950653ae8212f079c56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e585a583f4fe9d225c13c40d08137090d4a6bc9f92ae19e27a5b82822a8a9aef1e53a4be5519170374f0995837d09e8d8dc1670be469c56a71a267a7e7dd1896541ba3a3b32e153f050e631ade79;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7d412e48729f67314be0b04eca45640d4605677055d3984ee4b47ba58fbb13d23c13ad69f7de45c54052c24670be44531cd63c568cd95d547dfd8301a2f8d22d1f0adbeaeee57e28159ffe95141;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1424fbbc126a464fd61d95c50516b532678fa3f5c055921602784ab8198f0ee11d87551e66a542a9ee0abfa474769c4cc9bdd7fbb5575a7c72374a8a2b0838d0bdfc1b22610b8358c792f39bcf8c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21f923d3e21d31bad948fb6c6e1537be45e9d073d048c50786af13efc730c7ca100b8dec80cae7273cd664e5a1dd0168d564a3e16fc03f3e90410f6eba60adf48b67b99019ae2fc675066c1a78c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17aa4058abad738e2baf623783d8f5abb34d8da7e7087021deea2ab9de91d1dc6000f41456511bcc8e232f74f394ec60b996b00aae068559b79a1341e56e32f835e6f93e5b641a44acfa07ff9dbb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b46d6077f46f818adfa51b9801e0e0c3372e1dfd25baeb2b060524c1427df34f9893556b4c5716392a4f49706555c71b0ad3f791d8a9fee3816181c610a9163c9ffb4a13a9453b9f2b94643dc19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4075f843ef7ee46a3c9810a60d8d6e0bfc8a3ee15c2d4fabe29d5b953bc419ba1e180f6f8c4e01e12373818cb2b80e2bc58ae15cead3a9d114ca7b730d88d388bb7a928792b093279bf61b059466;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb06bc2cd4bca125be7bde0d35467abc586ca3a51aa9dce91241fb1397960686665fe83988252826103672299f166e5049abf919ab795a1173b017f504753b2983f7888013902d7b2adec1f1c98d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had714c19b09349b7dcb453160a386cd7a961c777e7881443a18437c0566c327cd515519751b4a4a4c8fa06b7dad0482e97a3b9fcd1ea9afe1eb557e66823bdffb3eb491c93c545e18439946726b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faf128aae4f390db0fa03289c25ecc89f62286af848eed0eb4bdbdf6388a915993643954bdc78b21ccb2b3f0f5d7e1dafc94633662fdc9d77fc62ad9cd8ba77314c52ef38372888619f8d777e609;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4fc12387b0a271e04caf323124a26842d130cc620504f393123bb758cdbbd33d0d138a9463838ca01e80e68ba7129417bc6dc39e00674c062e6d45f18c54e3395201ff5d9ed11c546c08ee09660;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h335bdae61675dac318d76f2d477a9a3e589aae1943e6c3fe9706993568f549116d9d48a89fa713d29a8e55bbd7f477e0478982de570106f5593ba7d70070edc5da251cb4d385f3c76a73248a5d41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1404569af7c49d8a02f2c18394e3b0ab157ebe480d31869b19140a42a463f4ce6add76ccc40fa17a6d19aa163ccc770e6c345e31fdf0ac6745e662d089c06797fb86029765afed5de5f690d3cb10a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1624befbc89ac7e7bbe703bd76dfd1204077d141b9be5ca05352f9e6e59ef51e1df6e2ef6516e7b8543df9537ffae8d67784ac8354b0b24d1a470e72d4b7ef20c10570790e5205a7565d864025295;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9cfc5a7f197bc79996c1fced357679466c67056f6f38141167858e23aa1875d654eff2b836a956b3c62882589feea632ac20eeeb42ccd0d604c273f8ebc9a174d4829c28a0272c810d675818e0af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eddbea00f4e59b680beaf4be8d98473232b83345aa0af5070d232ed913069c18828cb59ce3f9ebe90d5894eefd5f7acdae08f6f4cb219cd13e9dfb1706ac69af0de152abb50b8a1af53ee0270217;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf59fa48f884eed9708c10ea0c9de81365fa9f017329155646e4a854f7f9e715c53f1b805e9592fdb941fd12de5e271120159213dfc38fca2f1b395a6224c236fa08354bebcf1892452daf7763cb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a810da5e65f42936e90ff93a3394b68b501364606f0320018d9c7918516a4796eb4da7894619bb17b8fdbf8fb4d508bd54afd975d04740c1258f6045f59fb1aaa0bcb261dc769f58c8f6bff5e56a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc20379f978513a79828f76acec949f409c942a78929551ad1e34a30e3eee18fced95c92944865124ba986a0ab50aba54cff1c805d43d04ad62e61a1457826534951cdae4351909c106b671e3677;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3c52ce384efb3ac3df5c021aeae2c230937793d3461f822a1dc11cc5daf0bf0190a87b715c164589e8ea76446e0b7f941384e8776a5c7a5eba8e33044e16a693c3009f1ccde44c5fce5eea0fb4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6a5817051c2c9f87ad9295fc8be629f283761827efa956fdd8122dd404294ece985db9d8ccec1ac6c29b38897234c26196bf0a9b0be69a5d5af43c19f0ac3ff5ba6b88682c9e2152d29745a53d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b82134174434bf89095ec834eae4c47a88b7f329e42a25ca8c3da15574edad2ed99d6a0becd0abb144a364669de258fd84f6e7d2e5faa024033b00cd4bc935c784d633483c91f4c7acf57b2f4c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13aa8513f590838e32e2b4b8d6a84f076c20cb9bf8b3bca6caf544ecaf10cfcc21501517c732961e3d43b409efc69018d5e39db6ca0acf00a006fccee5b52576e7f56a683902130f8518e1ef329eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36d06d4da40017d63ae523f988fb0d0a062eadd13677e9130fc7acb293ca0f0d2e1f340da337d317e1a01d5254ee9a2b8c4874375a6cbb46043784c322148c155898288f64efd9a4431a349b1dab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb85907b7303f17842c35985bc3eea4548a7351b7575a134868f68b935a31754c5f4be5d9176c1628901082ddda382599eacd7f6459bf2f5f829a7429162443d886fa2453c175a22a99ef855b39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ac0e80e4c10b4b5b093623a50e4ba92fda6440cccf5a050f1e7bd973c5aa5d096bd78b28b8724c4997eccf1aef68f51bdb1495711f52f614fe9e5765520c0f3dd27c807c972e92d69efc6946207;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bcba6cad6ad094731581884b41e5770fb7dd51fa413355aa55e3a61e181f15fc22af39253621fe8d9043300e6f6db9898e19352fcbfa80804440fa9e234d7c70befc66c3c53218ec32fa05bd4f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4aba4383d2aef8b66b228a07c32fe71ec00f376c05fb6d02d8289f04695b08f86a7f7944bd5645d5b0fb0bf96367773063c24b5672196c319f9a5530e70b41953adb6bcbc50a2954899d42992fe5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12344ffa4f9a585f6e6b9e5aa6439a31e7eb7d6b2f0a9c3aa024b7142909261b51f7c20d8aee0f3abf9a26834f05c84d5069884bd1bd95ef3b1f3dba26eaa69e94cf16a46a4fd17eb16cb1569bd97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71750c237723628f84f93ccb3fefb68228039896cccb5e7062bbb548fe40a4eb02fbf29abc21ba11ea56d3ba5b7fd409c3d32da6495769c22c1c9514256d878ab0ff498439123b709634077d5341;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a32a45e98f4a85b13e808a8cbba2563ce48926e0940420b6e8601c9c7f3908d6a98533fcb6a9b117f11bb611641b831670c19de5f66625a4b0ed223a46ceab4082815ec9581b2e78ae0b2d49c44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1545fcc5bd340b5a025841f6c019cbf686f1a20010034d2e3a9133dae59c956cec5ab3663bac6aac35c5d82f614d781027a21f7893f4cd150d46cba867bfdcd1bceeff5e60a762d036d27d194755d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16099712de750638c0ccb6bd162851a03213f3aab808d098d150b227f760a005596c6ad8d7f681e2ce8a36d5ddd5efa5b5eb131e69e9053b47537f87a76f233647f51584ac080eaaa437fcac62c24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a58feb589278f1b9d25036de280b31d794be2e7434ecf24201c88d0a48b0e83d24932114a53194b1d45d7c6be665046f6848ae3ad124fcb8787e68bbdb4ce9aa631a97e85a2f48e2e1ed567daa6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ad0ef638e72bfcd9bbeba63e966af61b0cdf6e7c170bd7a2787ee43f5903201b19c78b088d23097e07b2f45852cd21223a7fbfa56721ee96371d9c15e2f0fc895c7f58c2f966259f3299eff9e70;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5af42c7397ad5560e4bb02715358a5d035c7505b746f77fd8fba8aad0e7d4b9661d0a59ea65319ef9e3cf71e24c4b9710a0a81eb2b752564e4be6a8be300944ae39dc5370c8db694a6c3add0c17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e399be6cbaa5d943687b43835b701a0bb951f84c3753a7b81919c53622370fc138556be237ee36e3c7f4a7304f27ff675425f0ff4c19d182df7bd19cbe5ddb54542f1ff5ee8ff6a3a429e5bafca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fb230b4edd78fa98702065112c6cf591a649a281a3d214554f6bc46ab915f2202b3043ab94f60fe7546f27f2fb7926add07ed2c83a36c98aff84b2cc5c20f1ac59ce4baaf467724f7df77be63a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123b6fb9d97693921f0c82f4547d68ba89a27151afa15f8dbaf8e0268c76e7ea5c460bf1380c7af34ef4090fb9f39780f486d5ac837028d7b882506a16ef531e9bcd829ed234f4bf55f6f279d5e4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h535dd039cbdc6c3f8d8039c2fcfc220477b219fdf8ced312537951af9e59aa2bba8f212ab33a35013898f233d33a39e77ed8eff9c69d838aaec08a041cf27abb2f48afb24aff99bfbc70ed78ebfa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he11147fdb3dd970acd9f691ab585eb68a056e87a84b9916d3216223ff27bc412ceeecc878a36369b5304400c201721159fa1aab008727d37e32eec0018dc5c5aa74aafb4ba16a5c17297adfc4973;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17404200d3f3b868367f3daa7da5b84c598f698e7ae1fb1e01b8c328c8d207628a718b0f4bdf88fdc3a5514babe63bb9af5b79516e76d8f27079e55419eb613c4f9213eed6d212c24b62ce0edffc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h993fda4821deb97a437fd8dcfe8d9373466f266798768526d492f2bebe4a76483c0a2cd25c9d4b1bab34fa4496ceddc70dd93a0f996910d120d6376294d4ced8004d222e1ceec2c1ca48fa03b9e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da39ac3b378d0b9819ae9954c9bbab0dd49db522d1c34654f6c8e39d4ef115d1418bcd0d6858f9b1c9535e1a2fc7bceb71b128da3ce77d730ab0fade9be4d27bec2b49ecbdc2fde91bf1f2d92986;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb41cda81d9b564083fd8b5064c9d7bbab7dd7e787808bfdb84d6aeae223f74648eb898046124146ee5b4306745ec717e9cdd7ec9354c09060862ecc2245facbb809ade867ae6f38be89eff18bf36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15441906f5cd4f48291d65a289a7a35eb61f2f73bd06e9879933f61fc3f7755363f29cee8fbd03689717423847b18a086f141d9e176d32a54c754f4da446dc53f002ab3e9ec5fdb23f565fe8d12f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2d21f9f2440709108f4970d9346d99ffbab6b87a0c5441fadef6920c56e4c42d337173ac308c448be18292e1debf7d19ecc0d682677c5e4730070a46b3bd46e57b52557862c1ec5943cb9daab77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a511f47e66824d2d5fae26c11e3410c51680a43b549d46120f7cd40df2936d284bfe4e0d5a192da1a6e1f61b583087a96c333720b7222a74b6c0944a36ebe5e52141873b9483da9c0d0f1de0467;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18946f3dc0d0f434a1b28c6a80e4d5de469be0e8b804fea4cf61faa9679385c4659e117d3237fb604447a5dca44dfdbddce3e75fcd44cba51e0bbd917fbc93c471c09078005139563efcf4a07586e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14331b499ec619acdf1c53110bab5ada79b840cca101acd7b8e00cd7edc819a47ad279beb46e0b08175996fb97207c172c1d685d5bc67a0a170add50fe481fd18fdf6d933d19cfa289f8741c5d8dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h993e56e14fc80e89b882a30e8356a5a88afd9232cab3bba7ae93bc9607cb33faa9a61b5a7f2054d8c09386b9f25fc571e3e7f0d9c43ccf6637a2a0eca099f2d7b2fca538095046498af17c7dd1be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc74a96c6d9b0411bb0b5b6b8f5a78490daf2ad5ab31c9cb3e56631df4fc2dc0099141d8944ffbcb20e55206fe359b5843d93dbba9a67d70a66ed2f5d385c056c635e3b6c2f42c390a8a52ba57d30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cdedc397e8340d98adadc7e30bed581b84ac0f29bfbfd239a9e4b8f8f0218866ec0458ba4290ef9b10e8e6030aa4baee30a4d4d1cdf41e2ea67db766befe40d2ccf9ac171ac91ace89476d2de7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h435771e70b1b01b56c366e60a854ac0147308a2ad832fb81fe493b535b9470ee613eda9090205da779230f4816284f06244661258edd24a4125966eaa1611e6b80893f26701a7cdfdf26f00ffd61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52995eadcdfe5726ec94209c1d47d27a36061a76771dd67a57b2426d32b89bf0ffc81ec015187513bb71a49b6ff34642b73b5c433b6f21bb2d55f9f27bf55862e2b10d36d3da0cc60732064393a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12dea65fe7314df272ec5153f89cc3af9d6f57fdd0d140d4e2a59406d0058e4d6b87559e1d3683216b27a079ef6ae12040f7fe8f308edeee67c42f7096b0d882cdc27ec12f0132b175d3dd51ce517;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef558c44170aec65f783a526cc3a7519b27b81c31d41a5385295ee1adbd377692cd09f116a3ff4e6e830c05ac24631e6b0c810e2fdc26c47e6040ee8b706e3e37f6a351772104267393ad489021b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcefd3fa473e419de1c5517d3d27677843c1a7341640d6fe2e1888273e2f28e610b6d9722828ef2adcc38a4f39e84dfba38cea228345a08ea9df0ec8d96e70f2782ae2c7a6560862c9f490d6d2aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5307b42420448f0b2d5f570d9d3c3b72e995026cdad194b2b4f0c4d5a941ff5cd1604d6a56b7f8ad9220789af65d1b080f27dbdfd6d987750b37b0893f722a1fdedc132f8d203c2e504093969fa2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c64326ca444ba249446eec85c546ec9406610f5a7aa145f7aa00045ffc10e4631616ed39997b13ca12a162fd479644e394038e4baf7d25b4c937cf133ba1932eeaa0e94c4a2d324061592b9225af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha315c6f276eb0a089b320d2d8eb41449f9719728078118bac95b49896f12ecfc04a7a48bd75f9a11f61b7ec3fde24395160539d42c3a4856aca7852702974e3462bc7309fa54c80e89d3953c6a99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5714c0d6b44ed12af401e6997bfe36ac0398d9fe1c8665eb6f48db407a6978317e684135932ffe4959bb048bf7aaa86d7956b3731fdfe7336933efb449edc2fd3dd719834443fbe2b7f9cdb27359;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab16dc5798f6a325756f6aa43659b260b75fde16f24a906d5006aa05d00e54c2f62034d81f3e0a1514824ac35ed658144193dafb585e260dbd23ec5d02a92b7e9d5b24c1b08dcaacf7a0410474f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h925a313bfc72946bfc3c60b4460be9bd1f19228dc900aa5cb2a9eca6f3e9679194a5389251f3879bd4ba6b9b4b0ead515145cd65308fd1740c977395e166e6c65824af2fff4aa6075f9ebc8aaa1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c0e49d7e1d07264d626fa1396e4527aa472e26fe7c576cc8c826985533d2a47d2aeea8780ef8844954f7b4301e6d325174521937982139d2573cea49f0b4f0a19a10613b2409b715fc7bbbc3646;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe35e085ba289339eda91247495ffda387625b1cfbd9ab0dbba0568ddc910c10f210552a97c7d4e6592e2f8091e824637bc967c1efd2957627fdcd74f0902a3cd1350a91217b7c5ec34e2d69a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a235dfd8c69e4f623b2f03aa48693fe7c600f081e724ae6344096fc5873868f57964cf04559a42e093247b82b8ec1cf4658dfa6908e39347851dea8db9daeebbf8304952d0712a3a25b1946fe71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a4d28fbc28cb0d984cacd55678addad2981963ff75877db2132ce91e75af2285e1b599f5e39fe72d7341e1785047a0abfa5bc67247e30700c7b689f979243ea6616982d351c6a4c895d1f967b68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cfb5e0d99575ca4ee7e5dd11e19edc21308fd8ba4ff1498d80dc5eebe8c7e617ff828261e7f0fac4d3d72b00ecff612a4600967e633255c33624741aaea3af65aabe1c5c6fde34c9393d4472f7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d79645757971c460e412df0300426c5957917e06d7612fe239ad98ee3b00918882b12d84daef22cf7338c2772b0e0a9b6229a09489239c609d3e8b40416a43cfde95f34ee0bd9396219c08d6dab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5578a731462155ef3fdab50f88cd4bfdda1cdc4a971970c590ab19f5b1a7b22ef75892651cf28e088c6ee9fdf7e5854039675876095c99794d2cad3b18e79a0ab041bd8c36acd7fd652abe5047a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5704f27c51eaaa7373c88adba08a82b0d567827ab65234a553d55cb8871e50e19b2daa44d1017ed22dc2cda33b115cbd4f2d5b645611ab3f031f74d059d25ae75b9203c2e092163136257bc273d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha16f99a14d55538e18450717bd68637922be0f56671bc83c4aa98023b79921675b41779f1374d6677eef5f5c2e6dad63ed7230c11552cc961ed021de874e0eee97dc657397b321172c87146fc172;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bb3994115223c1890793c997634c2e091b86e56245af092424482c024f2227419e459df2a12b105167f64ae8e55b55c5cca538450b95f674a5d5d3797be2b20e08c57543d09ad7964afea671d58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he78be89b7927a794685eb2189eba7604d8aa25cfcf8c98b441192442af5c4f7e364b7b1ae82c036e51a789657a5f5a0a051702ffc0c4b76114b59fba2340987ea5d83aa0392dfa332cbe2f6a72c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec3554388147714bdff459be9fbb28963f80796aaafb3914df4b7c4fc43e505ad377ec8880277f6a733bc481a31207ba2a2673dfa676ec675776c77e329697f6d218580ef449d9266feb68628612;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb3ebbf53aaec1f5d46ddaa8b1ddcf1df7f6ee969c89f7478cf3d1e4c69e04609d62fa7372cbc9f7a5da2bf28bd4c6712cba3380f5ad7f30ef4285e9e5cae04e5b5614494edbad26322a168ac16c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4cd6a41483bb17e5253457dda391bb4dc3b8109df99446d2f571004f75248769e124b72d12b1e06cef08df4935a711b6246b1a374a1de47a5ff010d1eef1c4e2fb3e09a3a8e29304e14a0817b2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf0c8d842390717878f7b5f003115ecb6e2d90f53481bbb5b58d5bfb38d5751573c8014efce99eb1a9c631d77b5936f7dcbcec5201fb986649ad70d317942fe58c1685035db2658b189dc441b22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b35444debff8f5b04f470a9a35eca1c0b42b0fd0e998d88961a2884f428bee9469b19232fbc723836c6d846ef07792923d1626e181cd6b7610816d73fc040139aef4fabe7d54cdbb697a98ff30c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18463157ffb91f3debef0d4d4caf91c2f49072cdbd1b9688d94d50324c5b7f71fcfb1463a91f005f8055ef66bbb6fe91d4775b232a623a072e30bf93451b344ea7a215a69375444f62144df307af3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14cc6dbcfdc537c7aee5874a22a1916d9201aebbebf2155f57f555ef8e157c45116e821455e87d04331e235483beb34d58395a1313f16bf768da56ae2c6dc91b7d547b7db33dcb221e35e6f5bcba2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h156f9d81ffc2a95c6e2611bb6aa1a3af811e86a2edb3160bc5d633c2f7b6feddba05bab2caf96af1153955c0b24be7afe141f92dc79b3099f68337e2c74822772a25bb5f30df116cbe43c9ef002a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa9b57bf5d35d61739e9fdedc46084537f7fea35a79caf954c2b0f580460167f56670e3e0d8a8f2a6b1b39f3d2df0361afc84bf3ef6cc02484fb35e1c57f6e27075871643b398776ccea18920f19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67960eb30d6bb7efdd40405b23b25acd3f2b20439942d4c5ce22536df13a821b187c2b829569b257a7f26b1cc3877605812ab91079cb19e420d87bec04b35da5193dab133681d38e8c0768241d21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120dbd88ecb3ec7e288f74379597a0eedfdcd9987137f1d0f49fcb07ad3675b413e09ec2299d91264cab146199f441757e815d992897f4c629e85e6675c1e671167830af08fb5e3591bc42ddeac34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda677bc31511ca6d3133f5b44fc412a1ac43e0ed22ed87d959d929570ec61347c0a935e960a9abb91c62bd929f9ec3c1d6e49cf4e7dc8a293c12abd77fda1a13752dd9163d4a22750ff37b3693b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfc2a95098cae260b9ab2a1bb7a0578022138d2eb5d874d56184c9aa68a1950b0a21110dbb48deeae0f498582c42a5f9bd1d18cdda75b1d45dfda704f387f7a9e04e275535435f1913266b6b77e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9aedc51ceb8afe835ed8fb78acff3d7386a5f9e84bdcf5436e853e566050843ce520a94a0470c3d8342a4bad5399fcec86429215d29960ea2df16530a5b8bd7db69c80d67c7f0c857ab072e03342;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d1235e6ea9f5927a236c310c53956035baf3807e560bdc2ee434e5995c0f905898ac60d735de488f99a42b298f78c9fda9135d8e938eb02197b40eb8a662f066d97bf26011cca3f7e8841688bff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4399a6ffe72accdb141ec5cc86af8b5c5a06e6f11cf174bf83c001c3770d9373d1931376ff4b9d6bedde2c88b0ec97ff47fddd1863cdf44452737f9eab0d2688748360861e3d181983dd27739ed2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbce97ff8bb1218feeb4792fcb579f650bb4ec55ed07fda2005c0551d8eb355358aaa623efd99adf4fa949500eddc1bae5814ba504b8b74a7ea471358d667aa83950934b861dba22408212f54294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16511158169399769fd8b6f4df0da61599b608a7ca7629d204800c3aa2ed27b09fb5768037435b215163252c078456759f61c7e4aff76b2ad2c85ea47c8bb0a7951190899f745b8c3b075b77bb944;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101a44b66f57fb9d59672f2d828a351c0309c557918490b0a3ce8c44d32211a4be2a49c88120e6446c5d074b3f538ec062daf120070425bc88951331837d6547bf188990f35d7f219ec1003e711d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bd2bae2d409237e1b0232a7ba8d207a51c209a7e53f2cb5d5956eda1c37169b3d2701cf370d74543e52087c42542ba0e60c5297c21ccf59087c0a64479d64afc0551852007a184c3512284c9d5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h468b4bac5c6121be27d7200df4342d839ded1a197ad5aeef2c0999dca803ae7d313b4a0c1b5649824c8d5841faceaa16398b56d312c9baebdcc19c234490354a1d183f8c5c6adada6d5c435d3835;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a41ccf49f80ef8712cc27af5c5e0adc241762cf3546d7792d9c8e73069c45b0685a03acf2e6b0191b82af2f42d4ddf40978f271d24babc7202a8c63d3423e26392603e5efecf6a54e82c2333bf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h802aa0eb46cd9cce25b6fd681f26123b56ebad4cdfbb2cb21c0bfd5a385ed02bcfa4f287f298457cc3f9263b284c0a378af072d1896e941da3786c1eb536399acb97fe85195303e008b4d687b2a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd09aa378c078dacbc8f2d72c0b3956aa315db9df5b5578c4763eb7c401d3a33d30d6ee56ca7fbef62eefbc05dd622eb091b85119cb7c052898bb3733d691acd66bd071cba763880a67358c45b02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3838a232928936ecbea8fc26efc19be0e1012a1295592913f303581e9d78c6363c343bce16765384160ce0b8e291e8fa38a6b80c300ad0a89ca5ff6c40747a224d8cef3b1923348912891155010;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1911b285c171353956afbccc75c76ee4d04213e53438d4b431ea496167715394fa2bef070f6be27ab65836501e4188cb8a943449972a5ec27efe013cd23956339490f0b7f0e73ae97bb43fc495d80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb308f249579df13daf0cc5890e28ecc412e135612d5cbebca5a75a2aa5ed50d2b128cd3e6d654da431e3af44a92be0f0af6f161423e80719d1b52c13b480112df12f29e6afecb796f54779619d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104b4853e09a8ca8d4a69588de3efab2a24a913472bec4107fb2d6fdebb2eec3f50f118ccf7498e9e7da644e3ccde762db7e670a4e39d6d79eb4f0648b3a6e02050d1f1853a5dc07b503057e0036f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f48dcd878ff6a3dca947a52049f63083c50e25686e5697250f5628066310b9359056f11e0b47ba90f7f5212258c021e126900a7fc8141af75bf4051e1d8b98d514a0b96581f11f1ba4356cb184f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83107d07b6e7fd428504a117fa810f75473585c9dfbc015058ffcabc5876aa7ed51dfb2d4bed7755a7177e5ece62a93a2e23388aa9f25d80810abcabd7125692341c6fa94b58541295216d75b8ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h522d0085221b5ad951e4ddae575b60d7e68f427211d49565077c67f054003c6a589109b9c2f4ec7d815da6fae445869b9b1a74b6d2ed7d80c3a3a0ba40dc48755b834b878f195c5c0ec4da7c363e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d51d06061b052f6c6cc7c0b9d69a9bc09e7cbbae167ada7f4153893546fddfd5aac38047af0ad7236efd5108ae8ab1cfadb96f97aa0f20d0929aac669c1aab51d199751991ed4a0b4cc5a3adcd33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc73e376a781ea199bec23580bc4791db2de304f67905a3ab07812a8c2ca461025e6544f8f0d7c04a6e353a949b9ede494e1f86734b628bb782cd45f9551a10f158154724d6459d4699198ef6631;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12737d46107b4096839d7ca8bde4e5b2f1d78a7bc3408992a43a4908391e3fa17a78b5b592c231e2148c69964cfe094a417624350ebfc4bf1061a6fad58c040d7184292fe5a9d6e67fb8da1880c4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f1b3df5211b937ef07139513def60e01fda9bbbe3e684b5a374a14a9f325926c6ef61b746f4fece2d1b6638c870c6741fad7453d5c946a6538c1e52703eccb413208fcd334f8f818eb13f02e98d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b83b6f2119f412eabb24a87698731b2038941c11e9fd546d5d7df42b6b7c99931744814124badc551ba9c1a0030d78539ee33aa02d09ad14390e0e1fe6b0cc3a44d9f36db523f12729baf2329dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176f566490647659ae55676b318a90d1c6d03ee5adea67ffbb0aa483afd15a36dc774bba3f029093174398aec8ab0efc876c2fe02d58b8be591e4ea443e1c51ebaae109353fa7e775c0d62a3929f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1309d15e4202cbbd4957ca3594551f0120f9600d5cb81c4a4c2c175dd6104fd08714155f8da2ecc65ad2bdf9663faf3e8bbd7c08fa09ba8436036de0ee7e3b5c166154c7bd8edc6200a6f1d3470ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16afd9de61598fb98c9f6f85510df5d03c3b758ecc70631770a5085546a3b654b51d7581a80e64e2ea787f7c1125a696b1d75a4761fe59e9e6ec071ad66deaa93ea3cbf4298018498c068ead55b16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83080e460ca343874145cefa16fd56874f3bcafc39751b078161f211610d3e0f7e8a6b79cc17fa1d845447d1ffbde1b5418372b575fd574448d612e967ba73b1f6add2ef836d9fdc875743fc4713;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3d2e358d181f7f37751a4046ba7d93a2cacc8fd7e28ca4e6700f59b1022a3f499de7d16668c67668914ddc96a1004bf20e9eba711032feb1058f818b855aa73e2d8b5e236da643eae532e73bb39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78900b2b48a2100a74205ce3bb314af66ef720b860f379e2892fdd4002f548f6d318ac78bb6afaf28df4ecd49c8d3d1767c7ea6e81077ce2f58f8c4097574fe2bf53b27fc82767300537b1c3f758;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0ef2de01143faa77f8dcf4de988a0b761b6459f2e3ad7a0457da110f52fc74c772a956474ead9e08fb921d837991b7630cdfb4c1a1108694426312b930928c7e4def33fea163362efe78cc80d25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bd3aa119b576ad34247a5c34aa93c0cca670079de4fccf627729ada7b390f7495600349a1c06615afbc229f0a0c86dc59ad3e102305d110c2b890a54d9d1a5b9c1afb072efe48435531935ae551;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f56350929d69115cd8678c7d0218b19c5ba30b48744312e16a877bb296730ee8c4d08ac794d134f78407c6880e5f95e6a21b2929c2aa2f6639ffc336c5c32ecb21f00c91406a6f7ca2f160a1e7fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10324e2407668a1d2d12a57bad6c2ca2d4da7b44d9c82e030a0288089726573cc3dc909940452c4b29420e34c443be66aef25d606adb0e52985b52ce390f6ed57ce5d41bebf29e0a8bd78d5150748;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb66d3793e436b89c6f846f1d5de6ee23949820852697e9d820038dff042e60b9fc96711ae15c64e3e4db2e67ac7f37d3cdc2878d165248dfa0afe46e561220916dec08c22c0221fdbb7ff2b348f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d659bd69966800089f89c9d8e9421237bea2e8e18e2974249f8ebd9a3604ead5c2c70c9002f588f09a96e7d0674892f587f396fb972ec6dbc24426dc9ce51502bd2b2a9383f9d2e19c66194f1aff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1edecb4a5cb6409ee6104407d88f1b7fb8cf3bb5a9a56e903be2d64a0d7af4d6ab2c240ebf799f8c9fcdb20a27a42cc039a867b8b19e051a046084bc5611fda382a31e2e28dee0afccdd134c2cdcd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8472de2328f3999bb5a8132ec831166f28aced7ee63fccedd0eb9f8497faa7222f0d4fc3bc610aefd2d94c5a62152b83805af24e8a58060c1a7b862dedb24f451220ebba046bbeac9e5911fc287f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1416f167e45f2334ad88c084303835090a57cca24bad5044b34546a359110d888935cf31d2276a5eee8427c6f57cc1b7b2030d1fac69910c48c200bbc447f873b6e96329ca57db087fc996be59164;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e84332bc330f058eaf158dc5dffd33a198e0480b3c8fc67c0704d517e18d458d7efc6e976fa387138dd955d1d94ef0f884dcbc35e29652a2c284c8aac3fc0effd8d912b5f7f0c6dc7e41c929b5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b988efa1994ef4b16d4de68071924419d1ac7ca2ea1ea4b4b8906918b3429cd0099fb1637c6747ca846db1a35e7507b0d6df72b747c373a75d5d17f19f970b58b2c0e35cf13d4dd62be1ba2509a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f0b6b70f79721ab6ec02dce2650c28b04963d7ee49de1763a80322d53cbc545c40fd9a3e9041b678d405e6b19c95cb835eb1b2fee038f95dab1dfae72cf552692c27e2d2020162f577d91a7b67e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b96e892003449bbce4bc453d3252563cc35c91beaa67e451c7cb7d90fc2e41cb8196c50dcc327536e06ed967b759e64d0ed60bb931d82b92990ecfe0a06f6973eecf2dfd24471b956ce0b8e1d0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff0c01b3dc8f964ec460eac397b609e202f97f281bc912fb315da29751dd37e4f89f221369bbab6cd8b8d217a5cdb21f0e4ec5114cfbf4e773a857a05cf587e549e28266357f1279352c7d25efdc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca98ede7144ec7936222cc7e6b924f8b0f22e168501b37b35328e23e5f464092bda32c3c6b26934886e899dc17a8024866903dcd676097bea89d8e04a962f67e02f61438281d7fb4d246adc88f79;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1433a64f726937a46fd7c53999cb533f819aa9776d6db347af5f87cc86b89a7f8426f1e1d5ac774e3f3476d6337866ac5f3a21d25d1c6443b9dab9247a7a85e3e1964ec8437de1d8530591e60a7b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9eb37d61a34c4dca8cd707f2595ebe93b172250487be24efd53a3485188ad22f92c087e57f1930e58e3fd96472228d420c06cff615a2835485d2c46d163758b0295ee1621b20464bfdbb86eef6ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b79de27af672a826fb44e7cd898d23f569a92798b8741c70ae94483cc94eda01fa31d91e89418698dd448335e10c71d257b9f84bba0b73433a5396ba1b1eaa5f9d4ecc01d12ae8f41db03a82a323;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82f6d93a4e8a81209c3c19b550e18b03815d3d6c0f7536ec53aaa5a4636ae5111a1a00e6022916606b9648d400cfc4fe4dfa1b6d56d890613974297e79e2fcd0997e2265ed22d83a51e5cfe1819c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6d4c08692e0e3edb6ed6cffecb68f0c2e79a75957f6dfb3474d0d4119e834e5ef3d2ee0bb27df6ab971e9f5662b89bb54ac4b3f30d5ee4796e71b8cff7140e2a4067bd4922dba670b3c0fe2d786;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd401faae13bca46f69919cf68704f440bb6bf87d2a7a829dd2b000a0e99ffa99944d2d0bc39840a3c1fac488440de2174c212b79f55593bc0f4e290873ff545d03c40bd9dac11a8a10774e533956;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f958472784cc070ae7d7c13fdbdd24c8434f15cbaec45a92dd1650335aed55c68a371fa767955d9c52d281542d77b5571be23bd4fe8974d55d54479af5b897c4fa8f6c49f92efce6904cf279ca6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdea066f2cc6e09e120f3ce67e9f9208b3f2bfa93bffbfa85f04d605b370dcb94c1f197361ae1b169224dfe2c4e001b43cf8f3142d56116e4f0ec6f9e7616351dfdbd08cf461dc2b2c8f47d6a9bd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19269ae9c4c9a8ab7fb8a3898fe33d1e14d6161ecfe57ca12b25ab068ac63b4871fb3567ab182283fb30af946bc68a0055a2bf629f931104bdf69f65add1ab3d982a37c9377745ca2591eacd77d3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf2e13461fdb6cdd9efbfdc4610c639feaa83dcef87fb03d136b32ee3c8e4f5a337a4b5e520cbb8730764d7eb3c42e3893ebe185d06419baea0790ee3dfc4043866d5549edc85feb5119e2a04a03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31ffd19184d3ed218d65f766016a0a6ff7c74351d464a8965ccff4ee7e3e67b2e6f0cd19f802d53a72d9886f07c14713996e45c020c797603bee4adae90d1dfd30f596e32682e2393de027617bd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121b04f652c0ab989c6869a6f1fd29ee420c9c3794a5148c3b3e17076879ffcdcb679ade107249d167c419a96a0df301db0b58e21c1bbed650d8416fcfc269c1df93b7f127fceb4ee1e8ce9bf913e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e643f04bd0cab59abc6aeb88e8b86a7a8a5dfc409ef32813b7749ee6fc009814f76d5a69c350d0b5b95887e9c16f43b1be7e4618285c04279b96a4b98982eb1eefc7aa97df5745f0ee43a3dc5736;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1931bc7ab4a35a8a80b435167e09b23d3afdcaf2fef6fbbf908a54980c79d97a5eedee4109871a39db419c5b4c25cb5ecf3d99e024fbc6d1a85cf38b0abdef8dc818b69519c6acd96b1eb29bb27a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11aa3cbd015ab0a63278ee187743d323a483ae43534d8eb8a9c0dbdb384812593db44903c2bc07acd6f9c84afc021050ef56a8287a1f1b8ffde8c152b0dd683b808650022d425dda7fa6b002ad13a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5479b7bc7cc4d22ef9fa70d587903505442e2935e3291b870b2cb21965b83539db5e230d85a9a971af040ec70af928d6c11b1afdb5b41e7e9858b9d55315195ed02983f6325f4c5da796afa9524;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13475f9257c96eebe6cdff0b333ba0418322e6156ccc37c58633a08683754ea4aece8e5c196d086d7d35ab05765925b64872dbebeec452e428fd26a59cb5aa3decdde2b04ada8f88ef5847ad04f3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f97081727bd700b438ad23d4153a9e6e24daa973f546cb9b20d5042e8422ea68ec90ce8da3a3a25c37e248f1f758de4be58f0406ebe7dedfc6925d4f282b4e2f5217b547ce8e90a7e6ad0c569e48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h272f1563bd25cc8a8bfd5da4d6567aae8bb468d2cb566625101f1388bbc42d8eb8543d1279676d715afcda6370a1a3aae193a0af4f59ad2aedd1cdde10df84d70aaed4291df069c2850063ac358e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4810d01a63414bd8376b789954322c2a060f49c4fef212a0b341d459d79731dbd9b78935a654a2cdd9e7416dc4f98d9733dd47e791591f7745dffe39354dcb979b90361ac3a0168f0838d34c8db7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd10f57f71041dc1d8ddfdbdf6a1c141b852da5cd4ef4a07d41d1df9d60987b83cf40bfc548898764f9b3988e63a8e69d66239e63b130d8cab4711b189e64f3a255671a5dfbbf67c967659ac0b4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3601401de8f4cd52c6aa21797564bf98be6e36382458c094ba3a673657bb1507e70067df1968d0f2e01caf3b40cecf2f7277f516591ae6d1c25afa7834b1e9776ffa3851ea5c9641d62818ca041;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c14c46cb63465fb564108c1f39ba16f54bfa646e7329eb1fe5fa1f445758d2d0318f279e99f8bd60c584e210881e5a4364d3dd182501dd5f9286fea4a421e9eb368cbdf5f8bfaaf6a267e2b88ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50eb953492bf0133a60c39e2a70103954104172a42e864ae52c4db225c9362ade13ec735e3e3c89395a4a4fbf49b6a569c0187fe83cda97f6a3811f75419fdb3b0e8e56952899efd82b42732902f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h938e0afe4a18b057aaf182261ff33ade6c2cd526bbe8c7df7f8250262b2512d98b8d0839390b37046803ced8ee5887de2fd3435ab901d02fadd83f0001bc4daec3e2358219b18ddbc7a2b74e5b0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121b5a69cd1b612d5c947e7003560c6bb98181e56db2d08aeae2bfec66114853db5c25a557820384a3efeb687220c2f4d78949ead08bf18deb27c6fcb0b9196351b17e075862ef7055983c1865d9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea1c15a499552179fc803ae2c758ab3ecd770309d0cac89b6ee4f6206d90ad1674ba4cb5cb9cd1a76a5072d78c3e655530464207d0a0516eb9f33b28c0f20e0288784a70ff5addb2b07ac9d0085c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h550c7f36bc6028b98c826dc0053b70c643013440d644028674d96cfdd8b0b4ed656835bbd2f4e523e14bfc30eb29ded2d61db3009de0e80ca5e37ec00b6acb6c934037f61cac2947986ece9c5fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h51f1dfe16852375afbc68ee8dff6553fea9236cd648f0f6f1decf9e61f71dc007598633535d95319f3df72ae2c755ae9b3fcb7aa2831f64b5a50c6dd9578ecf8d0c25a0dab32072791277d33727a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46be7b81d62919d77cad6f103c1472d6a66c398765b6d8eec267d7a7c458100ccd0b5bb07a3f2c53d8570ea0f13c9dd17d13aae839435d57c13929abe662f9e776838cb55ff0bbd690e6fe9a5fa4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h884d016236ff9239e9df18f16c97f7d1552270e5f8a720b20e68fc4f90e7e1786e70bd4ac358d836f70c1ef7dfbb5c0e6372947fb21b96855c6a8c0a3ebf42aba6dbecf4b453c1888d9a117716bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f10a96beb13e33ab2bd3ed2a3737962b036fccecbe06606d94c4584a6f70edf7be7829801206227a7bf5bbdff488f7d6bc32a149f0be050960ab2a20edf5091c3be6a769286b241e37ef9652f22f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c923b1043f4d825b4249232ed8c4f94490e118a7019bd0cf5b71db6664e5ae056a4daa57f493d705444c72790b987516e995b81b3e920adea630a080491068d55a9668b4fbc72b64ab91d9c10f01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa27bde094cb486ed824b9e1c57cb2e528d173117f70e8e1690ec866d7d918905caa8d0d56d19d7f409fe88385b84e6761a3cda4716e90e34f1f8876306d9a652f55d90d3ec8b4caee711ff9966e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e73ace02e01e4e7073e35dab2d525fe4d89b783b180004294ee44a91c1ab03bc1cc210c670b1cba66932eaad14a2ecd3ef54bf8f349688dc8ce4dd9e4a395a0402f24149ebe97963c484d07bd8f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1923166a2ee1a5f8abfd4e354cd44521ad475808e7c07b1d1dbaf5f4ec67642b0183fa9895ff690bdb67ec16b1643bedbc5c3bb06fd66c75e4ed229c61a07d49b686245749034f6c49532d3825;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12bcfdbcfb3beffd259870a1c600d94e8a747ee13501070a01a47809904ab56e5c1ec1aedc0e4be1859105f1e3ed4654386647ef45d0f3fb7db5cad9f01eae7ef52549033b3d6d4e7292597f4a37c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f26601b10b30cf4193e83e62249156bcc46f3323f56d0b0fceb9eab529b4d74ece9342b9f1db4ceaa2a0598dd021da8d226d258d87364c6f1bb1b109f8a17dcb0f19b415ae5ad3dfadc6ed71234;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h184935f64c3529d34eb6afcf0ee213f978d1f6a6bd99602aa9d7e96cc73ed1b35291af8f672fca0a6ffcc0f8ee6f7ef41cadc1f0f2e32f342e4582e14facc83625ab876aca68628b8966bd295793c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b4df8b8c2c7d240da491c5113fc95aa88bc2956a0211288e31548a92bd1fe2e80eb0d68193b812bdada152592f5b9630dc25bdd3128dda70e09c6aca9e689d8004a96d436a76d3cdb06c229ed53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e3e6b84a6185f05111763658fe02bcb9a5c18ffed3331fb4320d73d98e760ebea016b6079dd20c0eeaaf50c856d753c1ea0a5e759a36289d0eff539d6a4f60936a6c9e3f09535d58c82c7a035f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcdd2c0394a8ae7fda6e55abbe416135e71b8a92685df518089ba260cb6e7c9cad66bbc5ced53c65f7992c407ef549579c14e46b448d351f6111af590670e4011204fa269544700cba029e0e6827;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71644f8406a53b4becd4f0654c6e27377061b89776eb845ada50b6effd5c66200731e94a8e8c4bf95f0c226ea20b32430ddce0e82ff8f5cf78a50c38aee33cc4efcd0a07f7e74bc1d23083d0e98e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6183cace4bc99bdb6dbce7a5aba25e1923439bc99f8e9ab75a192563d2ad0d2ff1e6df568dea774bd96af5a594f317fc69a702f6255423865da01c01078ec0eae9d13f9ac53be0d95e55b129e3e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6044f9b61b4f8699ee321cd9056f6e5f1c59b96df1cb167b091997e7ae65102751193a14fc1c018357550c238febd01af2d384150ecf8c69fd1025f9f1f65d292bc18ce42add09c86474d2f4524f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179ab272831b954130bb7011c2b68e7bf283b8a150f06837f9db203ea2dd981c6086188bccd41ca16997717b04b5984acb538dfbc23f6648bbc0a1eb8260c610f7d2e6b5725456a30365a41c1cdc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b352e06dcd42e8823768873a73bd3e6891bfb3511fd6bf243aa8d32fff0f392c7d2050fbe2f38ca77ad92461af7591f4620e6b2369e848e63b7b5720940f4caa3a852dbb27b12490063fdc62039;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16209e854993779a3536b5f348d8176665d7e3b24c0763266007c57c0eb4ae47ac1162775e880b201806a01c78b5e6423118b3a15964ba0fb3fdd40b76f0615cf770ddcd6c2c0d40b58b13c5f9925;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8343e73f4ee5cda3aaf444a7657be5aca39edcc1059c044a88787de52750fa3e8890ce2a46d4f0efac9472fb806f9ac389ec5bb7b09591f9fcda7bf44f1db38614df660ebc0e64a460f06f2280a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b023cf4bace87413e21a627aed3b9af2147096317a50fa61b584d3b0f8f3a12ea39e80db69f0ad15256cdafe53b9f1e9ad28a80204b4313ebcfe047b001a03485a38a98bf214ce0756644b525d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bd503b6ec059c251708121e525880171aea3ff94c1c495a222a35d931ef0d72164d70fa922fbf74e4d037e53d0ef39ade62835ed73558038bf69b93951837ab9a1a942f401a5cc5a1c14e76cfb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heaaf236f321c96a64250551df24bf6dc1a56a9593342454edb9f2fc21846b00e828e99085e63d061e123f05431b5c06eba2377045cf7ba87c7bab5fcab647f9be58f1ae57942fd4f7b668dc9fd18;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bcb463441bb5a1a37baa6236520ca1b04742c0ae6fb4dde5e8a316d4fafc311d772e69d0fb078abc584c452c04b35914ec07c431fad03855450c196647efb97c6a36c025d884e3eb232c96c9a52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3c44f095ada5882c92bb837570994eb212df9a53e767ddec78b036368372fc7cd2488f7e9b20a81a367e2051f40402ba6536cd499fb030d787b2fc0124c6155baebb0407cde3abd1d9d0509b167;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e28259938d366e546b2328281deb4c36df53e3afdb60b0aa58c30298ee1cb9d8d261eb5daaf5817771b32b694167185f8a4776ac48e5522130f32041b7d618caa82ec425a15032e7a3998ba600ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177468b0cb191fa74c0b8e0efb8da1d8719451376dc632efc7247901fa4ab732935a9cc9dafe3efd5bc9e22c1308dc8dde5078874866c1dae8414522dae6a6c198dc5d5a8551e9d817d709eaa1e67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43a4c2b88308ef67b637becdc803999d77a9721d38f86b9b2f5a0febceca9b834ffad63e27fd87fcc759386f890a4a296197e98921806e81760f32b55eb44f9b43d3b78a9d5284d5866bb2e5de43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19176fa0e3680a88304597b732841aeb9d9ec89b9c66b5ea99fd62f1de5cfca83ec364110328e35d9f40312a4ac0cbfcd650aafb710870c47b9fc206621af1d243901d1890a6db62eb8d9e3fe7a6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h151a60a3414c5e545b59ecfc927c17e97a4019a98284126fb1c09e70e8eca0f2470e8c19d62e5845e7e6dd5bddc6da7540b4c0032c2c044e5057f70c15822bc2d9e15a4ee8bc4e137231c613d3866;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3edc4bdf458122a33117b467733d6a1f940d3efd6adc053abd4abc290638bc921679b1b864311443c0d0d685568bac31800b49380d5e101388b4e2fa13260219406e29f2495a8c3d02caa1bc500f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bbcc315c941731ce34bf96ad3a5845024ada9563a5415604e451be7351d6f623e9da039f7e073b53f9560e9823ec29b25633ba8815e1084620441ea49eff67874ac8605dadb9dd706d440cd9b8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95b632e3d8924e70d2ccb72d9914383423a292a9a3b9f566438cb325dd8bc58e4b4647040ffb0665fcb0894e722f5f4ff7fc2bf4811cf5b11df60491b1bf46f5ef3640258597ee93b51f57a0845f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa98043a2d367defe7b8cd590b215319b289d132eed9dad1392983557a627e5df690dde9116be8124633fc6e86b8479e15bded4c3211095cf768504eb6c49f6c0963459a01b940eb083a0b361474;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdeed013a62ea84b49afdf31395e3d4525735773efcebe5d42865b25630af816562f5b740e3fb51b3958cd4c9081c0a5128233bba07887013f6fa53b3fca35db6de096f35efdb1cc947a1d96e4ee5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h982316548ce8b094a992131a7d000a61f34ca7c9f42a97ecc8bdbe6a51fcfc87ea9247ee20e4caf6a6a378c9214b9312ca34688d9b972c53838a677cc83eb0026e8d3f1466d74c238ba67d439a44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81c0c87e5f44121ce778e18751007a252d7493d361325d398cd82ce7623395b6b792127c57e699453b9750c62852de2b2fcc29c7c25f4600afe1eef8a95f04cfff241673f0975d218f845e8aee9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd94249f35532ba14c131fbcbcbe194efe745ebc5bc20f6e19dee6a0e3ab249d1e4de56ef701987716df7bc1d000d9a7214aaf9c570ff036d532c716e5222a042948179cf9ddf390935b22ccd7b44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4561d9a750397bfad51ecbd1e8c49572518c52a40e253f0796516d9494b04631d5e2e14a81caa512dc2c39917f77b53315a6be2506c9b437493a5eb33b6171dbd170b45129d9a7d682cdc5985b85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9045bc5f396f358827b884427c6478b817bf8b037f84a1abfe741127b9953993f09c480c261d10eb0b2d061e4d7162ec9a258036379671222fcde13796e79c3b56644b9110ea13e418511e62d2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16144f04731314ef2917fea51125969d87fa38801b84a42d271b3661a19712991c8c75187e2caeb3f4a2049bfb8bc7ae7a1ecf5f45064a2b16b99548316a450d0b2a9169c0a1e1ef20d6c33178c95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122178f8ebd3213b82d216baa25bbb48dbbd813ab39e80b14df529cbfc39dc37b05f7a049df825dc5170b7a8dac316943bb6bd2365862027c525adec537c14138e9aaa508bd9b009da4df9b45d3fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20a707765e68edfdfdbb037f5d765529d88ccc166e83afe5f5bb435d7ad73138b1d78792e039a13bb26bde8577a9d9affb7520553651d5281c461f0f90b17c9013e8eb4cbc503241ac4cbbcedf5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1220cb3eddc148c97428ad4a9449994658f19e53a82f1732d3fd203accfcc1dd7ea67994458185c9d756d398c14cd9936422086725d3c7deb70e35ffa22e4d2db52b5eec92c924b9469f95943a84a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6d5205fc3ea5f56519e39ea2b1d46f8c6dfd83de5eff084f5de7ce0fa6c1c2b5fb81c992ca24235f22512c409e7adfa26a9cfa328125ac7a28b04577b60bece274b173b07e8f739a9d8de978402;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebbf96caa32b17c726f07fe950a6892aec401967adb77e4b5fcba363a211b7c795294fa6c9fab17684df0a90ac1c5089ca9dc8c12dfe370ba9aa9b2c90152ca7e13e221cddf2cd24131cf5c5d3b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ac3c6e78bc1fac9678fa23b3edfb09c7674285b41ba609d9ccf29df7f9091ca89a3ba201ecfc96af028fab9ff2b05153e77c4228a1a252df9e9a986260d13216679b60baf74c2bf74ef5caea706;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1817251e6c89815170efe495e5051e97389131b8e25f009255f30cdefabf9a8daff700f189592645054e907ac9342cb24580bc2b1c54561169f26b220c3fbeb5a131a3ef30c1a1afda3ce131097a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h345481a63ae7d002372376fb70a45183c1c481ddbb76197b45fcc5df2448efa28aa504be57bab15b7206984d7cfd18a90fd93ab2d33e1c55744fd2c27df30b8adfcf06c1c9a8fa7b99235cadbfbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15aaa0a790d9cb35213c547f71c24500c94615b33f00c14185bcd1e45876316cbf53e3e30e3538fc5ce3f696060f4a7dfc13eb8a393fc55a84a2848bd39b02e139a46b2a4f6df80b31d0664058bab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127da54d0ee0dd4e9c97bed3af3b9b0cc041ac4dcc87915b4b0f5c432f8ce9546adbfc95665ae70db45ab05a0c97ff33c0a06687896d3e9c839bf3afdd98e6358519afa4d7877e10735c12a2c83aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191f1e2d1e8083818907f7e9aa6cd4ac295d953cafde5bafc22598be96dcd2c2c83803b6e626aa281ccc8eda5b2ae490ab2f2f3e45a2621477df4da256a14c755a031e3e2ce28323e91053d44eb1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf32cee9ce873eedba77c274b8323d90ee4d58a139b6bcf1d3ae8c2713ab8eb02942ccca979414e491cb455b946b3aa368deeedcc0d1ef233326f86dd33c67e7d057812b049907007bfcbdc4b4aa3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b7a51bf8cd4c0c764c566d157061c41b4efe501e366a8252dcae7381108dd197c4922e1144791dfbfe13c2789c6910342e15ba2a9153d68c242ece38a7b73b64536f0b3faf762236d911886a1ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbe57f44db5f93c3d5fc6dab860bfd7d3e29ee3f27df8a5e50bfecaf522fafdbc81cb2e651c809480ca7a99f0ed78b1b6a9092038f28283056edba4f342cabd2bf16de23079bf26280f7ac767265;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197eea20881b8e503772370b6cd4f0fa4b3315cc662fea9de4d40764cd8af068cabe3fb7c8daac6f7ee2925ebaf70f33b1d2ec721f85e058f61e33c82cc502208e30d07e081bcd389e335e5f62095;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d0f4c07fea471327216a98f1124b2b1e2c94045722c2b88281c34ede5d6b5951af90668f2ff37eb51d99d34f6f572b0e2041e900458ecbab0c9e2eff46a22676476523824ba5a48f16993918281;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6dbdb04f77b489485ec4e6bb68db243987cae2a8fe699351eceed84752eee098cd1f0e04c7bd91b23ebb128599c2f6db3fc103f273c0633d0315d11bfd70b9ba273938aee21f5760bfd6e2c2104;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7922dfb1496bb8e0d11bb09350b46112d4311076b345bb8459f76698c6d617fe4c6a4e2ce9ae1c34082483e0f4a9b2f55bcde282bc6643e52f8de00397322e4487ad9ca1457d8824179f5b6b3b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbce892eb9a07d9d5a7479690775c1a8b3ee4d8ba23caf4424c53b056166e4bb5df0c0a16a433149f8b8ae929af16752111bb75f50a3e9801d2c5e6c0f25317777d8baaa84ac690a3a0745313b6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha14219da820d8359a77a82048e1aefb07598bc1e49a64d71166940d3bfd08e00e02d7cdf191803f66c198d726480388bc074155ea739b097c2d998a4bd85d582fc9b9d712a3b06497f8a7f079b2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d229ee7d3b61ea9471b2ec0f4e27f64125c9edee13db165bc3b29364b8f34b8ffc744ae89c403c98b512f32b3a69c43f29d7582be70755eabb537c8a94f277d2ca0df02e8714c0b0d1fd1cd78239;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12aee81984e95aea8a2778cb6eef8f17a9bac9ff3d35bdddab5baa82892998efd182517f5b26bfd9854cf0700db8305ab65cb4844a1e78e20326039c6569377553e7c95077843303bfc7659f3c542;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heee33273d6a40a122df483efcea723442ab8a32896c8fd17dc4a6a31538b3aa837318bc6360dc0955e869c1cf2255cd82978a81a71f7a043c018b653087d9012250c0f7438086f4d09e8bf65a83a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba1afe2cc4c12310b43e0d770484494cc69b04d136a0dff4430abc7bf746becf1f55f21e7212a01ac60cda42373bdec2afdf2153119f61b6493bfe7d53b6ab68dd0f94cbe2f8622a566b424a74bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66393bb76ed094b3997dcee174cce47e8e06981a2c5c023bd3024a116fc9b7885fe2c7705e4ac69fb81db22f9f622d3f54e34e82bdd5acadd4cf13a16ccd4d40f9d3e406aa7c1ff6fea6f6fb1f1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6044f33c3a31811fbfdb55e1c5453bb74f6d38a658c08601583cfb0b86db4e644db37649aaae8726409b3846cad857967d611c1074fb48f6a35f5cd5a799cf6ee86dcb7b348cdd030eedecb56b75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb797523fd4c09875f581e99fc7a6dfa14fb1fe3fb156611fe045a4c25dca1a853834e70170984a571eb1ba500c66730342ca74a4a5a2bc8fe2ca03ce731d1266d67bcfadae03a545f898252797f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17cc56ee9ad9c1d669f8a007150c4715de60d56d3d42a3ff3481719dcfa702e8e416c37a73e341de0178de9a971d33b798e94ff16ef60a0680993155581a51ac19cb79b7c8317a37fbe080856db57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10666445a4f8673f66ae3eeedcb240bb63b43092ab737cd8fcc68fe66bd9e2ba4f5628976eb305a47791316244d1736effeb185dffa9eabd7093702cc11bf585909249c72850467091aa3da0d6c82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ef647fbf87a561ae5296296dfe069b2a93dd24cd53b39eb0b010430ff790bf25cd15cec0485f443ef5758d56755ea9472e13060b87c370119b23595fa2885b321451ea9cad6c8b1c3a7c6c4e07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de39e4713b73f153ecaaeb07bed88430eb3ca71b86442b136b2de63b3bb286554416d49c9d3e5a6cdea838c83ad2a9dfd3d3040016ab64ed38a0026da7036cfa600513997e0192a08619e848dd19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dddc0f13a78601d3b7582e7de8716102b7cc00474ac248d90072e1817765ad48ecb42e60f2b7ca8e78e07322f8586b6dba1ab169a33d46d51748a16c1973f4755b042812d0d1f45e818e2048580;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b700acfdbf829b888961e5c6d03262ccbe3ca31183099e03f7d786c053a1875474b02b9bc7b55796199a127e5b32a1b703078aa34bb8c497cbe01f297990afd0a65c83e078b00bd38b6f45a72319;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a24e03ff903dbc6ec68f88e1dab9c2da42d5ca0129c831fea3d4933953bfc299281efcc684ec914d3767b1454fa87a24c8d8271bb10926932542a65a11a9493bc323fbb92c820dca372ef2b8ac5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2cf6c8de77e9e01000818e482175993134768d189df38375753a277c6e62cfeb4fa2f313762b53549c7573c6edc23566fd1eba9b463894d837ff61cf40dcac3b654e5629c56cc0aca573f94eb83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109ed907e1d35c7d90b7cdc0d55e59b040f432b836d9e0e0027e4d80aa6e4d0b9b00094a3e0d6c0a71f85181a36d41d4f68f5b3603550fade5da494b1bd5d4828a62d1801a0dc54b59c16409d2567;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c17cee21de95cc40f4c126f1e0eb4ff2ac9792cf22f1e9d0d23caca380f94b6929be48016978d9a98afebe2ce9fe9f1de50658dfce22531161a47bfc597e70d7398b080fa0121c3854fffbfe636;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21eafd2970434a59ce2ae0623e18ec1acb8b7f55c7b7f826a4360645cf83587159c048bf0a66000e94fefe84d90e03699410fe1a6d0f3797dd3630ea77d84dec68c4a06fbb37a6c0ef0e889a508a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b20fadf4c2875f9f0a3f3bd98b13c60d81725dd21ec8bb0e251bfa3bb1318011d114dcaab0583b7dded1f9db8d4191522ded886da3d62e076af7703c1353653de54f43ec68b66aa86a6f9c770e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he75b3070265641ba33205508a64c5b1bdec83702de689800e3a4958695d209a9fef04bd3fa38acedea2db80f926788bb62ab8d6aa99580664bc877a0633a289f394cdf4477a327e5649bb585eb96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8778971053e6db423f1f34bb8f798948036416aa1b68ac75f34cc145584787ca762fed46c3ca61777fbc424185f4597397c2e3f1a22876dcb844d9fffa45a46b30f37cc90a5f4659c25f1f22fbe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d81a640ab62027b75f9ac68ba4fcad9f549913d652e24de2cf07a00a093f68fcbc1def614bbf8cc876e606316e0d5b545da42dd0c0e2a3ba57b12214f3754558d005b998d88ec1cd32b9c3a06b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19871b3ebc7d3b2322b9db343acabea47a82b51037efa1dcb841e91849906048e2c7e59bae0041b6e82f14bd19e94c6d7adcd22e2159f8d0c4ff2f47125be7c21b9b181fa79ed02e5a4ca5172f4b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc39cd2f3a1513d5fb8aa599fb12a7f3a7348b1006f3a198a8ac8032bd7741f614014d46061e8862e0f064619049556c98a134f30e80bbaa83a9430c610c777a6684c0e2ba6e3526884877106fc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76e61a9cd90b0787226c4d5f370bdd1ae6ca88c3b6a9d5b4250380ddc00927127a1a3253a2d1bf37897ed94bb0bc6c6683436e88908fb0e18606f1a2857442ce9869ebd98ea759753f3dcb636a3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ea1805cec3de16b9964fd32fe776ae6532c8588e337bfb8f6fcec33d35b05eaec76975eec058ab10a4ec07670403a0a818fa4b417b51b72acd320b907d9e80c044d2b258fc5bebe02a422bd6b29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b20540f6f1ebdb7399846fe9c5530473b64babea8dc5891a2fe8db4006c28610f3cff9bce7a0ca0d5677b12cb51771dbab1ed572de906e751725719ff58878044d7b5a26538ee9642cf70000797e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db953ef4d061e7fb632c28b938ead9413b9ccec3da1f4f075105c2b8b51543ad502363dd92a476e06a7f50bc79c27f62e183c4a27b82fe2ca8e024698c0eb602543d448c6e0cd04e704d6d4b92be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb04ce2318fc848c5962b8a057d7a6ad45a21db63c834e4876053c4a8e93f89bb6ed0c5adee9f2e621ab5cb172f92ab210e1cff9c6c83be4fcd79342359f23f0fefef657b01bd2976133b850b15f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0d1dac6515f9504a282235f9ae3684d1d9a94dac624ab01acbff4d310e12475e02d4d1a63472ff0b088c7a807b658c933e5d2d44127d576d6d564a0baa8ec089a66568ea14271b81cd5c6feece8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122ddb56cff4f74e9909415e201fcae3c7566ccfeb2902f57829a331fe144b1697ae42ea9922fb264bbd8fcae5effbef9487de0d13806281b0e0635404c16daec4636a697bea4309e609928fc3da2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9aad7d73f49e5ab134b014f136575b63098b229e554416cf51a77ab95f55a1310349d2410b1e840e3809edd1d130018663d8b52ca0961d6e778ee4732f27c741486182fb48ea4e920017717e25a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1247a7f80895483df6448ff1d772c73fa742bf2f775d157d5653174e7c33c85aede35e981a5044d008b02ff457619b6f84c6bf6e17757fc8bb82ccb4ce48795f7cfcf58819ec66d7012c67bdf649f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78e0a6083c44ced0de146793ab5509b0d332788e42308f1d4aeb529372d91bfd1bc42de32513b9379ded12da59633cf095083a8a67be942ce4d8023a439a7aa19a06b9bd6b4179092565c6441f7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1410f4ac8de47106ee74f1bc0cbecac5ea41061de784f3c0f579d88e19a5b37dd39aaf9e1771c86475d42f17297d5a664ccb62f06d22debe2b54aa3958bbc7680d7d152564274aec1ea4f9651541e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191c9a5df4dda152c5e4c0036be24c66cdff4580af8a65ba3c77790be786e0fbca14918750cf4d1b947b00fd78b242811d5a870be5f6067fe3f6fc0a61fb5282131281b16f5d398bddb4540ecaf0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6ed1d4a0f72ecafb502e65ba14014bbd3659e194fa3f4dcc7c1fa4422326cc4c2a6df2235b033732e6fb5f9154adfe06c601d1878439b2f63bd8c33d0daa43169140c090b1dd3d14917ecdea3b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14092acd2645752364e65299edea2c651ddf39d9b150c9be30d4f879553db628ec6ae2421247e3b07e11c9e1d54df6ef6877d50833bd62cb31baebf39b33d7ee865bd97c8bc7247c38f001a3cb12d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16eaefdc8c49e4bf4a09e97f74ac931ab6b021c8a01811d7f2ae5606a1a2ce0e24428578b7a338343cad4346a9e78177c8164294191d89fbda9cc44f06ee704eab83ca18bcfc80941258b73450fc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b5dd9a66001212b9841a50da174ac08fff4b03af5374059f0d84f8ffc9b425ec87d1c72aed37e64aec379c473bfc3224ab04d812fe5c2f31d8c10aa8767c326efbbaa38a469430602087700d335;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f033b5f0fafcf21d5ae70ead68c5807433222845e5fd947e3ea785b089c7aab17d75be7e593bc09ecb4da4b33b7eb92172b9bacc34c642d67fae90c9d82a518e534ff312a39b8889b2932e3b6d70;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b5ecf501fd453f0715f689693ab988dcd2607f34e8e69e1e7938137f40b5d2b4a0817862c58c6ad94a81bfbc887c0a128ceb8383e55cff5f348cd6aa1bc1d1f689ee6cf40e0c9a75f276bcb63a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff9e6932bc6dec5a7441e200a7bf55b31d75f0e836bf7d2a983f8ebe86d99bfd5185a1c2af2063298e441029d3bcf6da0a329a3e03ee0459b9fefbff1541359dfd6f324b88e5d565e33c6a7c750;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106f2562aca33184562e0d41f6f3869f8cd409194f60114cb2e998f225d9e533c3281c7e7aeb373de149ec378009e60f8334786019419501d19543d8e59169e913d43ffc687cf85ef17c02ba71737;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf0fc3064d12ffd0246ebc9504c6b8b048e491f147f0f62d566ccd03d796cf8c10770e4336bdf3b554750e55ba1732c2c3e8689af9e2dd7f0bc865ca8b41146395c8f93e78cb3f07533e7df37e12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1109f56ebee5507eaf1f1446c2eb0d71f7bc6ae7e386db5b14b4ae16e71f7c0b8679d03acb9effdd36028d1fe960ef4075a59ad57900b0247be7da4b388583a00f11291e0adfea862dc324a440f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h618df7cdcf3032d308433225d4233d5b4257136a16607fddc426f2620ffb67051f70d0137f9896011d8a3680b580bcc8294c02461abdb8081b0cc5e8a50490a821c0ea7d18c2cdf51a14f1d1681d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f32aaf85b5e4563ebebff39a6c83a8fe15ceb3172c46830ba48275796b48be01b43ebfc5a87f577bb5d8d05f47ef44bf247799ba8a8e41f8d03782aada7f35f0f907523169acf7f06f8b0596cee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1191bf60614d5f0061ab5d57a96a48bc3e982a52fa6caf341356705c93f9eb621fd82b5e3923039a52a9959c129fa64b050a39f9fff92ecdb480a4f0b1eaf1dd9f00b92185191ad671290e470bd41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c9720d8dff495d958e03cc507d4b966c0244f602f648152dae2f8a10899eb7bfc63ecfc868206a477a26a0ccd2d0a7d662880066afb3dfed6a0cdcfb29d72939a839ec0821f440d13a663c94bae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c886960b07b60d1c0ed655618a62709ecd7df4a2088bb0b0716a070569666b75ed292b836d8061390918c4d440b23b9359fbade9c0f8686a80e8a8c1d4360e2f9145867d277b77ca2ce723b217a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180d9b7e883759a21df6422673855c284dd62a6b94323ba742fe0c395282694d94b4ba34b25467815e789b1b7563b1a21ded124c64a318ca2782de53ceac778aaca456d18e9272485dc20bcbea68d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8306c3017594c47775474b56e45c96b5cde6641e3587d4f683ae0138150fb2596e47afd8a39d09478eda5b2430c21ebd756c021a56b07086b3d34bd06f1c0b92553eb42c091d4dd79734df579552;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4930662add80bb6df25c7433ba37e8f9ee2b690ca929836cf96c39507e02f9b5aac5855edb65d533005acb1f52a3eb776cb5d054a598139f80988d0822444e53b1d0c76553259a8dff15720881bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe1db2b3a203558fc84a7a3d959ffc1eb00ded7c337dd6ab4d6390635f28bb821e2d5922040a4965b33a5ea93f84ce529080e9b3b26c461db5b2f8daf6764ec89e4483d3c1540941f3fc5b3aee2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b4dac31ef12762aef69033f8e5f52bc3de51d69fa87346636617605f413284f078577a8ddaf93c6f0db22d72ae8097cf0b1ebbcba306714154c64a1bcc28099c6e927f17e4209971e15ba835410;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd53e9dc1d6f033861bd122fa37aa8643ca077b2bda40760df3b7e23c9d5989d3ceba862b878912dd71236d0e7589d1ac809642b6cd39139ad32962154be2df786e047e098e8293a5b8b1ddfd4d73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8cb05cc0633246939bb67392eb98fc873255938436e51f0390e95fdcf68c7c72399282bada1094526ae256ee1495f5ce1c95e63cb5cd194820de9cc107deabac51eaa6bb1fce324dba40e1df213;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c0a1ba1ec4cad39752554821bcb59218588e00295dcb3b93295bb21e1b665f4723fd0cfed996248bb0eb93cb2413f6aa7af4e5447b0336a5f43a0c429aa7eb423c82f663ea8e28f5e8a36bb0f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad53a1691d3bd26ab09da341f5b3f5586d22cede7e7c84e5e957dcac23868c19921253854c1fcc924124af8255d2d036c992d983997e65e768abad32797543ccadf52da56b57b8e82cf3a36923f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79bbab717d1cfcd6a1bdb575e5bf2206ccf2cc3de66a07b3793b7e7f249bdca357a4465797d7080a09b75ebb99d7e8073a3ca10bb9610270e769b0e06963935dbda43f1ae9162eacab4273ddd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf94292e26919994ad3191c9c2566d84e7484f47b66ccfe63a4356097a0d9d17758fafe3a40df6adc08e6142c9ee13f40513b08330795f441fa05edaa6a2adba4359c79c0e0c4d48d267df7d4655;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hecbad9e8b7d98d46d173472c68f52a1cc7eba52fca901a7959d7c88517b98a1bc5877bf026d71d6e7eb41dc78670af34ce0e95f51fff48e64268c7eaf666b4a082f9f399da2056aa8fa405b02cd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17253efd090a5b2a1d9ca5582f8849f26bce4d3342a5632305feca2e5e5e091c12472c6067e7f3903445c424bd228450b1f205e8e038cd0174f87c69fea330bf74a876717ec5017ce75869377b86f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc5f8972309b79dac40a50042b1afd48be70e9399484d6b2d7b5de84873012130b4f09f566eb59e188208d9aed2142f42e35de2a68638e4dddd76f8c62affaf75f431074dd8c22241935442fbeee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2e6dd27cdf8bc39d1ae1fdfe5dd8ee8a3f79f4b86c3bdb5da33cbe9806b694b13524de868ccb779c3949298e7a44f324ec14de3a15ec5c2a0be416ad717f6330f02088ad67780047006527d6cff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h739b141e94531229e25029fd7554961c49829146292394208f2934d537efac46ebfcf20e09fc13feddc815eb4ec4c6835cc736d0ec52c9e3887acf1e9debe0176e0e2d160cdda0b8efdfc8e9ada7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1de3bc961d337e6e863462248946ea1500c5aa4571ea0ad7ca80f567a44d8b68ebd5ca6b9a8e7c06fc10a1d838e661d10ddeb6e66634a331bae6356192a74124a55fb1393eb5d103bf6b4ba087a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a4b87d5ba151514396a47e89735c404b752ceca91fb494c9a334fdafc2f8d36767f8b6c61c94c143d109adc138367864490bd7f9f9ba210ccc1a7590c7c01ad365b82ce1f922c6cf631ab07c4a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfdb6042d8915f1372676808a541abf01c5950a11dbd14732b6c0c192249df9ae798f94339d364c81c6cdf810ceae4e2d7de82e4a0173243416dc71d9711aeee23ce3c2b41c910d4664f7de41641;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d653b0d99b26edeadad53e3e3f18118e3334055de023470178f4579e681d1d937ec31a942a360826504fe154e64773eb54234f92da1f332b1bf7d9136aa10a4ceaf3131ae98d4dd4df3a5f5f1a4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dc94b34006c94fa1cd0828e80f9f24486b70ce367799489dd659a2934f95296f2578304b70926fa1f6fb21cc1653b3ee572421558f8e64e5bf205906e12b1c18b283785a4010f283e7505476b77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a8e3b733bd865b0f862610fbe5dc21ebb4fdaf835cd36397e22bc0ff1f88985eea73e512d6c18c598a704c1f7d96693b35de0b84c32eee465c962701db2fd45c62bd312c0f51bc1a0c89d60126a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f76f1b562deaab52b9af46e8598a5a5d050e8e8bc7c608e29cae9da5a03240f22628a30613958934c3c0e8b481fb134f11e36446a0fe8983bff6a9481b0df60c1256293d495bb3a1238a31d3c0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119172665930bcfe05bd7a4570a977b29cb6d5867f04cdec6d9176b99d344611c18369ec6a7bcc3c57eac52ea5fb3f637c07c9345a7d30606ba01e08c30d699a3e9a0a4bf0a45f2e97c6450f45a62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2750857292572aeda465c4d238b88290990981ca9caa540a12eb5feaf662c35773c8965d2f0c97b3afcb4b2f750d9a23b926349c51f15f97c87ff047348705245c77979c14dadf91167a2a4bbcdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bc21890edbd6e6f0b803a35bf3abe901d777fef99affb33be5755bb2f029de7c4aa435980a72ef3a4a5560cdd866ef689fda5b15e86e6539892d669e8eae078bc9bd709ce29d133a6dffa25e8ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c3692eb93638bb637ca8fcbebac492c19f9a297a1bf2af68239ba1f4b82a9e531cbb8a9b1b87c6fbc5003103e4cc90387bc0319d769027fab78bcf2cb5cd038812e665d639530261abd18d4e6d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7de0dc27e2f5abc6fce3fb49891f49094eb17e2ef7cdec1f9d4151188880d6af91c4a0a8897b797ac557add49e3ec4d2cd0cf7183c70aa9f285fa37176f379c00ce2da9c8c916504b97f390c2b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91f5b13f7a947e5830d77fe3112e1360f37109eb29d53221f370455b4c0b7d7d9fcd6a99e7ef627727ff26db47bb45bbed339b8bf57d31f67f50e9d4c0efd52bc6cfb6bf68b722becbdd0b6f144d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d592880a7fe1d72221713cac5eba6717a55cba0c9d1ff9cbf5f6e56457d469de59eb41af0bac0a4df46c1c0d75fa68acb951bf2268402a91db804eecc546fbc61d670489ab9906c80ae670a2247e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c78050304ac6ab61da4c2955c70ef77007e6031c1133a4b083dfea538688af9a08a0b7ac560808583befdf701fbf42d0e751e81cd98daed2efc4d2eae7644dbde50d055355c85d7a823eb222c0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18041fe7f381621a496ecfe8db8835ba5399ddf74872a8b3c2af17044f14ad2b57fb00fdb1a5c6e9c621ff4c246549913817c0fd005665307e2ea64761dfbc1e1b9fa7edbf8208962f1076e61874f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2141a7053b299bf866aa0262e3b38b9f111b42b0ce227facb949dcad5329524b9478e427ec0635125a428cb7fed7fe5f019f335e225c6ce58c829b481190710ad7f76977c9900d04f6f22fdbf99d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e31da128573113530a44a40f94c685d1dd3fc28f06bb068982e779e8120f0a2f97b98b4c01f45969c8eff2c3b77ef8f50846a1e359011dfc1748022a5f288a5760552c73d9bb30d499a76c80868;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162e87f3bf251a71143d32319a14f93ddf818588bd43815b9b71ad87630781cb1e66a9bba0eabbc979146497abddcbdcc5ba5107ae89c29d68f9758da6d6628b69afac12861f1621d8baf3619832;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f81849ebd0ff04d3fd5985a0bc8a54978297f1f333c86c21f8b20c9455664adc518f3ca1f4145e17bab37c858a5dd107c494994af41663020557ea28d02f4853dbae30c644fd253dac2efa8a4186;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13851c9c2c86a66179d9979c661b74e9f4809bbe3bcb01c14afdc8f52f7ab99670b09d3c4e082a600b74faddbde4fbc677be0c0d92487ad834e315be53ec98257fc61f5a84e42adcbbfbf13451683;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb55be16aa3e9ada7cfe521514b454f533f7d637aabc17177ba3e10f488224cc613957b1e3148c36dbed3fd7bad049e1a422c5936719ca71992c8978a63ee103cd4cf00c3be41e6d05ae4094bd4cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4545e5cc22d1e8a7843653b706e3d5ddc50eae01b7f82d08b5c40fb12096aac1b2b82b0777b252bbc5659d9996f949dbc1f1cf0e5b9e13c857ac86c74a9e214f43542af34c75945228f61580023;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2348d5d02df2a74581fc84ee6afa8151e6b72df991118707bdcb2096800ab7ae31efe398856691d6110b4d07620b0453a09e4973b205ce7cd2ea1b0eef8d537f80a3199c0bd0a09979616f34eb09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9659926fcdf094662b34db1cf58c003b54b5fb3b2f50fce5bff2c85d48ca3fe55db8525d83157b50ae541ad90071bb9a262ab866500957e4efc582f64ffaf6407c3851185896b87a97cc1c1937ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72e1750ce59bfd22790d91e2b749b66dd47878591d1c5bfab3a6c7ab97ef49c461872250b131bb8d9c9ddb1f377c47eafc97802abc7a6280d836e70dac8c7ea02d314a76a9bb874cfbd7dd61be4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109c9e025eda17a38eff14c640c03550391fc188dff9cbcd8d27dc08203cb58a898f0b5d7db0432672c7d3de4b6fad16bfd1edc020e5c6b5fec195c74c3abbecf8c978834793aa9880787aeb531dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1345b139fd152bb6188182136d99bbf016e3a33d4700c6b4e735d5d1638449d1d0ac1ce672766612a9a6e2d6200a2866bc4db01e496083dacf7853afed8a6c501e0d31f42757bdd3c7bcfe3e0ceb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7916721ee5c88d08f62a7298c2438d0799365dd1152801d2826fe44e1eae1a8c8e0d05aabda21a06c5832c75f673a07de11f644d41d941e5c6c46e1a85992fc53563ccdbc5b60dd85975e230766;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da179b957d187512fdb5de09f4efc0bdfbbce97efb4606548117b4ba6b62a229c16d5119af42001ed76c2204258dbeb7ce81a6a6ea979d974dd1314cd5f6ffc3f10de18a70229d644e9d9f17e0ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8469c2bf9ed15c97464b01db2f90d008c15177287bd02a39b27b3404b8decde47f69670500f605558eb345b05f880dfa0d0bc4fb63e753c1afa08fff90df835c70a299bafe7731ad1256756e66d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf43a1b1ca33a6c4bef409fe5767a4d17bc5afaa9e10aa32544baac4b8f290ab4ed1f312a2f96f65794c54751e2dc0ea856eca0c94a32d39bd8d744951bbca59776a11f4bbf984e4dff5b74985033;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed192042560355bcb80fa154d702e00e11930de8d66474a96b84c241d5de1b6315339a8ad23e22e1854c762fdaac1206eed1477d72f95eb0f021b5b3b48d3f30f8dec8a2dc111ccf7a6ebcc5db22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf3c92f8388f6d7c4167bd3303f0d86c8f60e29e25133f81c79fd1fca692576b51be67ac577c890f476db795333124936102e7ffa30c1098bc61d7eef29d5869c8f5ed355eeb4d8588b33f535b2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4026472bf5c848e969d6ace0fc31b9de764e747d44d47b248b63bebf084bc9596219cabd6cead08688ebc3c07ed250d1fb11191ed8edca5b930ba73c5c61b5f46eb59433195646f9097a9438ace3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h642af93e254ad22f907fbe987a9efb979903429532a93780b1473a01af4862703b2e78c71cbfbc5a151df263d71d184d2a4f2dafccc2758036e11bc5b802b739f64de6ff6b14d66c2337daa67e48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176dcc9e1bc813861722a59c088386d441a15bb50c00bf0952add6b9e06816b7ceaa7df2ec9d968a6d47f39c9de21b00bcabd6ca5b36e5b691cc41602c860bf6f62e269c0e5e42073cf0f3c7a5c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc13a5bf52e608f987275f2a9c0f3a6f623755710ed42328d4331744e960c0a5b329f65b13a65fa5a7463fc3dc4744be23a4b1376d071e44b5cc0657a92b563aceab38cd8fc31ae7811c93e4d56bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139d4f973d8a8159496001a56634ffc096b079f1ebafd1beb5bcafe7a60864d1d7239f5872173386e76327f153dd89e155076e0f265d764f7b7fbac6d8423339bf969ee47a9394dd8a2f956409d92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11860c11c6774d446083dbf0f5110fa52ba831a7c87045fff10b97d432016a3c19f048710ca42f7db3e69f43993be5fd4c5a0ac9c707c471601a785e39482add68efbdb532579dc93e323146475b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e84a80c5f8057678f4abd4e72d1d409d008a3b1f65ab569b968935b6c203407089ec02b1425e9eb324e63f59a9cc47fd1f4dc68923275cc628b2e153fa177349e3bbb7b0a578e08e64c2228a4a5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1349150fe7226413f78439a100e52b121731f2a65c1677508e85fe9d33f020263ea23f76490050b9cbbd0f5906b566b791382b3ab56e7e4b3736e9e671c05de8476aaf17b46f5157e79ef9554f2fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad455d5cb11f5338ff0490283c1099f2f9e1b36a5463e22f8004e58a2b59a1c60d74df4c70484ffe45fef8c01763ae03777cc9db27fa693c20c852f2fa5fc63664560d64a2fad26a5a93818c8d5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4184c9e484eae0153c438ffad3aaabc49876a171e9bfdb5a5fefa7d392bd8d5850c309d4c0a5e5e19d868be61472f3fc416e1424441affda406b0db6494d0dc8e3a6635a8dba455c4248bd5cb4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19465394f1efd9b72b541b3c7833e3aea26be98df79ee96bd955bcfd21d8e656570c80fc6bf7e27eddad9255e9925d616c194313c9a3424b9d02c7821a54201d502ce581ed2d15f8e737ba62e2a83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146e35cf9089b8c8c3cd6c09e5e06e7f46d545f0ba4bfd132a0cbb57960c18cc2356948cd7b3cee8fc5ee3137a85f5d600c3ec2aa80dce83db938923edf49f18eb5609f3610a0a37d6644e88ed534;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2127b29739910f59a0cc3b963e62cc1077278439f001445ae680387065579245111c7a9b7e7b675a8146ad869f204a638d499c5057c740063bfefab574e2c275720cf711560a2fd09370b3d634b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd45662d30378b5c1a23ef37c3151c55eeb2d33b165c098c9739a34aba5961c1570394d7dab407ecb12c204aeba1e32039be7ffcf95eddc80ad5d8f6eea3147c3e42a9fd5a4c7b5d79f952b3d6df8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11288293c64de56c77597180e2c2eeb2a84d9a51aaae1947c4d847fb8929918c31069d45bae6f15aa46191f918cd4fa5eaad2e719a6efa27b41c3b558b8237f38bd31ce47c03cbee89e74d91fcf89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b9a0e13064644cf6f51099feade5e8ee4d6269a0748341975ddba9ebd3453ad521faa54d9bbdb20607e438a4a96d159c671b1b69e478aff27e8fb095ed08023dc07e10586efe593a67859d96be8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa28429bac220c8a438890b80010b52782803bfb6308cc613b015b28a12d1e93937ff8017720575b96d529b12e33a54eac458d3f9a00564ed246fd460d48bbdeef970f5b1b663299dae1b5795564;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67981e183724c88177fd2dab08791b2e59ed7e750d9439a069ef64babbd9e79bfc3a322beb9de8aa5f5444c6e3fb0fc099907f0049e9759b5d7f6911afc9cbd3dc4da744ef4432a0c4714570b7ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16dedf82dd8c2d65e5aa61add2df075a7865ddc550a923c67adb7a92016d42cccf5c6c3c6890ddfbdbdaa1a79af905888257819129f6756122ccf97c82514c228baa33979625e9f8d80b581a5907a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1468e6db1e2826cfdb510885dbfcff71a013aab4adea7e717fb18d409836ad59ddcb063a12b9665f5c5d927097ba8931415c5fa901a601fa37ca654f86b92b59be2121c2d08db7461858001c71843;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb16c64c2e24a0c18211539cbb1e327df427122f67761d32a7c21822774a858db37782601f8f661a435563b4b0dc1d6b8c6ee905ab5182fde83caa051f4b5a5bd914947153deb47e484c584c0e73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fe12151e3cbc00eded579a7d58da207784b42964d5064e0e50f019765926ac1b1d90b7c7a0085234e2113e3fa895bc2a763d60149f78975dfa791a1a3b8c65b0859ea5ccae75e8612e4bc3328c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff5b07de43346dc7433aa2d571a7e8b60c8cc9f791d2266b28f69d8e932578497a4cc27693559bf424458339830ebd00647311836dc99d10635e2227db27b2915b7125f97de2983112757e94c5e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd901fe0e07b0222b02bd93eed33761c4e255fc611ad7a09cb158086bd1c9bd8be4ec2ed6d4393151a95028403ea660b2ed49317b349a2e5335411b556ae638361453e7d8fbb6237b952128c56bb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4da12aeb8166e22211169d8a48342c3f4f01c2509240a658af8e353ba477d67a45ebb606d6a96791609391570a17419f56efe57fb7948997c33cd80e609218d2bb96948c0f993b1d216b81d1adc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b82b5a1299fc30bd08e1925cdcde0a0f2b42014c14b08b2a9a9175a70561870acaef15c2b9455708870e673195bbda0cfff33434ce12826d4c730f0c31fa5388fe0ba82eee0b51478e7b1b43777;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0ee4df4957c89d714c9f9c22a6a3964294ebd8b3c707126563b06b9bc7cc86f1dce6776a4ee8d8010ce0a4ff7b461af7906d6f5ba0e24b5a5688dc18844a14b3cefaf6150ff3be8bd92a44125d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hade318d64c9ff88dd6500071dd0930667dba5dabda258d0575696eb2e3a616e4ddf5081045df06f9b40ea0f567ed25584c893ba90047246811343687b7ac741eeaee73ed17801cb8975f73b1d923;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37ff47e8a1bd489ac5b926199c0ffce330f5314f465a5d7f4b2e24d5bfd04f2c232918a06714b266490d6856934d4e5c45ec1707a28326fb2ea217e274d4af91ff91b80ee5f2a8b2a02c04e8b671;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a35c4890ebbfa3b3f5ae6b58b8557da7fa2133971683588635e360f8028a17d7c6cc401a09c0570f237c220495dd12de5615c6e00814bb11ba89116d90c4a833a9a369f8034db116d547c6d955c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a8cb4a280996d2e410cfce1e7597205ff6233af921850ef3f4abe25eaa366b0c73e7297a424be63e55e45c5af4d84d64a079da0b702d667cb549d980152cf60ec13001a746edc4566980a82deee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9db5f3ea6fe4443f8290918e3750c7e9b91400320ec3f315f9a49a44270fb6c5040d471ce3351f5f4a3d36bbd294b7cf43391ea55f667b4f946d87538a699fb3b98f2f6c23ee14e3016721d746a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h775881c47bf12cb1dcc5b4e81db7776ebd5c40c535afbf505809944a1c9dbf56750ea643d247302ee9bdf3b223ac4166b8f2fed8bb335c634771a7fbb3a79813f7995e6bb47030efe02a6216c8db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ab666591efecc8c0ae06c1630792192ec9a99c67837076b52834106b8cde076f2d7ff38dce430766094cdfacb213e15515c36999f18dab3ca53602b133d34569a67b6f4e0fe10650d86a5c5254b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117ea85dd509c11f0adc28d064e96483d6021280904e78eba239836ecba5e67668028497086b5c8061f891f59b2a4e8ffc1d0b6cd69513cd6658fc9fc4ea428b2d4e302a4f2441c0ea62716b080af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4d134ce4d742c94f1112d7a6ecf81d644348ac30242dd3b3206ad7a922a235b4442c6f8530de53d16fe78977812ad9f72ad502d75d881e2f7453a6ba4979d40122e6ee35414bc8d8ae7b56fccdc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fd35a1035b361124598967543d1365d6b5f76b183fdc32368eb17a72ab6e8bd22a52649dd344eb96ed6e82565787e4e15df2bb3f6c0e5eff837423452d99a65b6d63c8596eb58a937336e46a167;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85fb92ad6d6056eea3322c0df24a7c9c4bc48680fbedbf7b8abfd1a5495ceee0d548f3d5a431428f9a94ad33e1d069539f14d70b274212e72ac671d08678d3f67ca190b19ba0aaf4aa5edbf12441;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3fcd6baf9e56451f60c88189f2fe0a83a12a30404c522475ed770ec6f0a4466c05f86691874f487b3726208dcc2f391d37cad889d5b8445932ce933eca9b9305d91f11487a2f1da74aac91a6d2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a4da0736fb083acddd9edea469f55424be9e8c5b1f3c0d4bbf404316394ade8a1e70b71bd3dcb26dcda8b73378f2565a41b8981502e7361226d2c39cc1b09f9a298487d3ef908e99dc96a600f3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0e66310aeb7719d051a3f0a7a2d43403fea2f3ee9cccdb0e888352d5ccfc2934979b29e753781473d2c43b2f3554072bbefe79858e16b242c6e7f0cedd7aac21e1da060d2ebb6f68fd1e77da813;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c24dc40d5b4875a2ff66d55bf2f6befc7a881d51b1814f9abd19472cd408094b91528e8c24fe00501606603ded41ccb3de7d0f6b506c731eb7aa63f467b56b431a66e7ad5c7faa51cf48ee065ef0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb2144b42bf27af9b104ffeffcba4895de7b6d0f802323ff8e3c80c4521254ad2c756381312125d7cdc0aae4681f0ea07ab52e6de22405b9719f45bb6c2d5604ee76d4353164d8572fc34584414d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ac2db93650501be79773edeed673d8d04118cacbe0154c6cc4ba8869d5d063da737a11c8ddba1aeb6b0a5df62dcc01e219321ab723208f16e4f94637e1dbdf3f9caf071b71d3d094cf05365a7cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac2433b1160856c9cbba497c22828e26150ca24ea2e31bbc9230f41e1c83f6274a4d4f127695638e8dc7b8f496cc8d5018375b1efd3d45b2500f6b68c4d8e21fee6cd25ba1adcdb2f9c72be3331b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b00876192aef24ae689ada06a08188bfe26b212d0377986c81f4d6fcbed883abbc12bd6c258ac574dedc3826d6dceaf1a0c11c41561f3b967ce3fdef395c2d0b40179070efa0102b82933c452fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f8fe27095f511f765c589da7f989369177794c8fc47d0ada2a0198025da4e62e90c4f01aa53791fc63622cf39e419a3a8520cc7369eab82907d8239a0df01e5ec22ed9a35b16ca4277511986e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f2503b24ab2a49ad8af9085ece549872bb78cc665d08e6f5eaca1006d8a2280a96588f45e47e756916d2959f5b90a0f1c87339b0851b25e7233634bfb08fc8973e2b4bfc88974031b8c6481cf86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h73886949e646b27dd93189815c3fce23a3df5386c8799b999a71dc19baacd27090004c94abecff2a0060e8902791fedd07720b9d56844b0e356341235e3629da2d827969e6581fa23d74ce9ca632;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102eee9debba7a8ae77d5221a719820a5938a2e60410852a1bc09fb068bdf47c0f48ae3bb896fa16175f725d56836ecd8e0872d0a5e6663a40d23a1012a6557f9aa21d09a9954c16593d27d608b51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18df2c9cf158b2e37dd496a484d84b3177ddbaeab902f2bdf7b30f1d7030d52b935979a6113cca9e89a7872f58634f9ed38bf90d84ef3ed50ea8721dbe3928ad3046bc7e27424af7197c894cb993;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c06b33ac720faadde16f5f7ad48031e5e59d12fe9bab99ff2d9bc2d57ab0798d77376257ae48700d2ceb45940dfcd94bc111a55af0cbb0ea5fde594a458e84b5df317cfbf0a541c5b3d61a58cf92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1221c9313823809011670ba37c383cb822eef40407ed6480aaeb17929373b5e32126092ffdf2e7003002bbcfe137db38d9879ccbbfe26f8ff6ffe77529af64f7cbf517377d5b602cf732ed45fa436;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a600d99e03b0fe1d5bd588ea199cc6d33073c580e149a32c199ede14009c4a159dde087c12675f6dbbf778818a5f92cb91be2d7b2a8df9508f38c03f306f65015dd1605e09795aac6e8ce87c0ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93a1e9c5c843cf76439c6eb722916e41e29efe3a1c0907c0a74f1019c3329780c4244c52e745eb7c7b977ebd68f13b82f3c539d3aee594e36f1609c738d003dad3fba66f36749ef82eebde3d6bb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16039960348584d653bc22dec45bc8561fa1fd75b6fec6b89e2ab8a830885d2a0598f9d1e0ecbc1477efbdeb8bf1865555b5a0ce9925bc31315d26b4526e56a25cf00762f4cc0c3ff605c2fa327ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf3a370cc26d8195ac742a6ffd3bb15ced1f05bada9d71b112297655d938989848e6c86c71b68929efc2f4365d5909931ef124d1a5863d7b769d04d46402512fcc0c410ef79f687ee5f14f3e8846;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5dadf9814ecb44d967b54ab0fe9b1d401e6840389fcf2c6e050851e4ad5354182a1742be84a1b1e76b30027d7ac83407f904c2915d0825a5ef9c50f2a60d415b130ee2ded90267682c4079cf2aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4afad90c514e33507cf1096ee1119efedeb2f85454909d3b92558025513bad30cca0a08639dd274eb0173d819dab7e561fdac4b3d99c648ecf568b7e2eff5077b0514ec212e70de2b058a1b7faca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99208380275da08bb2a295d48c8534b9eebaab4c88d537794350ab25526b886ef45173033da680ad753ed27b3db6ce03b73f15490606e6724141be635583467c6b0e67606056472b47eb94e97e0b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ea84d3e846f8d76217230b21fedd392bac340505c84599a9f65b5ad45636068d86e7f98e87c2a3ff5873884df1494a7b65a529d843a2e954c94ebddb93b1f15f8d05d9d2b2bc25bc85eb50461db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180727fab129429b93badb924ce1492c059a0a09858e8d112a48b1405ff9b35b633f0c4c99c233ec0619efda77dab970b4b0eaae1fff64542dff0b8ee984b319e8b5820514b213f3a684502364848;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1685df04bf90b4015b4fc006e80f25f5467223b8a35a577e0c7c3d8948984e4047c48a1276d3b1fbab886a32ecc78798401df0a5fe3b591a7e0aa3661cb4187dbfaf9bb62337dfc4de58f4241643e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h923bf8b1d758915affddeeba240270033358f707d25eb634481f7363b5a2003508b5c23843fa57819638fbe07dffa36232eb20022543868d51828c05acf7c53951919fb98a6a6327d4928136ea3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf68477afe6df44c1923e96b4282630e210e7a98236a217c214a5246f575a160a535e218ec17b7e56278b903fb61c2d2a27694f2b97c28bba3bc95f44d3fb0ae4f7106818e011f205b71cb081498;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5fb41abc00eccdfcabb62ea3c0cac85ef842ca6d864024e8b6f4670e4451a294efc284af564b55569de2d4f3981ee35a0394f848270c6638c28d4082d50d12b0f20b4030cd2e2d34f139b1e29dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1919bf3a0610a1f14d92d50bd2f8d2ebbe152052779a6dd8994318c5f7d359d800d8aef508ffba563e38a28e53acd0a72e4f648767eb8d6e508feb551ce599e6a2d5e33c49607553e5f01b68b85;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc16b93abe5ad325b9a60f9201a7ee79735e7fd906bfbc38ba21895467c8340559147bd28df35667765c13f4b1130680787a312be22c5bdc669b58956fa1fc95228bf9200c939db61238f05d55e76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4430ca82c290c06f702bc800bcbe71dd8522ece1348c753610167e0e9c8506109c91986c05583aa5f706d853ccabd3691867a3f6275cced6ab42990241713a5f924a210ec0525e5d690e53ee667c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d9f900285d798afdb093a2d3628bf1fe77d056774ef87045c12ff26954bdf5428fc6d01fd6952924dffa4245c3268fc4c0240dca5928fd030e5dd246e73d3461949bdbabf74f6135117da1f85d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a735eb00d784b667f1e8ed621571f639a967b2206be223d2f9b1487d02baee9fc0dd18152deb55db6c60816eee40a131987ab4b2de38be3f96bd22fb767f0ccfa9610c4d3079e8074229256b59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16dba13e4db9db48610ce12143d34576a91b2317c05259a571075b4a1a180347ec7cf9e143b7f0776ecd8a259a7914f5dd0dcf526d10e675cea2703483ffc27c2cbf3a2763a1dde8c7f84e4a51538;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17aa0026a80638853e9602ea324275201d24b653b5d45dfe506dfcbc877e99580e49732d9063b1bd4ff7ff3a6c87d4a2313832dd7175c9ec6bd69b48acdcbbc61b753bb334f09be1c434e0c70afbd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7af8ffaa5ab74e438b29516fa722058364ac4d97cede6f8e5858a13d117f36e5722f75f47f8a962a9396b20d8f462023b5576d2e6810ffb2a22dee8ed0500f84e87c71b832edc4be65ed53e78e57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc147b77b288ba7f9c2a92d806f17862e47712a0525f6eb9f26a9467ce2e813c19257cb530dbd21d5d10c64c86d284308a1f56e42738a784cde3970bfba4a3c319e4f3847d97591c88aad601d6189;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb105d427b9987fcaf745fe496d0b1ec9a3a6cfcedd8d4484e6beb518786dd3111b1432307a0201b03cfc8136c526c36ff3b99f552534310c694879502643dd8fcbfded70e9bcd4220ea3ec287c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h675ff5664ca32098390e99a55b735b7f02a92c62f556eec34411dde24ea48cdcaa9ec8767fb5c6f16ca82ec27db281e823cb4fee66075c1f63b7e2a4e551850b8d04a12733dd4353fa3daaadb460;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcc220b77980078c3dd173b8ab6cfa2e6af6adf5f2705aba517d42f469b0be244ea471562dcf6595ef5f18a982702413a254493cee7ee7a39f98e52bb8c8af559fb29d381608a6ea0a1ab070b851;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d95137b7e1c2a4e1caff129d84792784a4363eeb71ca4b8f1d78ad7fd5e27d13fd8931171b6078d1a73e1a7c32599359cf29ffbf9cc95417b80f2e992ffca7272663ad5494c6548cb781cae1f5c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4e806f55aeaf48502002a3157ead30ca1adce138a2a6ef5b5c65d1b96c5009c61c691538ad63f7cfaf09bb9bd695248f09b275d52466550320f944ab69ea3ad3a155778e20e90d01337f2fbb931;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a1c7989addacf487c2997117a60853dbc369015d331fe982037851805617b56a152653a14fe7b0ade3535b3bf5346a6454dc8fb8cc81fea703b3f524604d5bdcbf0fecd8a46a20590a5634124e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb366adeed78fa7ea71988442cebc9549aecb31582578339913d3e49438006981899ca6dd17c3f3952d6b25349b607679c580df179f1068206ea2fdd72ca3d12ecb2e1152e57309e2d52d089879bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52daa6753ab28f2b59bd686513c1a9f5ca1d1580fb637381c20e8a7feb5b22b77a95686f563ef140e8028247ab341b14e9224f4b143b7968182d0f16cf75c047a159098389d60110285d5bc334d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haeb38314624bd2009051e51b7273de354318b870965b8bed0b872d30a90ace8f2a75043e34d0230b7365a4836fa196b3190bd50fc3ca144cfb19161a0c3a8e408288038adf34dd0a0b03f80ef24a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193e358d5bf096c0d62dae21772caf8f8d078f6676b0d7062499434df7e01c28b203ad7de2157e68808a92324520251a024b3e3422fcad21fa26e73413db0256cac72e221567410fc11b5023ee7a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9b03c900a38894aafc8786ff8df6292ac50dc2309430129baf61c37da56b231d43c33cba808aacad74f975ee67e9035cf7ad2602d0323ba23b241dbf5094d6a71424dc280add463f76e56059837;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd81ec98441136b33ee9914dbe0a976c84a48ea269f5672507bccef33b21a595e8a26cba219b36eb768650c6b6a682eabd76e7fbb12bb0f47f335a7a2f8cb5dfdb0f8227c62e9f43de2b32dc982f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca64f032ab0eb769b3ef9054489a1e6b01319f7e8efb31e2753547c385d7bea37abb8320cce1846e9108ad625b2504e46dc6947073ed768cc9e0c7e33cac0a7c807c57b97dc6ba3b481b5daf5695;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3e3f8b21ef1f4b5fdce0e1ca442a50805c2257f1e7ab8696f45aa409e8ea0724385cf916131ab950eff562e2e7c4159c5c8fa3e9b7326d7f4c43088bbc2648c3f5e8415f93764091cbd798b4b7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e27508db7a6ad6a6b54ff7760411d7bff990103aadb245b40eafaa0e843f5362ebfd046ff9efaf589f79eb18705920543220663f7de43d1818432a0db1a879a91b6f1d2d4e97e6fbaf9db2a7420;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef31086e5071471c6bc02c53cd8f87e5e79576c421fe4a449e161478787d5467dab1bd2b12b2f573145ec9c064eb5c6ae2ca105dc44ee3309288e13b71ab5390553d47654afad9c24cf3f57e3394;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdbd1ba9a7a3b4d971f49f8cfa1b58edbc285cb17438b7f21b9e29fb8125b1994167ec8b05842a5711008fe6c3837c19de3b18f5d3cdcf18661d7c50983ccc81034be52cf5a807ed60e5f8806f96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha193429e5a044038950b658742b7c5ef31e36243da7b5a77bbc9abde2889db1a19983cef73ad76ded05d0a9018fbad3959f315107258f980fbb1007ad09204a8e41195cdeceba7f122c0b3058647;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a9add7654e984b3e0a9b6a09476707d35d8d7bd7db3ed240af005d9fe4f563e39609ed58a9f9722cc83137a80e5fd8779088938c00b2a2735a1272e327756b37f9d7cc2a97adb4e40202d5c0770;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h660eb9951bcefb6e0ba45ef983fcee096b9814098ce381333a37b20edec15c926e4fc24560b83ab11af4a8e7bab8e4880db384df5a9ac24af103fdc0f89dda3fbc9dfd077405f0d526326a39ac01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1931327ee50e25aa61e561f248b78591c100d8dddabd727d9eabccc6bd684d9eeaf87de6766bc8d625952042800619ac7546ec4e20ca1a2a406ea0cb4144b3b3857e25195540fda9a18333e20ce6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ffe152a0b0c592860141335426cdadc40d4ece878adcab1c353489b48173d2d011a2d680aace30e16f25d4dc41e8f21b169c1fa83aef3782ed7bbee16de7374bc3e796503406aa12a8da9892642;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7128ad5fdc545986e8d5f815d6ba72d87c0b81e1bbc79e188da8add73d18b0a20390827465b01ef3daffe4d07970cd6bf3cec796f9e7f55ec6f576749408bec99917d1a6718713185581a918a25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9145887ddbec9ba7dfad2beb527f98cd8fb6726df17ab1d89f966623320c3f108ed533ae12caf9ee7cde7b6e128321e19853f658ccb360d64bc5a864b1f60ba50072781af582c7eef28f5e5871eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80bf313d596a6bdc07644d585e231b3b90f2d758b6ee1d2470a4442b9089c3c7cad97c04e7cffddfc882c67e289f1b5eb65542c502f3c3046464847636454146bd972be9d7709739cfd2e8cfb804;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8cb57e60933a21161d33bcd301fac64995e47d953b3ed7ba8c76c303aea6b69a678a53f6a04ad3f5928ffebb942841e211a5c35502ab37c5500afa4c40cd50ddaf9761cba99ec5083511496228f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef01c98fba6a6c16e176ea1540f957458518da51324aad7dd2754d9f86a537be1d1406412a146ede6036fac531a67a3c65bd5a8a9bcfff6737b5e67da39f58d6735532718443fd18bbee5b1cd67d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd29f18a68862ce59f9f19b6bc8509857b7941a160238502728043f8dd34b356d42f6ee403f1330d1c0e7336e432fafb16ffdcb9c09f4541bd85f82af182b7c145eb3b573c247b56a09eaaa7d900e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f5400ad2be4b2acd26b51e99e2e73d587f308d9a0b15adbc5d287562c28cd1cd8fc8345f186dccb3f55955f9e25bd2861d64c35598b0c6eff576735054081ac1f727c6e28b94d463f870ec8f418;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f07b2d47e76ab61c7447ad8d3f950b476441af25fb82fdf2025c1419a11e0dd79f29aa75eb2f2fe538fc83ce777427c431dfe4b4db308f7d8105bf8b4ed10dc9fed79df5d4f090f30af9352a03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1641ae6f7683d7f11bde7eee6f723e975a08d46c47d9f38572b53c0248089de1ae992cfe0b369538f84df279e0996d715eb300f592c4eafc91bbf5a390cd276b47f350f8629e2fb7e1871151aee9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0899a8f48d23b5441cadc36ea8bef7e0a30325922f2648b96ed7777f38637eec6ada22318e5b24f06662e01cc14f373500773250ad8c78c87ce1430ccede1247af419b1a7c96cee845b1321be15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h604b2cd3122acff21e506829387bcff794675910f8d3f51c994a6d1954d2b177c82e99dede0e9a56857c2978a2b1f6769d40a4313d4e46a4daca8c5a15d73707677b328d6d11d9e6a28f84edf2f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbfbf964c94155c875a5b82fc2c5920b32f5ab02019bd8b082499f93ec6d5ee06e32d69a987bf67408136c239c0c6affdd92905e0d66311df90c86083e5cf0386c42d86dfd981079399aa047647b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87deddcb3bd737780aeb35a24c37b34e91e0a8821e6caf87c3c0eedc3268d4cf8cc728a18aec2ca5f64c99446426dd470591570a0ff6914e178e342074164fb0de3a903f484e64e8143a4b891080;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf39c6069b5636b1a4bd48cce42346a5bebfe37ade1b4f911dc8d7b3f3919b5859c6dfc3491caaa6870cde42ee8ae5ad827a034e40627093db0a352f1289d3de5f93dd85c496a87d4210863c8829;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4605dd759070c70603cfb0b277c9a3da4429ccd9e300da08cc3ec88779f3a214348be7d6e59d93d311b0498ca0035b81bc2d580c252530eef423b72ea9fe550dc9cba9e6c31c7d8c754f379c59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbfe23c40a9a627c8840c80098ee4b46a352bcc5a104ea957a8c71c0035a1403e9255bb8bdf20a5fba2af9dff842023481e413067a2c37a4bcf501c15eff63172d033cd134634c77dc027855eb89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5cc78f50763d192b532f4ae29a02eb92947cdedcee8761640b8c8bbca3e1f5d33c81d0d1709b4a0e73a5d8c82b2c12815ab024b25abbce63dbb56425b2f93f203594ebab80b40e3fc5a554bc18de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1c036b2ac79dca8164921e8e58653530ca015f2022cb267442ead80bada2df764eb4e952b23365239a7f14b5e2fa548b6c7dc51be855a78464da4214d45f51d968e32b6e680cb21dea28beda7ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d8fb091c74a17ecf5259cb7c9e6d880f99e56ad9e916d592fd8ef1b74d23ab542ec7c91d6ed5f9c9e11fb15f1d55da15737d158b6ca2b129ff33fad1f6ed6a269908e80b8b2567283b33b7f9e58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb03119859174568fdb1288082298e71b53adb642277579330ff69c61d8ac86b94abafef83efcf5849d9299ecf44d2667464721dba01c60ddabea89e4c47673d6e27895f03a307cbb72934feb8ad0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19866458b1524ce3c24c07de467c775e76480c329589e4d5201044e0bce285ac1640dcd9dc83082e1322296b4c2e4003c94f1a0c80daf7371fab6a778d1e05e1fc760807629fdb0ff9e825a867fa5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1691115bd192a45293ad920dae005eb68360904bfdb11bd76c4c334759a68d951e6c44c1c26db0194e209d80daaabe619d8ffb9301576d4af15d590507c091b7c8746c8a3362ee4d0c7ba1b8e2c65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a51bc64f7e989a878baad462e7ac976cd21f624598992e5a0c688df7665c274575b4b22ddab7d4e70cb5304f35903dc05a464a2679a6097b4b4a4e896a6291057bd980d7b84e5dfb11c21fa49299;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de8db56bcc2bcdc8cc30ae4c6d238680fe65ffeafc5a4c709257d7292639dc9bd0ea7a1ccf0d8cc107cb268e5636edadca949228b80c0d186fd0dda3d5cbc5fc9a50912f8b2d589d6e3c10ca7994;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1945fa0d0f0efd7d5aab1fc7aad22a6e0890fbc177e69eb8726458b44aeff70de35cdb6341623aee65b351611f49f77f74683c9d0d145ddf887eeec25bcac5d9299c531574dcb15b0009f7bb184f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hceda8cd715e8245b1148f8c846361b9c8c59dc74a7385b30bfc549744f96a91f977882260e3f406427a39566b5eab9fb652aeddb718ff0d234c04040d6e46be569159ab65402b57d76f694be90c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce91f132206f66ec01353aa31ba1b7eb7912fb752ad79d97eddd4185df95f3bb763d274d95f954d9679254b68a4b3d6f3e04a940635b324231036e7a0eec37b20e536451e3baf5972b6ff8d4752b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91331e1718efed7b0f2c386822794f62c02287c5219e98edbc4dbc44604b7c0195d958a5437fb814a19cf569e501ebfd24c87ff59b9399687131ce17c81b97410a5eef7220862d061ff057643f2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc17b2c182a361c224cb5f144509d85c80901f17d5f4b032386fd81dee29f5532f841896d2e212f8a444b9f5091553347a8ef3de56d712455250bf141dacf9d0185e09b700994e8fcf72a8ad5ce7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf0585b4861fe1b4488b40e77a162a798097a64b653165b2199ee8efefbba16d42d0e05cb1e2cf5627debd62e4d2e515c17802c2785ae15c05e9c5776a5c26ec3a463926cb1751613f8eb5feca51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c112950e5c9ea1a81578a65770d9ee360186d27384fe133ba7b1010ea2c232f50d65bd2a8276bcda7df4593b4c5f67840ee656ac914b39227e710f95473fe55ba9d0cb86469dd72e001f44d9e3ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117dbd0ba3261f150a81ab22bccf5ebaa672704171e6fcbea57e459e563638b71070bbd3748fd179cee85b7bd9f1a8005a2a5a29fd05742b07fdc997156cbdf3863ecfa089f30f85f922f223a6cca;
        #1
        $finish();
    end
endmodule
