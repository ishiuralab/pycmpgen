module testbench();
    reg [28:0] src0;
    reg [28:0] src1;
    reg [28:0] src2;
    reg [28:0] src3;
    reg [28:0] src4;
    reg [28:0] src5;
    reg [28:0] src6;
    reg [28:0] src7;
    reg [28:0] src8;
    reg [28:0] src9;
    reg [28:0] src10;
    reg [28:0] src11;
    reg [28:0] src12;
    reg [28:0] src13;
    reg [28:0] src14;
    reg [28:0] src15;
    reg [28:0] src16;
    reg [28:0] src17;
    reg [28:0] src18;
    reg [28:0] src19;
    reg [28:0] src20;
    reg [28:0] src21;
    reg [28:0] src22;
    reg [28:0] src23;
    reg [28:0] src24;
    reg [28:0] src25;
    reg [28:0] src26;
    reg [28:0] src27;
    reg [28:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce73c9057cc4fb6a4785e3b2c2afb30dd1d6da993ef8f9442e5a0bdffda7e832dacb99f0532850a1776e4b623d25d25ca9dde7265f01173ac92073faf759cb31164d80a2c12877dd1bc300ecc8d604968f2cab7a513f63ba31cd006df403d7891cd6e91c0c200972ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b7e62a015821318ee6c250ab2e246a9f117843a223d626c90c35498ebdc378688a63f902558234840e89bf964ef7b510aa7ef696eca6b2be392fbde27ad33e5d0767dad919476554d2e3e7a9274facbe8f8751a493c58e6cce0c7a8bd10a94d5c38de8aa346d768e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1668e1cf3f8a69d917614a7bf9aebaf45462dcd1109d78cb2102928821f67520516ad1953a9300dcf78840120341c169573f4fd6a5af98cacf2f3f6da3b6aadfe3b1ffc29cb7e7cf36f536830f5b91faf8d85ef0e81d9ef4da8ed28f4c6b5a27aad5c4553cb41ee8946;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f926c2b47c7bb4533bfa7681a6faaf5a7e6dcef3a56389b2ce61ab688f4769ef84d336afc7906aa03dad7b6637e3fce16af3ba4380ca7fd27849f6fd64c934ce5b0985be8e8390531b2c1934e08a1cea515b39120dfed7eeee118d9f1be504e878ec6e2769e66b08ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd8af72dee46c52a92b815427b9f39e73bf1dc45dd39cdeec5c5e9a8e8d2dc894018ccb7cd02b6abb464671a82152d7ce40c8d00d2b59a6fc249105649b2b1668ec2522baea11549993b933c1fd0c139eaaa0fe60e07c8a2fa33b53c56be1a8dc3dd85528090a4ad14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11564f2c29c4e00c3fd7f3b745d27974da83a856a4d438f8c2221b7958df10c0adef261fd87f022b71f2050326e8c2e8fcaface745186b356518ce826c71c4ff8fd88f9bf215bebf591dcbf4c4f32b19892df19904e49e19936caf17367e1f1c1e7e9a2c9586e7706aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15830f18920a0e71e1fa2361b92408ecda3c3bb142f8a67c7ea393b640e70f6f02d93b980e36daf975624c2488359d0b510de9ebecb6f2147a60ddd771284391430a168defcf92e15fbd3b564e742bef7827045f82ccb94dc965c00cba9bf8a2af0ea11fd05740c1159;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cde19aff74fe288779f2c203c51b9850f80e5ebf237d363073d466fc9916b8c266f9b7d7cb81dc635e5e0e9d67ac1583d0e865cc8b14a55105a95c9c295a855905e8ca187a33da39d4f42bd561470ec96de4050b4ff8feb61ce01bb32a59047ec31ed8e846ba401d1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138d11d61758f1effb6c746cebfc18a787dfdd81cdfb75141cc8bc5bcfb93f09fb522cf9010b7a6b018e70370a533d5d803fd4c3896ce8e59dd17b85957a98527c378a90a5f9cef76eab3c2c099ef1d7ff5c4fba07244fd014ebdc2ba735d2c89e7af1b281524d2ce3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5879bfde9ff7b9c02322546ee8a4593c85ff31729f89978f1984518b9521b0ad71bf7f6daadd7562e766701f2254cab1676820df04fc7481536f4085d323b4df86996ce3043a1271f302d08ca907798904e97d75918964c9788e33573cac9a3611eaa747fe0cba68ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1872ad90e9cf5f6217377b5252e25a19b6f239eba92bc640524d4878e5f0e74444e0a97c67b8ce2aa0a751aedf5640beccd71bbeef3221a524bd3b2d87918abe3819e56f7742fa86433e9d3c3e7b3187da05069703a35c9dd68a26f2df80ac4d7e8255d8b8298e01101;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba36bcc6959922818d422b206033c43600d917d6a0c001d88f1a74a52f946adb5dcf1dbc8a2c497df62ca7bd5cea2f9940b0ebf195d392fdab832d4b7eefd1d23cb7d0737478d9a5fb829c5f33a84d1366c83a933571b53437bb2a7552214be5709c8486a33b4d7f40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f33383cbbd27520d0f7a967c01127e84b62bcc81e594ead0f4595a97de21440fc7195a680690012c00686ffc9c888c41eb87e90dab64b8d3cc44e577e3b1a4a1ec610ec316fa6997352eeb9b6117f99648f2ae925bec56fdb5237edcd104456730e7915d914aea0d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfcfeefaab246b0e46c37ff770b961026bf5af5785a4a7fd1709be91447f05e5b816e037eeb5be95d64ed3fcc36bbf488ebc7c349b0fff6290f39dd418629ece2add22480c963e5c166f488048a2c65400a95b0da56b4efc4a68d3745ac79477f4d0c842a202447e523;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108d0de0d394ca0b71af92f1592b2b3f3ae5bab8169ff5a0d493c1540dc2bebb47326424174a2b1af5138143a4312e003510aa3835574595e99134da97f8ee9e58811cd10ea6a4ccadb5d2518a22afaf1b411bc5242fbc640ea6e86cbe78af43430d8412fd288e91e75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5eabd0ee21e5778c6c4e0c4082eec5fe2bdecd4e5a66f6862116ca574028c4b4dc9ef095a789734a40accbdd58e05dde2d9fb305c029df0bb72515c6f403ce45cde26984e344d03130d71c866c35acd8395408ddcfc6c2243191649003ae7d1ed08b421fd16e018a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19646d9fdb64cf62973b7e2fc074cafee913b141e11efdbbd6636d8d049125cad6b93949e23ee0b95da6bc8c3958b7d9a15ed0aeb72bbf679b605920270a8c61668adc9809d7b314afd06769f87d3a54135b44f2f4f18f9c39de5bae491c981e6433b2ca427f8a5e9fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21fa3e3ed34a61319e7b467d8f1d53a8b33ba686642fcc655b54abcd8c563148886d809eb76ba5431f1d382ccd7597aecb4c1ce0df179a1979418e018301cf8a3b417ac30b1ec1c8cee5769f3858448d4be823b3a05adcf2e60f2438fa2b557484a92b54d0a66ddbb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176a12a51554b2a6e0dc942f0c390e6544e35d4b647d8e4219bc67fc4a833c832d544bafa600ece75c0c6ac92088a752fc005e2c1faa8dc4b2d9b0e5b913335f255b4ca3d867a31cc689ffc6f44d04bf3e49d43dd2a6d546d91561bcd8b1933480474cabe7acf907df1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173882433c5e9c7e4810c8bd649e145b53cdd5e7b679b04ff26474363eeb31e5983cba7fe659019fba12482047cb0ee933ac8666548507569eef658b891ff692a4f51378885f93e8e83f4e717571b401970ad61639b596e11ab407c12b04f5b9fdc899e926f45f3eb64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18449977b82a20a31c7ffd53f04fe088ced363c11987de3ddd1da4452bf28029253fd540f08cdb9b82aa1fb9650da4ce3829f330444d21ed34e9e8f3527780d7cfbe8261afcecba44b747a948b25ebd538dd12d7d408b33b09df4253e47e00ce8babee9912a3fc9f36d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1e0b085fc06cbe92a1344ca271e7d48884ee54cf1840810d08af371b839a06e50ee098e0716f3eb7e1ffdc028267d7c0bf110f89d3e0eb725c2bed5efbff5c085d912906bf1e900319bb611cfd33993653a54a86e904970539adcb70ad55a43614c3bb7e830fd697d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be9d5273e12bd4f7fd8631f1a5a6b4b9e8c00e9bed3613bf50cf20e38a2c6b4bb82212bbeb0e9f52fa5e149d4f353a3c2cc5e2d97315471c0c23bce383c10da4ee7301a4952dbc595a65f5157afe5ca9b4d349462e028a70e67197c5a0a155028da3ad83976261485f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d43e9c249d890c0430a61d6c3b4a0efb175c2b08a1b2ce2e9494660fd7b8b52ac09599246c021850580280e966eec3f70bf966cc9ee480b4e832ea366b444fb7d86763550be5619ae2f6865239f45326afaed3711b5c4a6090302e3653c10d13a70e61aad035fb312;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b3ddff8a7ed16f74d57900625b78693f2e8d741eede335c0016c26b0250c9363160713609c3943cacbbdba7e84efd4b65981e26a6de8d836cd92434f9312c61ece41742ed0fe7e129434878d619b34168479d6f91c10383bd2fe79c31bacf2f639292dcebe697f984;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70f8bd307c46b193c951915860ed643050ed37d946dd9faa521bc676be97620f93117a031524d608a2632c71a2f2085ed0df2ebc3960381471f8e9018d94be44f77ecdd821a137da0e6ec66aa5ed52a352b4f33c88a2f0c453b35f2771d7a319da6b66297eccc14279;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1b85f1ccf9ecc186759355ab6dd9c7285ec7ca5fc63916c7e38ec2ed2ebccd8e7a65e406d7ac1b9a13593f7c019e958770ef62bffe12c43c8324edd8599ff0eba2a5954924a9d565905a36192b3ab918b6b026ae4ae63093fc1291ae2d5c48033e7631769e8ac9fbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fcdaa2ffe9d6f6f5e35b58987f2c5193db5eb5cd446caa55eb906731c09bd0349989f442378c1c7feddd34920186143266f49bf9cede0608ae842debeef1c43edb66ad77718691db3194388744112f31535c20d229bd3a770920e5972df711e64fab2d8dcecd458e25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb6df2888fb2c2fc5f0e5fb011d794418eff3ade75c12901950920b0a0a90c5430adab26a410cfc84bb17b9d9fafac9c5c1e7fc4242cebff902be5485aa0aae4821afb2174f60b8ff5738ee9c52f96ffd843f03fabb1014e88cb6d2e7b67af21c2891e504287d3fc85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1486775b1c6f4ea1b7ca97e3b7ff761dcedbf86e542979fe49188645be4d4b84044789dc513f02883c20a7c8e8287b21de3a48bef9b271069584f911f00a04fa0e925003b731c5e930db2f6ddfa704f57b5ec0c4b30df155bf9f5b47ffefed8c2cb1c6bfc5e9b380759;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d514d4537aabc00491d14d9a0c3226fa6a0f68b6d6887152b37780ee0dc3f4a865699343d491d1987bdca5c303f5a49a55b1842853f2ea541956cd8fa52972ca03ee81afbab296f5d3976eb677da0b2c42abe6e47b85afe7b71f5d1132a7aa88b67f2d3b21b82ba4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aca11bf19b1f5d6111da78c28ef17296ad20bbdeff5b5c0cf179cc7cf89e02af4db4ec9533f0f6d0b3d3e1d33321b2771f01bc07def28648ed081af3731635a01f5cd76e18010d573e83ded808410c566e96552b33470a79ce05bd9f19db7b99f314e016bd59030c06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee352026738a23ade55646d968ed91a69559a988edcda3cdaeb8481a440855e690c916c79743218ba9d285e139b3e9e2024e87dab0c392fb6fd219949774d679d0e74c9d73edade6e40042b6b145c3271eed4018aabc94e1b429bb434c5ab1c6e8a1edfdf7c3785e0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hade626ef81dc0f829dddbdda6c6e9f427b1d3a876c6b82ef10e9909212fee247bfd119708df1f66e8df93c983128abb9030fd54e5fe933b85230f325bb0f3e21122ed92f5a2ae3c1e7f73f38fd94d2e9f8d8d49e23188517965f82bea0b0a4c38314ab9b1ad0fdb598;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfe7f050a6073ba779884b298c3f0337f298a0fad6837a65fa1a1cadb18630ba2533b5ca9ecc71cba71c530d4abb7c1f1192b91411219add1c30de1f29fad667d59f20c5b545afc26139c3b9c50f9d8294f1adde10de4ace856ba1297b81696fdc0d7bfe33227d988d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da372d5abc51b04eb30fb9115f90d6f3ae0641497d54e4e631c3be4521f83d91bfc7aadab0009bb3e747342f842c4262323629c63b59837ffe87ee16b97cf6086b3a9184701b6e44fa1cb47667cfa74424aa58cd7ea566fd463aa9dce2fd658a1362c0678b5bf8ea56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42b9bfb9b93a3085ec4555974e8dc3293193885f1827ee7004d0edcccca1e551e812e5ccefb346f22b656cd2a415f405552be4e1b3c96252881ce3bd4359bd37c9dfc7324a65530aff3e6511ea49fe9833065fe68437fdb55aa7ebb8358fc2fcad5a725440495fee58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39b05a0ac5928158d8731b81a7cba0175b7e2d74896ae3d25490b51453ef0ef558ec06fc2390d267369aad46b7bab27b7d1842512cde9a8e798ea2fc1a4b2aeb3b3ffa6b9852fcdcdb1412ac13942efedb199d1ed35c54ecf7ecda75ef424b700225571d70d10f1dda;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134e3a3ef57ff692c8565a4ec0cf36ec25bbd23e18bea48a586df66568865b4ebbf9d6694a5aa8277b30b51d59ce4ad366001331fa22fff76c080a18a227a9c45f5ec364b457b7d93e24b81db1f25547fa92db996490a3c9df323f8b2ad86beac2f94ac9a368bf527d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ec241d98bf8b64c851bc8c07468a6cd2cce5db06479efc96255ed27f75f9558808c5d2a776e31557b7cb489c77fdd13dea536db4710ae77bd462e6cbdbef660171cf581bcf0fe0953bf8b07abf69ced25538d50eee0d3c6418454022b94b95d0b7b3eb57bf29dacb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4333390a184b10564de1ff065001dd7cb19a3feca4f8dd15a0c138ef5b1fe0c17a9ced84a45c30abebf2d7ec0bd8da4c36fd2872426c94e13c8bcf705966797553da52067abd5c2f10615322d81c4472f9e40e58a9a06fb257e00b082c8b6baef9cf66d96a7879554c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f15b371e868e897f9082d07d5ce0c320a8b81cbb58392a0b2df230744152c532f54f9be1d5df6bd0e2d376fea77a31e62b793ef47189a8bf7c21a57813f162340447717eb1b4c0d7d9eadc9bf8aa0d116935b4e79eb1917719d00891de13747f442ea66f579a00382d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a744400632ee569e9bdb6653349b032d1dab9ba056e0b330b41852794747b820e2865d8bcac0ae0ff72deaae73f1d13f3577368a6c6014ad15affa6b98ee417fbadaedc7065feba60eb5de8e748726d5cbb3bdf94407d5f11efc5a676f3a70be522109e39fdd035e19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14984054936121691e668fa577db9ef88d59890e0b65e9735b0e941e6ff837652bbe9485198503f2f4d2d4947f263765d3ca5593657b022bc15efec718af9fa6583aedfbdad997aeb8d03032a3cb038cf6dd97e7216890dc51bdb56300f71316d24d0af361a4c03137c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ea7ae7a0d80018306936146e61e4073796d63f7c86e64f49bf79c9b0ab1f30fbd483a5f8816abac204263047dffdab10c994b8d78e0773fe3237f16ed92e6a6e4e3015fa98508bad49639603b425c8c1e2a11c75d574c55dbd3f67623823dafe79e611e0b25109158;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19076478a44467c149e314961f4ae09c3d1ebf99673d41d8a6e43b53da7d7409ae30f7a3ba0ad8d928523064af03d6a8c025d798ba724c0935e3bd2be6d55f7d22ed01b552c7363a01950415d4c6009f59a38c84e44e43efd592c7e7baa64e2dfd1c3b9f8d5fee9c24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15413c20358c6189583e7693dcfbeec025aa4ef38a46cb3d1f6b8457a7e407ab19e2c169f4267856a381652b27e2b6d811d8fab07db62139914204c503568d70e1adc13ee3f862306a96d632f3e6024d6cf5b674d8013a31325e936534f70187150eea838d4b2686a1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2afa80f77e3766e78e32f570921d8971359a2a132d4192da92c93095f3023e520ee46299f74da5b7b6fd4ff0e065f318ca656f750ee9a22db394634b212e975a1c77654fc8ffb042af34d96e7d272c595b7a1aa8d9a7448d085c6f073706fc94a4f43362705ffcf88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0cfb5920d2b86886be57be24eca179a3a34f974e5deb2145e05d05ca93ba5811030acaf664f63add52cb826c9f2346d96ae2a95a5e3cfed4df3c34146c46ced188cf608d9043bfd5dbcdf7ac083b24a40152c1ed0d7df04e8b3c8a2e2bbb3454a064a9e9e798538db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he0cd095f96c9965d3768ffaf19825381881df004ec94b6b107e0649e4d74a4cd716a0826c14cb0a28b20df4f2048f6b4f808a881bfe01f505a56162d70c5dbf9b6a50935e62a2460b34567dd8995cd7440f09421c6c34a282f86988383f148fbf7f0792f026e05adf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e5090b6021a2bdc10c51427c9b9157ec88665004cde2467d02c48455d62e490c624cbd0bf801812eb47dc52497bd5ce55859045716e8255ed7b36e7cfb0fe2fe7b7b1d6e9fcbb6b4f5052574dcd904c1605791b2b01c0c6d1a07fa24352afcaba932ff12f5d14a371;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ad20169fd94098b3a8bc78189e64f6b3f60e048ff551a54ddaa05295e8dec5d54b02b8c21c2639ca4ebc1db4a2999657286b54c37932f8bd552e37a1d725679fdf064291200e0d61696b32c251c4e4e6162aa3ac2c884c317c15a604c8edfde13fdc79927e9d022b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c03c0f5d98161aa0298c6e88a4e15aa4795f4164ebcf9f42cbf7f97b1a8d208b2abd9bdeb2b254b3295ffd5c23cc78c77a83f9bdc1f6caa755bad0a2f098c48d9d85d8aee0a96d1933d78b2a00ebbf7fb9d4cc0db09ff1575bb29ec141e9089ce34b0a2e91a96b8109;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eab74e69b3da7f349bf2db15c29f12921368f0afc84fe5a36f1e7b89872fe9c96419c2956b635e1e7a1f613d499ced2f4f974cb118cc1babd12749f6310c1e29a6ed5c78db71a82c398b096ad20a8e1b3a48670a80cffb2ddfd981755644723ccc471c397d37cf3e18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d4dc208a2b2f193b8e28bb08217c87bd660f792bab971cb768036dc84ab7f003e6b9b76516b34b9f5539664e9fcc116a6476fe15576a16786d5b634b5d6bdbe4f38db21918ce41dc10b664e878b557b4b35fa81f06224723ebd2beb2ac7746108fc9ec9d14aeadd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9d345b31b6fbb19b85fb8d72635186d1568b6146c4c6f5eac923ab57b8d46ef8f64dafe563c60785f4289fadea30fa00006fb92d7db338030a9dcda523d071580337f5ce02e272b8a9f09b6012f5f1bdc7bf56c5189aa709ff594418a668ca8b0f4661efa857a5f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h612abf0df30e42dc1303a90add98a801b3148f3a047d786907d7e2240f65e111d4c1a7c24bb975696d814be9a10756522942aa4f6aa73c19c74f3c8d6855b907abb93ca8c3bab9e5ba057466b8665f4e84f714d255f811ae8296f47a069f4f81e6d9f41aed84f0240b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1c3210d00b4a6a0f862b1db677d7087d6dd805f158cd87a6ca81ce763f96383cbf79b0a7ff1da63f5947d55ac9183a6fd9669a5045a6f66c38fd9ef4ef5b47035f46c17dac696a69e796bdc37953638fe257edfba2c1a1e9e90ded742e893f849dbae3828f6f8d869;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd950014df348e36000436b5b136a9b20567c6ff3a3c5134ebad7574f1ba37eb7c680d11c92f85bacd1b750878c8a38938995a5f9061c6dae52fe4ae8da42c3203099174d9534acbe7d8041f9e543409017311a2d3bc3b28da0ef39d3a8f5634d0c620c3ad001ea3e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd267ee7405ecc59036d97692bd3b956ce9a4ad23e9f30b8cb0951fbc683aab8b91679a98c0a7aa2c44f7ceb8cfdb43f3bd0ab967cccea2a5417d0101efb92e9e2d9215b4345c30ce0ba701462b356ec807822b274ab32a570debc51dffd7200acb6fdeb7915f26c356;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a147e12c22d67b044f95f8f2f1e4ea55887be67d5a8e74c46babe66ec3c73e1f850382bb92c447c4821e360b1499f527d22bc3515768688413eed7b14ed3f9af8c68cf4788f4e15ca2dc384c24584369e7abe850a908eda795e2937698ecad8bba8775c3990802139;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d827c25fbe803f0f6663422e9e2dd22b075d583e79cec0c39ffc201a46186fcdf5ab1f5e27e28a09ff97acd0f7c9011b836609006ad95df50b3deae199e14e5c3605d9489b321c7d01ccfa8462ce571cb883d4fa97455364dc7acdd741f42d42d31492289bc3019c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187077be23b3cdcf6a731582228a49de85ecb4bfdf5bab39b8f7c38eda7e192cae59890a675e055a1c1d40fe09a901cfdc7bd948672e70474198e74ea383e7c1ddb92d03f04356015306a6ebda938dcd8f1c2ad71e27db50c6165613ca277629c6874e12496359af74a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c1df3c237ba018c58b57fcc50e56b735a30eeaa010964b967c01291f67823d81dad5ee0b87089e401d52cc17561d1d4756e44cfd8a892b33bf638cc884ab58b32a86bebde82d4d3a87e8d27505cd1b8457122934f3d03bab5d72e4086122d8f501a7c3c9eb8824cf2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c6067401c3e7d80bbf66a7d27a7bbacd70eea387f7de943594d997ddc6961627dedca192aa42c04d59b92aea8ea8f4ef34e89bf89f191a3df4dace170ecb88253f3d9a679e0cf641fff7287bdd28b3274d92933fb5f8ffc81774cae156177e946bc1423891a8a8dd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7df7e216a2525d05ea599267a51d8e73b5737d296dc688ab63849c8c198905cd5674fde77d8e388d588f8db4877df08407860bacea0921e54bc5009c67a2826db97e7b7d02e1191e9e58c22f4450b6c4ff1f2badeb17f7d4230246700ffbe3c46006ad28ccf4bfe7fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b49792e06f2a468c8f9427ea95181407c7fcc40428e45ddd3a385308f4e05e10cabe2c9926176a5465475543449647d12c1bfbd5b5bfdb5c82d60956f260e5273e87c89c024fd0f7681391e5b834f621b80d1d8883d3a3c90cb95e922f8eb6a4adbe6613c4826932a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1caf14d6f8ab1d6fa77e33c711c3b6ef306595ff1c6c9b7ec8fd9dd419635d907b1118213784fa6038a496baefe3fad01bb99f9de30c34fec8c94f55fa474c469c20bb7f0129e924ad36c9cf1bc737b6f4af1ce4d85252d83f8769a0c55cbc2436e0fa24e5a2e68bddd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dd3516348a9ed48d6d386528c0b4f24486a5a80e53653eaeaf84844e0130f0f3a1c373d2f1cbc43a0c454ab474dcfb22f0ca02f7165e38c6d1f4d8da1fa3dff18607b088d23696911c2cf7f0aeca748499ba8aeceb21d6842596d189444dd5566143216c89894fb6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8dbd8f34643640e2d23fe1c0dc74104fe60adb3266d2a711021a00f46f35e16731fe84c843ffa424e101db2498f4b1775f9b86df728d2099d6b86e03c1d0bed89614392e2ce009ae5bea57effe3fb6228a7e13c98d01aba08109d1190b65bc8157ada15a64b0c019d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164a6081bf858074893fc82f27fe817d7c729a6768773a87def87d3287ca3a4db217ce338c4d54317a23c035093ff7d39b14c5aec1a19bf3214db72a59bad782037bd78c6b21bc1efc44d0d6bfc6af416c21417341243adb0b03c4e3a75f7667724afcf832a4f3aa2bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c3ab1c5da6b0cc361bddb70e458b8ecd6d84928749935808c805ba2847fc8cf520a4f3784c2c6c2f97fc5a1944b507c1c6831deb3d850838afb5496bcbe257fd56cb50b46391dbd0a9a9ca03374c205b36fbaf16a7a70930d5db778ac42ffb0fe005b93f49efb3a32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188dbe010fae1beede221dbe796c391e2f38bc5d3411f452ed71a438079bfe984a463d19fdc9740457c853faef64be5353364b2ffeb9824763d50081ecd241f33ae64a6c209a7000f6d1ac982b57d818174fa3744a5d9c85da79c54ed929ba0929c1aeb29cbae6322f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a016ceefa5aa9300f329c73e16e2f8fc9815ab6d0d2ae21ee8a45943176f47c8ad458f9a83fb67384df7ed386cb9c3afbdfa5c709989975fa66ffad218533b2ad47e37c2611e058eb9ef2e0dc8e1f74ff2fa511e14f4c2e202a2a75a62395bb522a76ba3e867f9b120;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1486ca6caf5d0c9cff970b3f62905a09c2382d27ffe8fe9f17b39b6a18257edc21fb5e277973b800e9711a9dd6e549f6ce6da80cc790fb8077099a2242c19913e8bbb36417fac142e6df4d927dfa2ffce97dbe87ca50539fac0226cc050f88584627f088693ef27c55c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1edc10a4f6b38249721544b5d9cbfedc8013e5322951f7acce19867b58b6b873d92406343ecb5362d61f82b6607c1aacfb446196e0b050e37c360fa6acb7e6bf35b0d31ced2667d2da297bb525515a6645ca8184d11b42f9265d0741f5f88c096095a4a25c8d40bdd5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b927f052d9c0aa5e6be3e4dd80a6768431ca36058fee41e9a157c15469573f5d2bff8fad819b02ede0e61973b2c47b32b32cf94acf9e40885b23d44444f76356433cdd04a73c963b183e1ae80129bed2cff516705fef81002a37725936f3b775ad0db888a75feb19cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a063fbb7387d22de4abeee5bdb99c05b835dcf263b13c3b601b94b7f0da8fee51b8e561064b1697e2f1f1b0ba7af34c9705456969602670e13eb4ea9bb292c74511a1f7355c7c88c7647a1a6b49d23ec36cfd74fa07691cdead3379a769973f111ee208539753f919c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha888b3af01e9316071707cea5a41a1e079d963e37bba65ef17771d0e5819cc161bc0cc4185e074e1eecb8d2bf41fb0d45cb108ad47dd68ac1dda6d7139befb1a5bc14b916f0c54d2a379b3b4315cc36458e4447b02adf1d97f65be43b6f2cef4551fecf181771c13d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f94e3774198bb16ef72a386529a9924219573ccd7c1796bd928b9082c84f11bc36b1699b5619903cd6639452aaef65b41c95ba00208cc3ce6507aaba58f025ceac3e1dcfd1d00e536ed9a81f8f633d967919db4a916fde61f74aa7c61fca2a67b23361312c863157b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fc048b91b7e32870b6786167eed84a9c0c2cd0b2beed01aa6f40bb2692d3ab845974d086ee1ce99051b79967efeb9406dfa36378528d6bc120f6afd1c6463e610c083641f8f15899149595d1d62b65d862bde558657f8b77e7fb5bb26a6318e284510bb0f9a79ea59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1d9c4930902340dfb9eed95dd68723799f2f107bb289630210c1b0e8bde87ebd4833180abfc36a5782a0b2a4af9808ffa6f1ec762f43260f90d9872396753a028dbc151ee59b9fc3d5de68cd081068069c5921c04f133f691c3647f0ac78159526b509bbd2f5314ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d10a648debcb9863239bf160d272aac31b5c3eae49f1ff8b217da77fb69b8cb179327654043c4a9c396877346054af6bc66b100f7d5a6f862d2fd7ea4c4acf46a6aaf8962c1ac98c4a823c6fb769f142a6dfb6190f218e6a8c8a5e975670994ea699e523578bc27c84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7dcc1870d3fdd6ad3da439d2dde4e909ca3f64d50a5be0eb67701965862d102d79c4e2748d30e758c21f9e46fa1f6b42fab1e3984d70ae2bbc41db67a788378c4e945461d3a9578235f48e73e47a8af50928fc5416ecb6497a121d966cfc358b2286e31724cf697cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10821b6b73a8758c83f4e7dc8a609e9bdfce4ffb4e5ee9b6c2fa1c57bca808307cb25ac38636a9be7a05c80f3995eeaaec0c1231ef2130fea1397b138918bd1373b8131b7b708abef5cef4c8583938be7526f4267783c8b8c66e34b64baa9e7eb970c08c1df6e518d10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74c0b026d7783593ddd8934aa7c40cd761b72ad4d85b2a7299a031898ae1c1d760cbc325594bc858204546be26ae182a68a5a099d3cadb583a9aac42f534d55fb10cee6ab25b5cfa75aa247716dc0bfb0d63b1f79acdc3eb13698860455b7632afcbd8a84fc75aef25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d9bf1db3365d8308ce635a5a82b7c3650cc0e5b3f773f9c02b15ad8661e456390ca29667c5da833146cbaa3109b4745dc979ec7b113315d07822cbbe2473b21f5cc5bb59cdc5cc96a15bb3c15607522b2e1fd3a5e4d7e5d61f26f2232101856fb7b55dce0a432f1a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1604800e87ee4916f676e96f6c28be2f8040b27fa2f80a880b4cf3897179617830eaf5a2209894b8c4892c2fe17776c2aa211c5219ff02987a32cc2af441a1e6ee3e818ad7dd4617c3e6d2f1e69adc8eb9274a834d897483e3f8a5aeff65c7ab478b1baf513e239f52f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b80a4a4d802d8396a0d35d80e1eb3fd98c71a862ef9f113d9c8a0e6f65b063567647b7be9fe038440756a97304c621f92ca18f7586a06d8a62b7dec7aafbfc9e0af10437e2b4fe70739c4854d4c43ce78f585bdedd9422c52a88420ac89ba7abd54606c8c778605d76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43af5aa4e49029638e42ec50a7a58261b77408f9d49287dd03c593c56d38231ef4728452c06e8c285c6eca92769ecfed0fc4a91cd2e222630809ad274329a17291aa2413bbe54332a43d52660557547ecc8278472a17d0b5df9764d14d5000c68d877aa25bed2ade4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7438206037fc9ad81998db19150c8b8edf0b3b3b9f066bc49bb1e8ab4343e8c2a31795a3cf6cb45de4d5576328f47e6dedd629175f96799719238e67bc857c37c8ad47ab3949e882731181b16fc6be98f6abaad7e966d9e5bbfe6011a1f5073c9de64455b098c74c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff59cd41dd9abcbc9bae1024423d68792e20427af733f9afc32e163ff3336ed4c5093745384b9e5f688199db90a7ebe11dc59529de985195b38a4c8242fd9a2075dee30d3f5a6ed9061feec90dfb7677d423449db887c9bccfd4faf7f22726f4e2a68ce2113edd28ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b792147b63e5a576d9212563b6a69aeb49e4aba966f5d666be4d5036dad4eda56401a0de9e5909b9a955d88618bc0ceb59512aad84546b0963004fa86699df915efd0f9a11d5ad43908b7151f54ac0d2b5cb1edbd3b09614097406e13f0dd10254e575cc85bc1189e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he43847d157593b6c341a9e742da9fac61d279063d2dbc0dcb85c3520430dfe1a54ef7e25eb3d7b81ee985b2466f8556c721b164c6ee8d3cd069500e3029e63c9585c7e5907ede0dad6395e7d733b46ceaf62f2f51e4a3926a30ccf823ebfa8745844487c17987be874;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162a2551cfbe72f400dca7e3bee2e4a361ffa0567fb32c4d359aa43fe566fedb893414cd00b7d99f277b4a1fd8640322915b803e986142baed0af793a8abdec01e4e142d982346751db625a856150fdf0c33c8ae6da87fc222675103056b320e90e4cc671e04cddfb3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h301e65d33f11ba61c69ad8c1831667e2474f62bdd436bfefa68aabaab12d4f4eb45ad1529974302a6fd5c701aef165d753325a2adb3b4232b5f5585e315362d5a461600e80e13ed1a638005cfe9b11532b89a3e19871ca5a6e37248902e20e6bece29e5b3b32ca5a04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1002bac32f63a6446dfd26e662211ed7b3fb4e469cb70e03d61dffe5e594005e8092a5d51e4e5ca51054398e330cbbf97a28930fdcaef592b940c377bb6bc1a3ec9409355a6e349302d9329bf3b5ef8998f1bf8e415bbc2aba13af97b2269aec93943ba7543984b3bfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f26532b962d7bda2781fbfcb530dd47a9dec86943b80954ad6bcbee0883594892ef6ae304e046c643c068ef12cac0fd8c6939f96ed72dd160b0307987f870be933c17b09e1cfcdc1844cbd39d07f2e98c1a3e11d770ef73ce71d7f5a17cf03f3c934e80a0a23d90d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f31898a74922437ba42b4eee8ce109cb672abd1eb0f80830e7f928fa83e4db66d37156a6a7dae457c2dd1a61b16c7d1a81f21699ffb816d93939873121da3c8b84d1ab7c73aa61bfad087eefdcaf6e06ec4144ff6c5f4a5256efb826aedf5f569e697e1c9757945b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca82378e65e6adb31a3f880162be8062f1108e2830c6e9dc4502913ec2aa311fdff6ed69eea1e4afdf702c384528007c14f7a268e61474b31ab37a16aa44bb3ebc6e2254d5111949903d576efae5c8ed8592c30ce2ecfa1a4e3b82c9e89920451f562980a5ac4944a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea2a1e03d1439da0a499f8c128e30001df5076348a788564c5a6344596e65db5e6c6ed3cdb0217818467d9df55df786553eca4aee4dfd4d4984bddf08aa08f6c536d7255772fe0f2e516753da346538147a701a7ab8e0005d4ae542c78166467cf541fd52f3215875c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43113c3b34ca90356653f362f5d1b1f5b63b8e8161c124efe53fb4cbba47e09768219b00bd3841045fe08dbd2a676cbdcf942edf9f7b3fcfc9e3fe05f9725510a062902297986770e3718eb380d1193f461db68b048dc05dacb4d098d945489559b36e3971b3d8ad1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11782b9007780f1be52dca3cb803958fb57e8a76df847fdaa213da0a7c53b596d72ec89681b29fb466ae22d7ccaceae54a065411c54b96af59d7348847dfd998d39d0d3499e3b44e4ebbca50943216e3b6c47d140b43eac6a4ad791c8fff66093445e64d4db400de548;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a27ea12566b45b617d5825a3009fbb49ee0a5d537b558518e14562cacaf1f837a29fe32d14521b87db4b84fc822b16b469ddad4e5a50594bf72a76e59d11a9c1d48f1389e3f37e7c65336d61184bb76ec4db4ef96e82bf39192f85637c42f03cfa06100b30ce9d944;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h653b7980731110ff760e91fef977eaa07354b50ba49ae7ac268f357f9747018782a299643a3e8fd67eb53926f55d9a925a58cafbc6baf3395f0ff03ba3590d630383ffff482f6e26d6d9ce6c932ebaf51096e627e36e71114e15b21336a2e0d24c1cae4f537fd9ea34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e229f59ef330212f24df8b209b31cab271390e026f295009de9ebc74ff0e9683b45aa7a616cb8f6e53f7396aec23b8fff62326a877a8f2e6b26f5ddc34872ba04288c763026b3a7cb71f6fa14795851f100f745955b3e683438b7e9bb16698b0768d40267c0f2d91d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd52b90c05e5acf4c31c1a1cedbadb7717ff6715420ad9a0a31e949710d3f4fbb7140e837938f560a597cfb2dd529525622654ebf6c0df5d2b0c668c0b8ae84a88a0dd62f35f0ebf486ab38543bc4fc700014df0df58a6a3b1c30f4380b6af468a8f1f58fb4ce9187c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0f3f62a96a4e9236cd23ddddb65ea91fa88a2abfcb01b6eb2ce3502c6ad18c6f8751b54e7aefb11129c68dc061adb021c6131b78fb253634faddf35396be9afcbf77791b5bf9f87e157c277aebb25a1f209957b2f0b71040a428122dbeb4260db7ceed929da49e9c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4365a37d1a7a61c4bb88673a8da11303456f88cd036e600d93aac954020f2d24aea27cbb9c8aec06b9f39436cc64d5d93b9f29a6e45ffe4cf338046b24c63bdbaf1af41ae24d0328cb79e4294332c944e91edcde732cba7fb8f64282b7d7f64c756c909c3d0128840f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198a73738da0970202b5ae1238ad1154250ddd1391e6eb8f3f2ad5d36ab01036b32303e7db4038c7f0c746da561a03e35324db7a1ca72ef578e29d8b80b85bbcc1d404b4925e40998a6674a90613ef2cafed8ffe8e14212775c1a6359bbc1a7b9290452e307849a5c93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb524fc68e31626d1ae64f41c84efb2bda49344b26ea20da35b3bba154b78b8cff3ac6a025b4ca15b57f8261bda14c9debf5317fad3037cdf4c7e7e909d3086ffc9708d6b6a24c337a423fb1a5b36d48133beb4f23a958d20bf6dea5a448eaaea1a5db64a7b3857f2ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f9322d4200c46028d0a518292984ebf548a7a9eb0cfb5221919c50614f6f76c9ed04aee74ef9db1d242563f244cbbcbf9bfdc57c59deb39a301695c35bb28e1df80501bc45a5a64d82e68070d256a800f8e84be2755a459262a46c3dd1660bbe38af49c6ec2994e06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c87523a2b92126b773b94fcd62ce7ea9e330a598c5955d9835c1085c88bb9f930844ccfd86a467be59b5e9553c1fdc2763c26508c7aa73c5c5549291dc8f97c696fd1638de887d6edc7053fdba821f01ca77d26308f3c2314ef9a862e25496873028eca0aa660e56b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5d67e743c74213f5fcccb6e7754fdb4bb547a4f8f03a614d765ca87d7e2e4ea2f03f180cf9503ac00e9b43569cc383eb70e4a7dd358deab61a8cf1dc420716f5b44083db0852706e99d909de45e8553b9e389d9990edbb873cab477934db65fdda4ec49d34ccaeb4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had27d32d92d03b6eb14ad0a7030d045d9bc97fa26a338537740c9bdaed7e9c70bbbdc2435f75e482b7cac0454b368a4f718c1b6e158696fa68a872bc8e048eda106437b3524037655fc2186aba22655ddae8085684727156fe7fb3893750424a40233d63939c461bc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hebbc627b6fc99dbb30d5b5ebdef0a5e1c2f04ae44d85d53db1e9d54f6f17028571221c1144fb47eaf8c88f6df51a77a9389bba2a5c61240400ce17b2818ca375c569389815aaef080c981f663bdcc6f1e261a835bbe6f63bd1e6cef18cb83e1338ec5b2c22ca3d474a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1caf9ddcedcafb0b9e51c2d13a4ef07e55a1a5ad8be9d322658d2774f366ef056face9b237a2d5d600073edc89e77c2bd8f82e9d87792d200c971c1d03d013aeca39bcf78aa1838ac4f6d8b4a5588742c8f28373638e09234c7323586b61cbbd6d43f982a8e014ca4e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e1952865b729001e5a6f0ed655ef70ca08a14b2c612ff2015436cc5711770eee8e5365250fdf13843352a8a87b2468c3cfbdfd608938abf121e01442c11a29f7e8df5ad12cce74672ae3a82027839e0bef2f2df9b8ccaf1860203579c537214209f8b3229b56ff2f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146c27337817cebe02327c6ae8dde104fb2ae6546f3797513cffc04329693d6e8615bd9859c17079e0fb38cebbe855c1772afa4cd51bc3321a55dfb92635fada60dee5ff8601b946116013995a036da66b0e83f8384ad60b6eb0a296eaa52de600a7f98b74a2c29673d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109beb750a913cc7d05ae5f5027ea5032fb9f7c8b3139e9a874ffa84ca522c0a3851f21738945425eb732fd9e32991db23fe349eaee2d594e2cd41afdd9edc47cefcf5dcd3715cc0f4ef57e3387a0a9c61bf3c47bcc0860a3bf8bc22bdb5309594bc75de6c85a9a0ddb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa5e43ce96326212afb3ee64e0446a3664146f4ff3f776aa2c1b0fc238380fcdc06992090e527fd49ffb9a53464c5baec4dd9f6e366161a7b9aa9f08dda56c38f8dc48d7a212a8d441f4152566061c9f7abba9ae64670cd06bcd25986411f418b70e945cf1633c56a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h933eb02392f8d880ff3e85ae983755334e3244bb90b203cd9590bee224a1990d9651ca27f94d52cb5ade8cda2fa8141da683553a2ef2ed027847bd60155b065f45b449258872b8249508025e575ca3c0589bda90ec6bb016d2138918c3db27bb8b429667dcc97eba1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a694d8012864837675e946529526193549e3bdb367fb1e548db3a8df1972de91e22b6b079a2af36f38932e4284fc596e29926f9b26582b142d45960cb21ae32b4e5f8167472e38680047f763f6e030b07a159b3f0beb1890a44caa6a8d49b44477b611fd57bc624b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1715ce876db774b0405b76d22cf8fadd78ab57eeb0af819ea7b4555ffe3ce64bdbd1b229a6b003cf27e2a28060ce3f9ace4ed7881c4bd2dfdb041d3c2286eeb406c647a1a7582e5927222367266b1745c24918c1ddd69e7cbf186cea270f40e863387a7f6d8b6cda9ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136d4b291cb9ae48db248f45bd07e7cf94084e57121fc28d0bccf15f78198e1bc9f16747363f2be70b9adb693cb640fcc7cb928fb8f54359339d09d25ee72cf4ab1df688739919c3890a82867a44e91e18e14e6cbc22b7b07013f54099a094cc937fc09a5e9c6ee53d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13051ec2dc1f4036d560b581479d17d2c541d9be8dc315289b871ee7acf9ef1f9990e2747939ad46ecc1a68dbd791d6eb1633440adeef86e8bd44929c97bab6ec032563ece55394deac27919da2f39190cf923f528680578e9ac1eadcfed30e4e98d4308969ef944ccd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b09809518bd62b297090829f289eed9c52ab5283a23be6ba6072c31ffaae9aa6978f5d91879f74ec4f685295968c634bad3655057fbc8defde27d9d0d313b8278b53cf42686a2450001eab680c13fb365d4595dba93b4fed04aa0e1446f55358eb9fe8aa4665343af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd1c37e18df19f406f8d018ed4327cacdf8808fc4eab6d6d9692158ba08aef4d4d29258441fb4f3bccd754e35624c9ee3a0bad7771f70c8226436887772a7d3de5c177bedcf7eeabfd94ab2b6c8a1774ff4178dbbb537e69b60da2448b86a64352feaa13fe8aa7ac45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109905e8da559c2b02cfafe8397344e8aadf99dc22a6fa2e37abc7bf34eec89b83fc30760f9e34ba208218ed29aff88383959fa20a47c3c4f22fd39d696af9b6d85268876202ad074705062cd140237970583c64b7fb5e552d098d99ba14e8e2f88041f7b691aa6d1c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a087a56dcb47127c55c3f68c045c06d97a5a67c7e55744b24f0484099c198b192038b3de627665345bc0a1b8488a2407650ea4e84d723002219836189a62bf671e77df2aa80d68b74f25f1ec1145045bf2942c45258f71aa23a705812d570232b7269bcba6a9ad811f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1110a333d890ba55fc9c84d21c05c589e391d57c402fd3b4ecbf1d0f96d938fd0546877c5b8b19bcd87df19c0f6958f9e66b0bf03140e0f7051d3bb97f80644c6452607f2a1560fe0452e77fbd5ba1e8d8ea33588f5bd20cdc7ef8ccf250e1bc39290a9dd24fd500b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbdd621fd77e82ced245d6116f0c61af8803de04f7e9b3946fd8767ea5c70e6d511e535f44d59efffca3ab54489787e4c920c48291a11e855f48b363c30d2f3769db220b387fd4c2b802766517a53e8ec17efa8f7335c3afd66828a40873f34307d52a494196c95ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bce60c897f80ac1fad6c29d82ccdd5454b2685c1102eb68f21ba33375d1fab7cd5550c8ae6f3d0c4303f502289b1252983cd6acd336b73c2e527312ffca10738427b484a6949df206ff421df107f915219432766048457c51742cd45c732cdc1df5b760a0058b62d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a07fb0e970fa726ec88f029de7647a866ed6501ee50eabb18bfd87f1a15b1e9b175beba8e1f20d43a88f4516a841fa2fab28295c5ca2055a5ff83984839a0836e57bb00e45400c03b84af99ce2bab64c72284f506bd1ecee625536a0691ca1a232009714f7ca7b71e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3e5b6977680a064787c7f2d721902c7fd6de25ff97e9de3ab81eef0b9b2eac70053a76898320f48ab0637e1069fd07db2ffdae7834d48e51f8c97199ce0704eddc1e4a53b06c8b714205c3cd73833c7aac0ef75d46cf6293c156ec9702db62861c6edafcb68c6838f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9c49104a380c8d7153c03da11adb860f394fa4cf0c5d50d1bb867cf81a07503c2fe1ede39be8dd1beb99889f11b961aa4fa123a4ff47ac31cbda9c958c97870e5c8c41ea5dde607dca15eddc08f54958a77cbe221391b76dfa2a15818e9000edfb18d1f5bbe95ed45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9dd7cb28c7537890e71cc2db8b3953cedd4782974befebb9712e339c3a4ee0fae714966479510702b92a2ccb3b4650a65c095aa489dbf60153d93a5db6923383e1d50da825dea6101dba2efc0f34b742bffd9703060b965df1702d19bbe93a137633001425f21efb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eccd1436d43d25e0695a3cc53d94d5bf0b795b873ee74f0d45c46690e4b034df17723097a3977999f7998654c672d8cdfae1942e0bfadc28bc7f1658a7fc3c302018371732459241188378ec3c700ab3b9bb1b484d6c80cba400927248b000020e5d863b16f0ae46f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22009127d4ae2e4018b5b1a26499c406931ecb825108d753e4df9787bcf34bfed0763ba1fbb09a2bff18730fbf7e591da739d0f5dcc4c5d1897ba512af2137fec3da5a6937c119c6b3ee8013ba064c5a5f8c6a7e22635b3270f22c3a9c68b093310b225fcc0c57fbac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f03ab6cccf96c8223352b7cacc32f4d7915ef33978b25c51f0108f56f70a9a6bfc48fc68e7acd73c487d3e0b0f35445fb0c4c4e24ec37009d016d26d0043206ff81b8721404b77f1f309b9128b34527122e3cb7fe1fb64d271ac374cc6b0d65882739bdea419a4b6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1fbb9672619b4f0a0aa8942049aacf9d9a947b31274dc760c0e358072342f95e45bdce12bf2760895f3b420ff8f2769ddbab7b0e68faa6572005576666adac79baca5250cad5443c6e78331bcd86abf2d90e1d5240b3d2dd5131ed8bce8804146613508b8cd768b22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1907050dd00d0310527b1fa07c85ea9db179f2adacec9ba31785af641ee6168c11920b2e66b2585c1e21918f91a4ef992855d622b381b9ed3f80af7f50c81d9a104d3d9d9fb1128cdd110142c3e29df2958a7e728a635b7c355c22b928dc220d99d0102f1547a2966e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17798ea6502fb841324dbe326606acf68cc229187e67de5bd35d95dcc6d523eca81621ea5674f886453633f2cbc06a531dfc8adae7074b96f0bbd6381ce7675f207d39b865b3d2fd21e2a604eac6da4478bcc154ed4d835d5a4e7c260a459d7c134b04b52c7c4b63e32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4828d4df13f0e3af8991fcc519eeafcb428ed7270d7e4a7719f198d218ad977f16034f794cf8deb20c11ee1384e1f3af106c7480b2f4688f6953f2dfcf0b38dbe9d05f29f7bc5b85ce7c2625834122e257c4f1645390e8b487f6e00d2d11dca719ff22d06c5154e181;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4079044e41a80c943dfc91c5136c529f2ccc90d5cf291ef36fc98cda46de5703b6f7f2b60e35df0f667b4cf735dcb27aa973be1f73ab4b13770ebd4d223b1fe6c3f3a6693d3a93c256572ca292c82cffe1cfe2a48308fa4388e2dc8bd50d16f42801702ea181916104;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ba8edc1d8d23fb82e01372299d83361074800af948128568da450d61a370f9a97b5c1ae255a0e619972d3f058cef8c10d2afe17b9cd8e0500c3bb1e3d8b5ddf5ed21b12f772d182f5590e868628098f8988300a4096c1ed07fef7a9f00b35434fb68ea27964ac0911;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12496974e52c4d918aab6b0cfa78eca0a9394c25e6664c66ba3567200dfee09a5f8492558a04b4c516238d4ff39d00d12d6dd771f85791c9846147cec031be4c3821e00a2ae495f5ed2f484b94bf2e2d727f006a27d2f193765308e782541fd5214f0ee1aedc99f07b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab6e926eb161c400e9d309ef48995523b1348a75a68a9bf3530bba4630f95e25151ab6128e3d17781c4f5a665ce5d8d75c49d7f51dd3edb724f9ecb53426049f562d4308c156a75620d4b0f104b1bf779104530262fc9e681d53eb3928d70b4f33dae003e657a9b958;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f741a26826275f5fb71498f9b0ab670144b8779e9f06f7d46eb5d0bed69b4dea4ba988dd66137608e652bb73342d2a05497ea68ce852c03c85e02e1d476b352023af1e516a225c7eb6236f33f1a23886ddd90f4a9b96bf5740ae894dc0c9038f54d512b8b4750d1e0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b419ba3077c3fa5a4be429f21be40ea1d4aaaa424b3bf8bbc8be24b0f9f40861e7982e5c7b9a1886beef030cd9a0132c86e18bc37b04bbbebc103b2b80914c5f22e598044b7721874aa5d8cc25e01a9c7748675c70718abb3b9fc4078f3f980478996cd63c223ef850;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95ae77b608eabbf9ad2944a74036e7fcffc73e013cd3c05c2961f0f8d9bc3dbb4b8916df3c252072dc34715e1d8beaba5dcd4dbf0f5a3d562555c86404d06e3737b8217c3aca828cc0db820a4c5dde172c25012c2c526e6dc047335ada1ca31e6fe3d60274c56f5072;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe54fd858f8192156c6df50052d232db0717ac9ccbcb8ce5a22c5ca28b7f3789c4baadcf89fa8a0f27ab8a7c467bf4b1f00bb3f51fb35dea2df2a5bcae8e1f77aff7d6184047ac8edabf764c76b515e8a1c0763acb3e4c70c80493ce8dcfe16fac105f45129f8e3a60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b79d9a04366d5b5af3b1fe07f31c940f168e7a3628138dcf4f8f3ccaf3fe227e4b39b6973d12f046479f5901c352a5a6f3e83ac76fe49aa39a2e96efb9b32ea53dfbda158c7509c73283425931385ded517ef1966670b91a3bf8f18a86c5f8d29afb5cd59c9cd31692;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71710d8f93b1115975060e409e4b99bbbe506ab2cb545d6f44b9b756a27e4bebf5653368dff29c353c40169d0fd66f81fc0e653974384b517d254ca44d9293a116cb633c35a9796962fa7b9e589ceb436bb4059b047a1c08e07c02d2922e9c78da9e4701ee9dd094c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25facd3ce5a3b49d51d8dea44da3c0e726d28945605199c3c8e3971e1521d4f562c8df08fc85e493d9bc90e21e6236aa1b0601d963351d0ceb9cb6249abef3f8c3c952e99b7ef0750cd222c554b4ad794e2353320f4bd70b67bcced55932d23726386e4f198688f17d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffa8d4cc68b199abf154f6d701ae7f495a114c4fb1b8ee0031ef032aa1d5cada41204f96018e5bb3445459371d1bdb11036813f9b90e2e5ea110399489854b398781c547b75403c0f255ef878b70ed54e95d485e0bd083c719ae6261173db1f9674e022669efc1bed2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e128df20cad52f0d07a84dd2f007402df9068ae9c90542a768941c5aa79639594af5b085261b155df1639e78059b1bb8f8dbd7e6f530f9346a8e7442b978159696f7c8664a28794d09b8d8c8fb315bba0d777393215c9cab5586175f16548d1d1bc9b64c8747e20de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10865fd96a3e1cd3d189b948d011964a94f76222e6af003a7382207c5f1e4ece6cf909dfd0345755cb133e8f5fd6668c120efb898579ef87e5d312a632fbce2da9bfb06396bcbb1189262163f5ea2af016baa41cca9f990419b22c57d4fea2ddba43cdc7d7e82315ebf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h293db9c1949050919801f85c75b8050e5cc4b51da9f4665cac301d9cdbbe51d152f3836e18d1319091fa1c60f31c1672dac1d5323bd23dd0c72d971598f82777290bfa155a1d7a32d126633374c17c77aeed54746cd97a1044432d5ece222fc5e311eef7e9e7cf677f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17dc719538bdf137472940d4f1a8d1cc12d461e9baa3fa966f49648a312195952c207df8da856269d997822b61d06c02e480c204bd501cd613a68694066ccf7e478c23859fb3c4d64579e0b51e27901fa4328fb78975ce0bad4fd204db9049b0df15b6278c2916df4cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he609f0428eda92de4db96075a02351dfbe7202e3218b491188c215767b0301880931187a485fa416f262c4baed85c57975c32706d1ddcce0aaca8a4ae3d183e4598fcb788640f82787e6527b81bdf70930b34ba7760ffcc159450e04de17c6fc7bded6921cea76a03d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192677c8aa6ac7b613a25903c65ffbeb2a154a2779c4430703ec53c8cc07de235593c21ab152463c66bc311b6d8ab43d656deb0f0292f9420714ba08cdd6861e7ae27412ca3a910e1fa8e40a7f22259b7e73d82038266ce34940af417e2052dd541b267ea9f34bb65f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8906eb46f7b31b2b47b6d7a7574b23fae638b07dd3741e9be761f0c087f5ae6b66521fd0336d96b868ec28f335d8a49b59ee7ab6f26c5e2f1a76ffe9c263e14352078721cc54e372864c4fc576c24a73668c2839d4693c9aa8cf1d8455fd1d456f65bc896d4eaf20a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d574aa1a45d74d8ccc1fd5e36a749ccc92042f50ee8cd995751c85d433a587f91e66a19f6fabd666a8cda892e9fe3505548cccaf4e901e971e331e025a5805f0810b805829f1af5ae9b0b50da594c22a91753e851c83baf5153110fbcc7063134a01466f28c7c679d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111f24f3de138a8a4e3c4512207291c00b378482308452d4cb3b64cf27e4435fe0a1f64509133a3c7f5311ab123ea6fae594c11e1f83d147d7bb18079c6c3b0ad51f1ccc2bf46f0e1d60673be2db8ea4dfe0fdf27e100dc1c5d43f7bf2ebafed75549b75d5d145d2ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161f334c6d6f1af40b07dd732141a55987c567cf395205e389a3519f52d52cb09c515ee2c37b118eb40fde783154be8150e822b98272d7d476c2f8ff2dfc89912fda753131dd122044754da8d67c0eb6b06fae58b658dd24619ba107ef99771d3a2531159839697f68b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10974b26894c0f1cc31b46a57114e0a6dc672d3775ed90e33ad55e2abdb2f8d5948cf275ea1f6ac5e6860c8fc0cc01f42659419be836407ef8d8f3ff9576982cab142a1cf606885e5050a9a6f948f16cf7099ba123e06d11bf759fd7025e99e97b7f03d045f56d33148;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4f0ca3444abb0cfcfd2b2d7801c0b1e348db8704cff45749825d091e677b4683749c09ff6e28f69c5cd2655654f3bedd4e3b95d9da8fa761dc8b5d30ac35d7f8a34dbb000d242acab21d3fa49fe751602f57b1c2bd7b6497e6b7febd04c9d9d895ad5a81834dc88cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44d317d7ebc6efc38b82bbba74122bfa5424bebabe1820568a8802fb82d9b0ce1ffcb0a2d300738af97069e23e7f1bb97851bd098139efacc904c86c3429864cd16abd13c1e9cee463336249fd571dbd45c11e8b115771ca04c8ad9b2da37ea4d1339ec7af996a8607;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3f42d5db2587ead9c807142cd64243004f068b881e6d9c62e72f4e787379d21f79605be6f8bdf2f3354bf26c95b29a976324e7b3b28110f6d63fc9116358ed2f7c51e40b50e935dcff2c33f201cb531bae6f91dda17b0c90e6e9e6ad9e4bbdb9cc5a8953d7cb629c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e7178421c723830b2b1fa5c470e55be759a1053e7ee54ee8d7b084dd20ecbadd75860ead3ebbe6ffc61698603f03467cb3c4c1cbb315b329449f8d01754f88772983a625190a14d619bfd5d726f62aa251d26f3dcaa8853d74502b3a2ce519ef14778d54b7e6f0345;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11fa989465607b5516c2feced394424ce344015eaaef529ec58f2bf59cc036766dc97842fcb432cbed59a64df0e3db10a44cd166efad908581115aa3f8cd90bade691eee9bcfdffc36e17a5932fd37313e616ac913544195ef28d0be26478ff11a2bce80b20633de153;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f6d2e7e171750cb1f51022d586ba5baad0c5dfac86c10609fab6ac26e9dcb44cdf420f342b9a3b25cdf03841f1fd09ba764362429abcbda69d4aa9f9588da2ae939e18b13e1a5f3b757f5b61ae6e28e12da9014f690360f5eda114d02825349ba4c4bfa39a42f3148;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112e23260bb45f9ddd5fab8a4891a2998b45108fcbb0dd8c7d1b296852e436157d4f3a743495155bf871f9c56b8fce876bbb0bc200e7440f5dc287c549e488fae82a372776827b8a2d26d39271b40a020984a7bc86fcb2a74cbe6a29bded429797df53933eecb058b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1763366a606152fe3e95a4d912c90e538d950a042eb370d4e77a1bd4d8ce8fa85d848cdedad841f2755b727fb60db0d25df3b9963d801eb779f6b1544e8353b121870b0bf7ddc5b804eee518247c8d34fca37eacfa9e77cfbbc34cf44b1c61e79f0e217fe34bb27a919;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f8f5f1d46c936b8c602d1c82bf3bbca47d1e56b287bcbf507c08b89957950aa91782bfe069965cc3d651056efa364b66f6c10704e8dc083c7363679358a54f8567e34ecee76dad114689dc5f0af35dddb2282bdf49c06c1efebc3be83b171222ee0a66c2211ac41ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he188ff6ca10343bbee0b9cbba68da51864b7e258c3fd645b97961e7471f035768b4492391984d8197e757b089bbbdc1f5cb34c61e3e70a07762bd28fd746453bd2afc9ecea200193da33b69f4538637b7bb26f8ab8f48c10527629ca6017a782ef1d7dcfeeba91f136;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19aa37ee5d3ba1ee9593f21e5dc7bf29d1e554d0adb5599d74cfb5ce6385e405828c408125bc9e2f585e3214d1d4c85dd01a3dddcfa42ff78dd92ffc79afe72054d76eabe4cb922b21531166455c7e68aa9a50de7468460f54b1ec7ef90dc9a4914b2e5efd1bbb03f85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf03871c635aa991d8b8459c07a3642a0c898dae56d84d20045548965a90f0db4438f5eb582e1148440e2d45d4c0980f9e2e98d2e2147793919e1cc9db89c148eb95aea7f7395b7d9b31ea639cccfba7feb849178ccd8f1836af93ea4a900ce877ecfd1fe6dd9b3572;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180483807db7f36e6099921a249fa841077090706d8bbc5042e2d44c3b500b2536011b3ef8cc6c3e812c5e29896e3741118262048058ae3f70dec5f90c0159f78a4810947992fd2bb8928a4639c4448f52f8d94c550bf82a157ceb7c8f22b00f3e776a83fdf87647f99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h846f36dd73b1f2f62cac4a8e201008afb5699456be9e25bc8f6911e3964897a0c4e5a913a84d34ce3a0e9602f6a2a44ba8f249259eeb82763ed0e9c2518181a35591d12098be49eda223ff2efd151783eb4102f5dc2610ffc5e42532b11f2b3bcfc2af30a9390f5057;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161ee315109feb0d57c3cf75f0009368537b294fca3e7f2c2b7c0fdafbac4f9071ce70c5b52f4b878a0cc01a12d7acaa2a3926ac319fd6528dbe7dbbae7c5b999c275185863d207e5696c30a4f1c124ea5a07570f55ec59e0c74bcb250506d02cad14658a16f157d1a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f9e5a5414901e9475fdf1a8ce3b7e66f3925b02891ecdf999d654a19bab819b44ee5d7d28e7317d9ff78422fab00c7865e1c91a8cf12b603318c7ea52e7a477c163a4d33a7f6e7f8566468d89610c87a8173ebe48af4a4d50a9aa56f50b5984018bf1cf39dda61361;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf838fb5f8a2f16f01965f45fe23efa9feb65b4326c544264a9ebf5189467a0dbe750cf61e8194cec752f06bab53bcb6212cd94a6f43d7e3dce1ec1609c09e5b93d7f8945042ab59d1b4d43b0f118e6a184c427d7ec4718f499624c206a7fbc8536664633764bfc1441;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120b4e25f763153c590b4f3d0a22b437af584221197038e718d358128b99349a4e23020f48d7c0c2c3d69ed8f75615c7d842f8a75f5369fd2e1f9ceb26d3fffb1c5902df13b3f796d896c0b6779f82d7f2a40f62f778a084d59402d09992412b28134615c05cf63654a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b00013652629945e977f8fc62861b2d18beef65434d1cf4d2951e6083d08f4a5353d2aeb511c5d922e93f8294aeeeee9041b122b7a7cd0845eef298c73552a3a2f77419a7c2687be461dd296b449d1c0ffad3b42723b082d9e13a1ff85adc8ce427ff9d9096454250b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b56edb3fbfbf0d766ca78f8055970dfcd563c25c1216ded2fa60b2895d97923e675ac0f198254d5fa2c62b0d02ea699dc5429d90f37b3c9594790f0b9913a6a15cbf41da49efc273a3e4183a72d2b44a7e1d3f8b6ce6d864b2f69a5426043c2f72c4df0a273b0b4d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a194493e0b6bb8dc6c481c443a6051e7106af2bbb28e4b39ec14b49f65f831bed42ae0e79f16a06bcaf7c138a6f96992718143911f998d50d16d1b475957cd85925ce35656b735573ecbd651d51f385ce75af432e145ad230950762825942197f3bf9c5ba20757117;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a80a987a694c76aac05da696df8d67b9b7990cfe04e1218f1a533eb09dd8eebbcabe72fad0b539c3855146cd9319762c9167ce72d04078533f72e054a380d314bd3faf7b058489438fa8477c7df5769892a8ff12f262ef33b080e33f48eeb334fbaec5c62e21eb121;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff9c3a3fcf359ecd0faf74f1943935ce106723dae904075552e2512bb75a23738e8c85006fa23254fa97dedfcdf8581acc9d933c990c52c197c11c8049d4edd6934cac7814103ff6d2feb2fb91303e051ea851b8810e57eb79bf9cafc0f702cf85fa1b9e1aa785629f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b7aaeffbae2dbcbea49378b53f82e5d08148cb615f85a4072090f31b119957fb348269623a67f7277a96c8a61bf7f7b260571f0062ac556a6e74e698dd3ab7a1b3cd0d9c8e972d8db307d08fbddb051dc00ecb5b989097cbc17f7f01c5fe73dae1ef9e21e9363b612;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141502e7779e45afe1f3967ad23302ac26a1742b9adea4821da3a3b38190211dff275307f5b2d9e5951733b330e98c0edcc568e907ddbcab077f8c6bddd0c16505b2485cdf42e8ccda97bb7ac01cd57de486d45913b1832e5b64aa9d1df132a73cd952e59cfd997c290;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdca66ad4991c34f70e39d37b3145b3c607fe7afd8357c4232b023d34bf11ce68f718fe56286fbb51311156a78e9a1518da9d53c3978c68e78c54d4c7fe167b05ba790a455ebb80d8beb0f2f51a15d3184dad854a40c41efdfa3e359c7a0d7bfc05e87d4bf83e75d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4388636fa1a37e7def11db081b418046980a6dc97f9aa85d3c43b7cc2394618b61ba7698d50b31428b71f9be3fbea72218603a9aaf6cd4e80e6fcc11d323132f5ec2e9f0a05c9b4aa76cecc0b7bf78de1c7bd1e66aa74919d88f5f7d2aab09d20b82bb69f9f410696;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10196efa8cb91888b2124274f9c8219a3da50cbabd7d64405a6e5ab82030da8f06ed657f9a20d657b8d53a1cc8b9fdbb96081d225a24c20de6b987195d8caf0d5626e77398699dbd0a391807286c4f005cab7680fdc54ff479c4b2ecd6aedb9db937d047a03620b37ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8b82c4f5cbbae0da98e969b44936893a98b3047e114edd14846eb65b906c85727f988f6ff1bc06192141a5436c395bff5eb553c772facf0671c9e7578046e0c2a7b790cf9097d1797644e78f4ea19f17c9b371bd79a3d59f0ed25904c78d0d9aa2347d56d5e702a3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53dc436abf06c2c76379070748b7f383226fae7b944ae9a2105f394498943383c35cddeb3322193ed32d1ccb93e0c6227d94de017ea68aac764c2b13c1ba1a4947553d4aef2d0f559c7fb6c17411d30a48fabe8525028cc755977359de2e4be61ab32882d3022716b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5a28366a0c1fbd8ea286288ef48dd87bcd4cca611e30d2534f6fcb2f0cbcde71c98cae17f51d52c8df8f03c405ba7685c028ead3bdad2ff9779e87a3f38d3e467ca7b9e45f47e8cc7815feb2f12306333df60ae896515caff986f75cd119261b3220f3998f123c64b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da7759ea2c204fe5bfc6e98b5d17405e393880f6dc28baeef8243d7c5e2b9afadc90a4ae4cae55b8452589209e4d2cd9dfa7215ea9f20a3732bebaaa400b980c09d8f73606d318e9592788a9f38c994ee7fd5d471fbfe57f919f0d41fd522319e000391d7014f1660c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab5c4520f660ecfbfb04188c7b6f7f498f7f56b8c8f8304a418f24c7779f4be283f2d7f8e26bfda13edc0f0b85b611ae5a67f2662c326d95a3248937fd4196c5396705c91b7a85be35287fb56bebb5748a037726653be1e71e6c81197ac3c11c90a354b980121f6c07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15011a47fa8cb70361dcdddbf04c13f4a77f3556b1698bd9f531a9d4dc1daf5eb531fe7f16898c73c887bbb1e5ac83fa117c0390d21e77b842aee5c9b0c0dfb35dd3374ab9e5fcbd91ab2616d51c6bcdc484fa3528f365d9314f39493737903ddf108421ad129f09173;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146b1ba1f78c0cc5ccfe842a09f77e21608c7ccc67d5f43740249fba1c32fae4f9d59d0b1648001507f56fb3389b80bbafc8309e92659c3291cdb82c036d7ef9cad494fbda0abf049b6f16c7d4e5ecca77c033d5577256ce2165a69699eaa48a8e9e57f395fa8b8b7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h798a8329b33a5dba46a5924e1ced0b88ee596befd2d8c8fd89262afccd00a80fd053f9173143722138f1b08dd127fba8c4863532d90db7c46ba4729748581f6a3bd992bcd636a1a7b4cb6a2ed9d31bd2a29c9ef921ba98415f0818d0b387d2812b6357006990077b76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c59d0587218984c1d00ee295fc4abfe5022f21f490e4ccb00508be59f41e1945afa3c0def331d51e5a8937b487dcb02e54899673e79239a6872d9c80da0679600665e551f782439b42bcf8a551fa3cefe787491186b018bb41749ea5329fb03a1e3412aaac77d6b66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59d0895c57fcd509a00eb955599dd6f7e3b0d57d131e8a85c26ba8cc5f31568d284a898156601c1ecaea01038626ec34805dc2a83ede6b3493584cf02ba1ec7f5640bd2fea23398d542ba9d8b3206bf1f64cfbe08335dc814e54170d8d60e5096cc950846f84c65134;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7452647907c6a61398623b551dabe4c2e90a18ff2f24f71dbf37ead38a7bab4efc33504bb799df2cc41ec665e9e322060d07915593c51b4d4533fecb1a0dc662924f8b6d3bbcd91fb58e7015c1c6606264ac09bb6812acdf8959a8a1ef78cc1ced090ef537773bc2c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9e13002996360f31ec14d1aefed0189eac03abbbd68abd81bf3c173d28981e67e2d8c6f8b9e12f1c8f1fa43dbb78629446b6845259401d3da3a9acc823ea5ab8570b5d0841e5894bc1ef0a50eae13ecf020f1036d6d013dc5e9f0ad1a61b41942bfe75f583440e110;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c1a354502c70c425556491fa74ef2fe2a01fab95a3cd85e1cfce187d8a5f03cb032002523048eb4abe10d468d31e5ad161e569aa7dbe1b788e65d74ab59c16003e1cc70aead9cb5c9da1e93de3372adc02cb24e75a1bf395a3932e06d04a065c4808b70ace3f709ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50e03cdbc4e6978c93d5ac314a465597f0a0cdf2b5cd3518c28b3e898a42ff05f7c2f76fea5db761b8c15f46508dc23939de49a16b8dfd1fb4d0038a1cdac432826e56f6f03dd91516bede1c490a2e4ce1a126cfe214601ae256a4530143cefd9d3b734473935d28cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd610d23efd04cdab8a2ad1d28e0b2c7ee2dde456dc667caf3de79cc56781694d3e337d0a50b81a37f254267c52a89a0e0c0a30d6dedd11568d49bc99ed20ed6d63a9c07020c5359c508b1bcad0c5b294826bfbb95fb68d1a89a273a0694be75e4095def7ea4f02929e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152e93bfab9b0751428daaca8fd6296559197e4800a4d27b9af93eae50000c1b08997ddf7d855eabff2f3f9caf6616f6b4c510002726a515c4bd04bd12f07a239dfb02bac4610da4c0055ec4e29183ef378e368af7bd2708847388063142b84392fcd572e611d64554e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6030edd45c2bb017ec3cba423896d5fa15b156c4e4b8109bf4b189ce29f823ca75b6b8bc8a752bc133eaa2b50d2318d0d1368318a105a9134659bfdb80a9435eb7379725f695d0eba147529183afeb8d548f0b6cbb1cd12333bb1f75c4c95ea66b1331ec4490f2750d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d524d3946902c649b2659752fb20cfc6dbf6d2b4273acae96ac0ec167cba6a7d481c05c2b60223cf0573b6987ad9cdf2507c282898a384b0b3e90bc06a43f651507cfec541a1a1cead83fd524a46b5e71b4fc7aa3bcd5d057c9d56d7dd453f4aea2e89a5092cdab8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41597785ea3468dad77c115571b35b8b0a24c10c7ccdc1f98a2be5049c35d552691d60880ec840aed6ccc277d522cae83c43282a85006373c692800a0856f09f8e4711b847c6c7694838ce5936a8fbe801aa80cbde4f819cf5bd3abb42f2b053434a33bd9995c2a971;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d463a0d25a2835b0d44f11e6eca79febe9ec1c1ad0a01f9b1e8d8776e90ec1e9bdfebd71375e6c38cfc675f68cba2fddfec1a42e2c6584af5e07303d2da7deac65e2ad6cb79f95ef54afa714ecec9f16e5dfd12c018cf2077ab1fa25037adb2f4cc38ac31a4218124;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d5094082fee8ba9e0ae9c2f977796b565a3f70ebf1dab5221f0bbb83ab5c56986a0478d2dddf9fde4cb3d392de5cb3d0a0c45678faaa4029a1016e30ddfd868fafd4d1efaa8c1bb00ef3820ff3c09a2983236445d44aa2502fded8b9be3d4beb158902f257775561c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12fcb025ae39ea5be1f9d77531436c8f8f30cafff2cab4ebbf3365b8e3b253942e88d3053bf8002e1beb4cf8d788c455e55717118b26214862ddac0e799a41b0a0ec2b94b2360b598b5f41bfc0bdf1669eefa95143137a52c76e7833aeb285e756be5c16f2c1bcfb9f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4edeb6d4f180e718707c74675d56d42c3a731c5e4230f9cbe6509200856e950990c2fc97e7a3f58e5d38bb5d0a5975cadaa35ef3738cce3f03f2898206807da419b6283dd7f4f917da41dd5283eaeb12c4352932f1016b618e26fcc3ed2c3ade0bf5d27f3bb590c2f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc5137055677688c77fc56e51b36cec0d9f69c2584e84dd5929f2ee0fb01f14850e53ee9c1d7ca9ff2c6a2f68f28bafa10715297bdd9098bf290568a8f74b58955889543604a86a8332812457298089b87b23df736292c97e7fcca212c6ef8e85ad793990b3303197c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5f0cd555cdd02774283e8d4990878fd07816a9047eef0fd9ac0b07e21bf884ef5bf47f4d97a5c5d558d69654d88368c496e20f5decde3d16f36aa7d36519f2d52851e4035cd37fe5ad1081fb1a4d0771668cf3b54621d5fa854043d0003f64c5dc681710e5bc9f72b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0ae902edd758f73a594a9d681d6b632f65ee0b4aff783fb57c4016d070533294eefbeb72541e96e4ce68101c88c068cabc67bbfb4f6dc27eb616a3ae62e8e99867b8f641f2086e073dd688e0bc4bb701e0c44123e24db3e74f88cb78b9ea96c4772b748fc6d1264d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec9fff632e9452c9b20b911039050965742552441cdae0bb8ee4d199acbc09658757bc9734beb6ebc49d7886f59fecc929ede60da54f3799d31e6260caf572f276074d3626d020dd592a1ac7aa571eb8ae900b38438c2298ddf104d1ca2d6f35bc531dc90c14d7f5e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c4f14981fbed1bd03e94ad273de5b0538762ded30a4022b35c566c38115927208dcae34275674cc68a97bf1708c56552642e83e06775408c71c98fafc4377b0b226c5b65ffb7c9e1293b8fbe35a7dfaa870beb20c6484ba7144684a99cca8410214401c49279cf75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22833e0bba778b20d0dddc561395b27f7045e5f6b5d465cf168ea9af086c60a0c82b55725d4ccaea6e0b09bcc7f22921f7505dbc757b2ecde62bb59fcbb6d91e79e81da59c8a64d9a3e3a4d2d0af591668389e17bfefe068ff0511059a9867dcb3df4436587864543d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffaf7db69c2165b202a6ed90ef3fcb6742d1aecece9bcf90feed171efc388a97d6620abfc49db8145824ea4f2bc44e0b1a9f71b3efcc2065223239ccc8faf878c1887f6ff6b874cf67c1b89d9d884c63690cbbc1ddb37dcc91629e48619d0578231a7e7bad4077abcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89dd5dbcd7d98d91d8b588b6be69d443dd7d3d07a7293e13c8b7d71c85fed4212400e53cbe22f0852e50b8dbf8a5d7a1bc279e25e09e41dc693cc83c320a6a0cb4d990fe2c3268a1c7ee330271a414a4ae82f4757a06d7c6a01229a01117521920ff8dba247fdb7b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'habd4f669f3403ea26dae32f2d7d916e02009597407fabcfbcdea110c71b1201a51a801090d53b5620db67fabb665bc542f30e8d6c5ea4b909d2fe3443c97214bb7adb4e5aa405d907fdd268d683df03f8cbe2a17774c65d292be37c576c0e5f662033fbd037770f5ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82f934f8e314de4cdf316d37456cb77b51c0da902c7ac592be5c9d591b213dfa0fa415f3081122b65751999a37bbfe9c7d5ec799b2e70a1dd4a0adb19999b1c2b90ef42b64de2fa246fd860c4f0c331477a32ed8260c45871ccc29dcd0eccb03c73c949cdfd2b9744;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dd00c0012f828de79b2842c63bfb3e086020081f5317f2b44aa6d81364195a91251a0a8639f4dae55ab3a5d4fff9a57f9adb6478bd18927d6e8668c1573e2a8082ab3915ef724f4edff50190f62bd71a2e3d006b93cc52c0a319a3edf7d65b6db46ea5acd174889be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h659d38f80d98ef001c1b8a576b2475b2f1ce1f1ad417338cf3fe49ad31fb25473377de4b2bd6f0cdb58238da10aed9ebf2e8694cc5b60de4e0ac0d730ae702ae891846cfdd9b2c9b458590287a1e74ba223d28c1e36a7fce2c287544c3b749dfad4222f43dc827daf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108c1b356ed84eca0f4a309aa06e760ffbac00be9ee1695ab58eca2f499787c3241c8691ee74d16f687876408f57a16fe3cbc2820d79bfeb578dc1ee8646431d35f1b9823e398087c6c07b1f29c3a99223894f8d5cdaaf78e24a9fca7f651e3006cf77a212af643db92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111e1a575b07c2303c73fb39cdff030d9a27422c97dd96d6cd4b8567979b4558ac2ad032acffb0d7093514c0b7ede3eec712198609d39ed37393468980e331ac8da52e125e3b0c24e29889a8f90e02927394b181b723035b2776170eecdf6e6dc27248b4a6f7e6c95de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45bc0e05edf93b9c2d8e894d58e7f8302803b9b258b3ad371bcb35566d391e79fd2044e7d799f78b5b663d8d565d86f113130a654746b2ab01e21bd8d39656e3cccae6eaa3e27ff790f2a83a68691b675f3e1595c4ea6a89437b77aea0907ca6ded3429c44b3c21ed5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74f398ba5832084eb7bd4e6d27a8e39cfcf50242734afa1d293513a874e41d72f4bd13864dd31246b5793e7b9674b75ddf0a9eee604262711881b6b6db634242b45125197911e77c17ad4e746677dc1e862ebcfe9f5e8775041a2f88b0c51ab02d944ca0a721c28ed3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7eb5e5dd2c149a5ee6b16a1612ba6967325142388bf50e22e80d50b218c40a708689efb56de1bcdcc487960d550d9373802556218e411672743bbc4ef62dcb948c8f74d51c75932aaaf717487a8e6b5f30eb315f9bfd78265fb03ebeb6b9cd91489c8e886a4375f75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1267c018a8f4d724b461b642481a7a96f09a101deff23b51362b019ea624adee7bbdaf88fb22a27b0ffcf51a0ea8f66f3a3e18ebbc4aa5189fd79cf2ec213c70dee2f8adee1cb62819e1eee994f1ecc1a0694eb1a9a3a64d4cf512457de7bdba3566110c6240e5388e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1192f5ad80132eed3d0b681c4e512934c1e4f7c53c209db58575cc3b0a12e93025ef8efe5d85ec69bea70cbfd018e9911371e92ca7680ee46a0152a9990c60dbe3414cdb76a07ed847233ff9433b5c68b9ec063670c45c394670313b5ec4304f790cb33f7cee6c1d409;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ae9ee19e033904b0331999ecc7cf8865640896bdb78acde04bb54778b8d0bd7a513b29402491083f366fe435245ee3d2b3b137f974914ca92cb080c385ae0dcdbad98d38754e2f0ffb7967df87ec2801ec99afdb421e105e682f63d334cd087ea8531cc5edfeaf117;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1d460b926f0566630dd22308f4facaf0d37eb19da316f1646dade416eb60d02ed555b2f8be269a37a7acfa9c9cbe334b0642d4878752925a6d357b5ef033c963a4cab8c250cee1bc6f7811b6cfcd41316aaa423743a45256f6c03c1d89ab6d627135424ceb4ca283a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11edab633316978bbeac10d569eb09459a1096ed2b91779b490f8606c90dfb724ee9b3ba0640281dd40fe4f26c1c40f70ab9bcb60e0d1774eb1f7cd061bbe5f88df861e96d3d94cae38367cfd27998a91b8a1b1b9eeb9924c8d9470499ddcee985728f47b2a7ed0b349;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125c06605e9e063e827bef4eaf4f642c7c90809ef472358a5db50cd07899c7e85c16f9c757900edc51b7208931a3086b59f665094d7beb8308e70545df0399637b671ec0a67be609416e9feb9dcec4342e387fa410d2ae00a0c1c74eb5646a9957cb2b0c8e1c9ea3e3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16eb1c319a2be32c6577dfb54a419acc1972ff29e75a93f5e376dc0d6f38d8ccd9da3e94ecf33e92295ee5cee32774a6fd62bd6381a9a759e8524dc333262a1b0871f1a783471b2336cf43f6885b6063f704d62f05c624388089fa2a757dcac60ff5a168bafd3df118b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a13ee12cdba372d7577fa7b2f3b385b2acae6c43bf21da94d66afd897c4a5de333806d51aedb33430da2e184a17eaa18388e53c46f7a2aef78a98089e34e6b5e9218028023b2abd882912e071159908c49f77540a07e4f85ff73c9a39fc44de33ce39e33ca3d71ee1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16cc18205a58984880045eb0e38198f2173f1b06ce3aff43dd913a6a4905f171327c8186c48559b844cd2f1107cdf7262fc547ae2c50d02874f166a1c89df69e766a27d11571cf15eb851b9074a92d4831e9c6d2a3f5da98b202fb3562bf5e99c3339f00ce667f2e3f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h441dbda1a21255e2fee1fd65e983d0094050b9404ddde397664e90c35fc927db4b425b6604936dfcc918faff1b916c449312b604c734b3f5e86d18cd58265631229a76eaa3305c6f6d0ab841a86d5309678093e60366d585c5e16f264b516b5e78375f552b7c1d1d9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4035d499078a653dfb19f2c10a3b85814596ce2b330ce92b06a51232e3fe4ad22d4049b5ca3e495248ad7adb6e485bc6e039140e34f2dd9bdb47106b9626704dd845ed5eef7bf54073d36e1028b3f6aee119d5feac08327e2d7e499c0da282f2aa1424dde68c878520;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0bc955942a68447915a26ba42b3e57f7c4aa0197c9192d7344baeeeb7437a54cb5014dfff1e97220f21e612a46ee80d65b81e7ab9527a698ce92b3232dffae6331e744fb70bbafdb5b264121f2ec8a94ce709a4ee097f08c197fca877813ddbd07a0d4ab9da7b5b7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68fd2b4746c42e665263ea3eb736e73339f16074453974d654fd3c48eeed8b7d07366aa4fa77fcc430e8899a61949fff2b9473504b6ecaf818ac3f6a574892ad87a634bdb376cee186c42cafc3765e2149788691cd01fa0ee4ed19f18632251afece9eb7cfd0ad8f6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b628ab46bd90e8b88afea82cfee08454f7c5b09235ffc47ef4f6e3efbba361d5cf0c30fb7db0009cf28855dc77e202a8e72dd7379e57e42b20587e7af2da67a6bc83c2376be1b5f0ee874e09b9b3cb87963e32adfba65c1c3ce9f98b51822357dada9b94ce66efe77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f4f6622294b4b6d37b8ca7bbe3f78bf39157cbb45470bfd819e72fa81bc7ba9d0d40b3a6f4d886c92638549f9eca084e7a78b2d90ec7a86dc05a985b9a4466b6e827bf99e3f28f78ca95ff36a246869a9cceac6b7c9061a5d5ede8e953f428ba9fbb5510c7dcca082;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1906387188161b8f8ccfdee8ecc90a0463442c4267a22bef30ac858e0180553d7248254ba3c49780e2acefa122535e267923248433381d1c06ce8c89aaa65f7cbccf2a446a78b7b8c687f1e09ab96b4d23805c700351b4319adb1c7b8fcac632c974b899503b73a11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d885ea7fdf33b98d41cd2d3099083ccb82210f2f0970010d650096a1c0ca3548cb11369f5354e9693dfa49533de4c69af4092976e8e3c33402fb640bdbdef8915aca262a86605bea960bd53b221babea529759e6c3d413409cc5a302fe392e382b1f9abf48bedad6c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7749967038a2fab029b50cc34c9ab474df97d59376ffef5fd66ab7006f2ca90fbd97df42c37bcef0b29f4309bba3dab5f76c53a65e0d5ccd4c9338339d05708675f473507b72d5d7e2fa01ece84d2878dee25eb62f36dd36f256d47ad215b4cf52735f653d2abc4d4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166d64c58af3ae54bae4a3679b4e46d49f2add2eb949a30a3238711908c2d7c9cc8e847993fffe806c8ecb701296bc43cb06d2b145776dec2e54544afc2f988c293bb52f176b7db25791224b0d561df4636ed0ae8f5a2d25035dfd80a8cb200017863248a726ff9db62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118d8d4907b5c7664ecbef25f56378886a1aaeda1aa321f68ad539ca9d1dd359dc99bc2123d512e44d32efd9a9926186c169ac7e3a09bf25dcffe77bf05bfd027d76a4e34071dd41b8dae58c558d0cbf34bb7b912f4c5fbd35a520eaea94a45bd0f126a4dc2dec8415b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1bbdc1223b7d75c1711ad191c3645bb5c8b1c16c1a41db746319699ee354d77434a8868b28704d2649cbb66d0c66cae666d17f9dc128d4e7612e0c5fd266a15d6e711c775f83251d8d3b1de88c64543b7b5a5a423ca21d980356ae3f4c92100b163e64839a1671dc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1f7e2f3263f2298f190ccfd9524c8a26dd99751ed7a3fc53e2543a5861d4230a24ae0b05c35ca0b513de31f3fcfdf2ce1f89d2223bff7a1a485042160886ad4a7f32e2200226ebecf66737971508d0d7f68ffb5581058fd70cce17161f2a75cc317ec1d938d4930da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56f68d6c684c4a939c561245feb6c3931c2e8f8b9cdd6ae45bd09b80399b09d0b212d0894ffa66e2ce463c2f3c86fefe05e31de32e9c28e4c930d90477061059dda8f4819d0cf69c4ec79812b4fa221e8f648b79e94ef78688a1096380b8417bd382f6bf3889b71aba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0383f7e555997e6b1a82345c05203dc95cec533e86bd2913aaae031ca2a88e6d793573efb4eeabb330242081de0717add16e099a017880c9e97ad907299b957bb704653eba82a1d6894fc049fb4ab194cec0df9a19850ccb3220d0153307a439ba38a045a84728ea5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0318ebd6abc57cd16a2098603ac710c9fcf9c804f8f307e03b3e49fe48ae2f555cfe397e0522a2ee0fb14305fd997e6cd3d3d2135c6714854e96bee1ef472c4c297a30844cbc6dfd1c04f43d23af85e8614671fc023b3c4a3465cf7c570e1307c47b925173433596b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba6383e77abe8f0485ee673b7f1a5f2a6d31d25d9f2122da02db1d74f21e386e563f75d0cd89f6975d7a9ccc0aa3890c900424db826993ef936f770ecd6454dbd665f997a376c268f4b45b06e8e6422b80cacd6002618a7afda25d4d082ce90de399d48a325cdc55ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f48181fd2a7cf9937d63a7652fc1b27964fd92d475befc9a37c64fddda1eb748448658876a89bd636e5d447e4a67d61694ea066969b1b7d1e6fa924c0f81cb79656bdb55083f1f0b85e3cf9e027298ecd19311d4902d79b6b6441bc3399e95fb14311c1162f20f18d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1753b493d1b224dc3d62d4109213875f214db3278ee9d41b9b72072c04d3107cf895f5db69523ddcb8cce65e5404e846e5d3eabce8f7f36e20d6edc1d8d69e1831c936b5ef9065f9dc1b873795aac36711e42f0127300fab35cd45e3fc8e05da136e289489a444b3917;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1428708f6cb6398dd02a554c721b143c6200a57ca5375412a85320795849ac03ddc3d65157f40f45032d995a1f65dbb179209b01557926297f9dedd537a4b8c4c5f4abf2a337e0a305b4387f396ea78d291b18d09d01e7b956a2c816f1011b32ee86bdf7b1b1456c6ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155dbef2021aa3935596eae32f5654a0e50312df9046e3dec128476d45e47a76252167001423fa547bd1597d5514e4ee7560797fe9a0255e64d395466d0f6be4bd49c98594832e24be35bbf725c19d5d4cf9c06d5930bb719c3b2262e6981a6e77d867c8848932a0b1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c60c291747f240cc51bf67775c65b11dc4fa0af776c404b69d8cbb7f10cc7e75db55c57d260a1eed302887b56aab2cf6cef6d2454ab9ec0745041510d1e165fde1086915586d4de246c1bb6ea787ad715b0aac6c77dede9fd5ce92af77e48e9b4e562f03b8a83e583;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170cc011f9bf02ee43db855ffa84eea42933ee3993824816eda2a21b9c5ad00901504afc0e34ba62b5a39ae236176824f531f509c33bb588fdbc447ca06e69d772ddf34b873aef8095bb900de0d6e312dea9e9ef4c99ed39dcd7f0212761a993b17f9ce2070ec9be06e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a79bca99bd7886e8e3265938e9059661485d6c3fac840af98d27e0d73a9a6cc8d106fe775fe0e786b363112032a48d06af1b75b02a00124ae8ec15ae50e3ebd60923980ffee3b127374ce7b7636003ce09fe2afb8c45cebec1c3db83b1afa1f571f8738dad0a05eb0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147da3fdd91e5f69c0f78c079333d0c0c8493a622318eccb07fa714945bc15226a927315491b74afd09ee131c2b163ebbbb63187b274db451da766e058ca7b9c7c0841e255218b74bd784b996b21dcba3463dda2bec9490cc4153ead37c241dc5def54acbc1d266f7d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he732c23e329727ec75c51f4ab028be578c78e56d9205186f7301b64927d5efd6747a6cf4c7c7b84a58b519d0b500e2dbd61fd6327dffa82f1427e365081917853dece6a062161cc2084c779ddc025671d8b8fc36675d2700b65e5757c3605bba1be226dacc9d13432d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e527048afdb2b56f1b41862e99b201a709e0226c8fbbceb77b9587a4fafd741c0072da8d6a7224d9c86326fc6caf5a84b06e0ec5f348760aaf07829130266b2302aff4f5198ef7ff85690d98dfd3741b113c27fabcd36bb4b6522beea9bc26cb856f85f695acb1fa9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6f3347bd09f9fb511b45985e608c5bc5f62b5b45f03c5bf77ec833b20b33dca0a885cbe3b468577de90b0799ec87cb215c4c1832f6026537ad902090134277db7237387a89d8b8fe4a4dfbd060c6be5654971852af11bdee0d11cfccca7824bc43f445692169d4ffe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56ad3057f330ac0ce39bd03b1a763d51cc3db02bde8badfdff5c1edc49a959a017719d66ee152d008ec42441f831219e71b1f9224190409bd82f4fecc94eec1d618c0e2908ffa0d5734a18042e1280a52ff6d04131e3deb2fe142d34eeaac905c6cd4cf3696f19a11f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3c017540d7f96ef5485f3211cf8231878628a2fb23fdaf99943abe1f07057034aade9d747e80fb499bf921118d1ec216230779dcc31abd5f6be62371e638ee204cb52c8f5f00c36182fe355d1c815727a1a7b76849494481cb88149a7ac407b4d270673ebca1e6bfa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a05cdd6d51ef3ebc46eddd5a2ef7085f2f6a234a4cd2e5d0c7cc68f0d5e8c46594377b51f8714c58716e60aeb9b357407e03b42598c701c0729beadfade482a6a3ac01c3ec3513a982473e483f9786e8d38de84d3a2b54ac7caf12a47c1b8ca3add0b934f1978e1d47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10635cad039cb4f0fed8bb10250e2ada2eef5501cffc633fd985c273956d2b258e33d9060b19c471d742d1f4a0208b3864d771a5985aa9ca4c8628d60b1d393a3fb1c78c541cb8afcf0e6465e90d9a129dac7db1248b08f9e1ea647ee5fcdd168b925cb5ab0e9191ef4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1194c03e58598f75ace6ff0b835ed909105412b75a88c3c112861be8dcbbe11e861eeebc82efe6edc5648b3f373ca61a1d8f0575ad9d66cd61ddeaf36f507a12f61f19c8bc8e80078b10e38633a6cfc9a7b5490d4d44b2c3dbb4eb3632ad48f8d898d0e09d81419d163;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1201913f21e2242f6802f75a7fd7c865d31bb49201a7e39636efc5e12f2f71be97cf6991856703b63848494c019921b2355b6150f8fa8d7fdeecf21c7ecc1aae6f17bfab98907d3137c08a4cf3663d5e59a1674be5fa42e54a8a1cf68c05024cbed192090dacc621b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1805c447299198e59418533dadd1151425895be3fedac90fe45b93c7119105d38cc0f5aa55e754ce9c452815c31f264cd5bf3f831056364479bb1b9598edb66bc6d43dca00348605b78f21fd8699badfa7c115c8d5c59b56dc2fa2d610e52c6ea3354778041bbb074e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccebf84d5194e32f74c065418d745c60c9bfef2589476084bf594dc45d8748e0006c5470e9aae77f6c3fa2cadf4063948373189bd2fe43c467a9d5a08d9a288ceaaa69981983c9f58c28b28ee6855ea5a7ceb48c8544e133a1d866350d7c1759254f6844c8278cb42;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0420b2119380fd802b05448cc6dc90d582c6b04ec51e9c3ff2bee577bb96183d9d767d9e85e6359778881285549123ab266e3f1676eea38b24d05e19a6b8c756a307106e1933379ff51b5f3628f505baccf0b7c6bb951b4b47dbab7cb4167d9fb9d13d725e84a7a89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h256a26febb5a067398d09ffb042da6025657597f0b295b58cd531a8caea18b5952768b7ada7f816a3fb50825b48c2229ec02e9e1a7366aaafdc964c590ee191c0f6967ecbed6079d0213c1a147961cf33d751bd87396697ca96389597048636350d2b29014caefede;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f36b63ef788986415aa6b703137425f7ab31eb660da4a79d3d3679863018bc1f32876ecd38806b9c3ca7c35e17a2b739d8001ae0d0f235c5440d0dac46864be4c88307e0b8e445b923c5a6400dcbe2cb9f976bac08e4d6c1445f088c7fbbed51c3b7279cc2378b5a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h278b5fec65d42d8cd5eab71d08ae957772f32627d93c1fb6b623ea13e175d16f2090fb94066d55931d92b8b494291e6940f56171a0d4e49793fa768daa88dc9139ca7e43697e1d7d4a13ad49f9ed4ae37218427c368d2dcfb4c5433b55c6bbef00bde97d88e94780b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11de2e9931349db1642c6ca4f1c760b27eb6ed353a0aee694a903d2985baa6654789d0961dfbfb5a278fb1dacae92bd53c191072975af62f5c7e15e9f2015b3f35d8195af602cb715fc88e8bd984a7dcb0ed4e9dd3526ea857ed63883c95dd1565e6f32ae6771ad63d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34bc262b9f93efc805648e6399d859632ef9d9885a5b00e564ef631d8513e6d1525d232f4e488a2810512a97cebea3ef367311e836615afc02303a99f3705631bdae02236232b6f1b25bdbf5c9afc22afbc2d1a752597b415db7929ba51de1a06409df3dcda8a61a52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e57ce8763e17200ac4f554e3395e021c7e1824b76039763a222032245108bc5db1c4ff2403662b5de8d52c551c2957a11414245009dbceb80897bea6eeec097a548f8cb3c50b573352c4eeada5f0a0458b10474a09fe8620c3f66c9d1bc5f73597ad26a9bcf5c7cbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1749fa13a191443a8f231a56bc908a1f9957961c78eef5a490ce88d9f2ced6c8727540bcecd3717b9302827e0314396e4dbf2107c51c1faa2b73fc4659fcda37ade3272f9be2ca745cb735766e4cb93e1c5823bd115c4fc8aa755ec43adb92370857447fc024580c8eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5c159f51b341d80ed80cbdf4278e9852957477aeb999491498f59ee462a96af9a0745e8506ad5f4decf8ee1e290143bab1b07ed6c9e36ca1382d275d4a14ab876fd2ae9b398312918f2454382ac6fcf3ac25bc58e7480efc131eb8048e115f818b60e0d5df49d14e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42b4e96f9c239fb642651ae00e80d1816ffac2cc429aa96a032d4429e7de31ebc099e1afae9e79dc8056c5f6e66a835a467f93391ffb3da318d05ccd1b24e23a1fbe0fd5963abd7f5fd30a3f6a2a54820e0b5eba29f313df769ab655d2b1a3340f6ed2b7af9b56a794;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3518d1aebd0a740a0d8a0d4b8bbe038c3ed992b923d7903ae1b1d66689fbfcacfb3c5b0ab676afa57442a980016fafd35d0c66c9c5bf746b612fff6f6ba707df7bf6de6177e379f8e9879959f4ab38ff78bf5c68c2b9efdac37ab59a6a944f5f2ae2a4f5f8e7ba1a59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3f5a56badd0210bfa8a0a33ae180592e9960c07fea731b499dee8e8b8ee3064ddb6031b1947f20ea498bcaa03c4cc39cbad469bd08b0252819803ec58792780a10b80ce65e42f111e9c55941e615ed39eaafed019aa952dd48e9dc13efd54ecc50812f992c012c11a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12738c7daa02eb1658b86a09015a481d99c4dc8ff826b8a54e71c841404acf63d2c5292114ef578750175a46c987629ecd98555ec804f68e6d6025e9a715250865dfdd7ab939b5c2e87199edce025b2093b964c83c346543cd1965ed49ce04d06a200ce16eddf517f68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75d92df7a2f669a6d3c7dc7fc9afcfdfb9160d05a7bd48f79f7b37459a43586c18b91907e028a25c3a40163f4814e5d312a8e5c6da70ac5671adc79885119fa5b5fcd5092a069355ab1921b9a0bf1fde6e843eea258973d63b57ab7f0f2a968b40d4d7f59a623143dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1223e0c82a8ba27bcc33e8754e53e2e19c0a4b8819af2b04652f1b148aefb00c974ecdb30b70e5f11a299b3ffbc72eb13de5c227cc2470447ccc96e0a09544a4f1f4f947be44ad7da67d273e3f1226babc99f95f4acec7c25c6ffc7751dd62f68f705d7fe1215f50d49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6471e648bfcb14fec57eb37b7a7e6607d60ca2be755d86270f5fae5d5ce74fde35005e8b36d69e40bc426fdb99b168179f63b4aa6d23c979468c02647f8c6973a8e94e16735b3e37d57a11b30bae31b208d3ae263c1d0731d0f6c59a3ae68bd06888a718a3eac49088;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb4b1b2105dd5136ef2866dc00b9834b59a31db6f11562ed4b0dcbff77d0f8b87ca530056aae2b6b0278e1723f0bab23a88576d5e202bcc163886b39f8c149d643dc0218dc469101c631510cc23a5343125cce01b4c4f71e6fb4b175d9ced0771f6c0a975ebc147980;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118ffc3e7290a94aa831b303164e384292d2f49bfd3c744dc810fc121272e3b5c3953a9523d08215aa828b8ddb4cc2d8df0233d33bb50cf800ab03b25e8f1f9cb2b0540d235f41edbcd4aeb01fba13446c04dab88d094448e4427b74c757f7d8cb14f2f4d1ba0e40ab8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d8e7708824d7b3a9fa31bf022e4cf6fcee85fc02ffc3d5668449a1dce17de653f21054def86f60e508d87f5530afbb2acf9ce9be6d1d64cbe3037f9ec85d323c182b4bebd83b62d3590722646d784b7e815772a1d734798720dbc08817d24eaa9500b441daf1d8dfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e150feec5413e1245a1edc1e3fd2fa9e4b8ed91cac7d61831a973bafb9dfdcb984f55c5abdc79c5fae86af97792f958c094f07f4faf5eae12e4e512f5d463b4cdea43e6b1eba93bb93c0ccacfaded499502bc3600f82a08c83502673e78185f1376b9b52ccc296ef2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8165ab51e5dcddecd103af2f2d608393ebcf8c42a3cf906f9241eb7b00fc59c639727778af91cc5eb5693f4a93ac09b230bb976366ca36ac8fdee4d35ccbb8f8c9e1d7d41d08b22720ab50dbe003e797047b9662a0db633246ac3a0a16f7a195bcf9a58f4d2221d6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c2aa6262e6269cff0c49889a9c6f5e41672cfa15fcf202a56787149fffc17c9ba05b9d36446c8e286e042523cc828352a69337cd3bf8b0728c0f4a0f5dbb2a17f032061a55f23d544a9c9485f5a03a8b5c92abeaaa9bdd0e03addfc6902b25b80919688b31e62da5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb9cbe7153496b665a69840d50372ef354d5f8166d9529f6c4d3085ea990a8a564fc4c78c1631281b192176da38f96ff4a9669bc5cbe4897c65e7c449f524333a1f70fbc7e218791c5a7349f2ee5fb3c361b93dffe4cf9e05f3f39eb2d4212b603d40b7faaae87920c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54f281345d93dabe6838ed74c46b86c8e3e9a24800e4ab1057804e4b3675e05a7c84fbf00e9d6e52967d4b3803b265962c48ae2c34bda9c3ee14ea5fff75def6f7ebfa3f29b16264443b16ec944740af86a039ded0177869fe981dd4d50310f383c6181b9fe72838b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10672aeb9279a1483079aa3c1521671f63f941f9229c55b800eab9888029c1ee1fb8a6ac42b26907fc40bfa35f739aeeb4a4c4f47494cb4cf5f582f43c11a0c97a38d89e9f949864e72c658241f9c34fcac77200539a755465cfcfd175c8d8e7e7f4acc3e12be58875b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52187b41962e982cea5e821c082d95207cc94d02ff307a5940544d281d80f9d4ae561d8cf034fa9a5c74544fd65d77c6b99032c6c5baba4f769ea27dfa6995f9711977d1524ffae5caa908f9140379d8ea63adf402bc905c1f1e4ffe44708743fae13cfd1dcff7d6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142de655e51de405e4578d0ce9fdc03f0af717dbf6baebd751c9fe95c879d67b3df11281198e04e55b7f59c1a857c420a4f360285a366c84460eb8c2e0e1199c21fcf5e1460fbb6cb69b6075f4a1a3463ff23db69ddfb3b3c0bf75804d8d32b1467b80d2c2dc62351a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h49b28b5ef8415ce453eea717517d4d5c36bf8cc45cece61ee9b557c2edaec3b08298c3aaada72d0284fe9985c7c63770f2effea666daf54b39ba916637aa3033f164bbc2bc50c59183f154485bf2fdfdd1bc7897f413ffc89af64bb8ad64bb1ef2d1547d90be034038;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42c0cb146c5385177cfc155fd1fb6e59986e2544ae6616fd2cf4b6e657f6d3699f63a21b6634b2effd75bf01bb22deee64c16eef56afd2d5e96f852d067152fbf4051dd153ffce1ecef0f1618b2c758c9db3245762a90f2edfb3d769fbf59725ddc3c8db82ed41009f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2560b854938dc0ef8305ea2e1e84e37d6a1d4f0d2a4bff86654e488b85e923b5a8ea4e92e9af037e35f583d456e1957ad50a2dca5677835cf34f9dd52e403127288a4026853d1480ec8ba12a0a1844f1a4d8fac4f7e3f9b025dd4585f3c06fe917210295bddeb11b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f67d8e5dc76e15572954adc7ea100cc1aa83bd3bbcb6ee815e1f54a8b735db5613bbbb982a1c7d58703d0b398b8bfdb0f2cde16da2dca47328a27af20c02d0a910f654badd49f6e2cee4014ef734b6a6359efd312af3a97bc87c9fa324c466132557aec63b6a0a6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e9941dcdbee0a48da913ff491ed2189d395ba96555eb379324469b512ac560c17d4f090e512c44768cdeea4a94f109ab76f4331e0bfe9b82f03dbfc1c8c08d475a002261e460c111f83b2110b64fb9281776c9348295d3199d3d9d7c4bed80975c8f692b8c331a544;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155065bb9aa64830d9da0e403f9abb22c9a380de452c494b6dbc62e4553153d06b1b6b231f363888795060a2b92f95d63bfadc90d6c6c368532bfcc30487382d3c94a5bf0679512ae2e272a7b892d1c92acdae494685488610810b82b953ce189ef34bc402776c1da67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba703161bdeb482f39a730857bf3ee0d95dec7d05963521d06f6c5233ea05a4907a356ef107828d143f4f7569024ba806e3e8b3fc05acaab22c6e7c0d9e61c22efd98962a823e8f5719330ccfb48f1bb6cdbfb760d806cb5b8a700290a8961242ec498b20eeef3fbac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bce0a0ea3e66441c3041a6ffe9c7e41b8473b809f80895e4d4f1059e7e620bf8258d81f0b014a665dffe6c63551d131d4dcb8748736b81877209a3eb6fd961359fe3346cd1b15c32295dc79ce9653c09ac273961440d3e9e6944a48362e654e1b3d9d2d5a65d727ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ca6f0898f1919d11892a5039efcc03e296b84753fbf7e0a7775f64c4b7209acfb58759e8c629ffa2baf6bbb940fdb65007aeb58818a6d5f8433245190288fc209aad82c2fb6c579cc9479e457e52dc76f54aa8212913fe0d5c9de60e682cba2ceb7858f954c32346d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1201ac4352ec5ebef2a9bfd06cb7934e226176e65b9a5f410f4350fe71b97ceed9b85d4060c9bc97ea35b8f8f6e72b30c62b38692ead11fb8ce8eb6a4873f8fb81a61d27d327e9d9c26cf16266a87b164f30109cac11574d5046d25a151f5795f7a807f7105c2f713ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fecef259d2bbad16c7526dde7e59cb523aacafde0006424b4b2a0e647d0e4b8bfeb9984b9dc0839bf2fbe0bc2786006888bb68548b0224609236d9348b2b42f7d9801ead9d7ebfcdde64efa745c36c8d256156431c5805358618eaf48d0665837d114b228a91d2fc48;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17296cc9d906842f8aeda2b92ebc5741764209c1bbaae8c5527dce69df17ddabe28c22f5866dba18442bd15a0c9f7055be3eacb50d6750e6e1d5ed00b975b81426cbdfae4302a842cb91debd2c8942b62d117112d40a0e9309ec334962c17ff14e16b75c86b378e4549;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f730bc20addef20e13a29dab8b181d7ff17c37dca32452ebb0cad9939758482fbfa3631537af1061df08e1260eee937ebce267eab61884740f22168b7d2c851fea54e55f5abe16d46880e2e6c012bca17abd5aa3e7cf67508225b6dd9aabc0206762924c106fa55e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1611044792242bb97a0530bb8582a3799d8ddb4672cbbe0e64dc562599d3995380b0e2037c3a9a2d290e02ea71caa0145f7e816421c971c0d1d6a493e757ad81f55294c984ae3895cd1cc914461d5d927d1c4e484f480211bba29d771630e7537c204248fc049385378;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aff72d6960dbb3910b78dbf48242daade48f82003d2f61fc1f9fad15bfffa53ee7dabb279aa8847eb0515e84be4cd2914dbfe8d8eaa445e14b3723b1bd09aae1aee67bf7691b886ac9e2c796464b908046db336e42f48121ae1d9134217b57768e164b435432e35851;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1aab036585734a7cb9cd6193c62efe616b2ecd6f150e84d07bdb287f27f01571dbf13c234bb6edd6cc7eb8f0448541765fa3a2057c09690c8e4f0b5c0a82aeef808e055e3bd5453c17db270ecec04f307eee1ce61f6195d34f5b0f56046407edeefa06a3c8394dcad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bea4a3dbfe77f9b27d23e020ca42efbc36202701dd3360beecb05c9e803621e7073c40e036d05615a779a1e4702233b6b5edad51e7ff2e8e00a699a2d3fdee80e9ee2fa2389e208dae29b9f11fd817e64614845b0829442cd8bc7ce01f0a5af6b7852632183de1daa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h699cf47da87f7120a40df50c3727f4424a1ba613bbd5b8be9e726dc3a704511f3b5495a5b559669b247f46a985046a584ab64089cb7509f8b95899b7140217d1ca83734682f3de325fc96c304f90754309aef620759ff788efd9c699f0eadc471f38bff435a16d7b53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf380ab913fe42f5f3f7da3f6444bb2d195ef4c891734c68a862184ad8471e0001306ba1f1c6a3ef8a2c3b2541a82478fe8d1d5c9c0bf278909f0c28e9af7094788de3d0109b9c2f019870ff1a16813c0cd3eafb5d98ab37ac5a8d2d84f47fcb1eb7f4265b4d114012;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0a4bee3051210b56154bd208d0ef3e34d780cc9a2a02e9ac8ed7e3888debad4782d4bc13fc30404e166b87ae5dc031708dee454f7b908ef38584cf490943190a5032e3eef08b99726ae4ab7c068a9d5131c9f5b23f3d2991add1666c42f7ad85811d0bf4057b1e284;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h726e57e59dc4d6070a369a09b44baafe91436ac5880e97d091f810bdcfae36af4ab37be85853cc7106d3ceea7e44bbeb86594e005e8a27e1bc2a1b264b52b9bf61bda5335f57322e10738161b3b10d1e28edc8e6f7bee33a39db8c4d4ee68dcbdf67e238ee3714d012;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he62a6e6d0446e669da77498b98f7f8be5f45c81da9557260356c35c9bdb60dd4255c35583cad3257a5b0e69fda5be2463390aa05d189f25326e068df1d2db7351d2655cf5d40be5c1a1e528c3423568ae5c7b55f81cf76629f57e9610ddf8446dc8e54fd23cca76585;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb35f6be4c92612aa344c6d4a7fb3fd3532905ac63fbfcf7e2033af750f90c4a5c86e494fbcab9f1aca5ceaab3d9cb09bccba50e991ce72d2bc6ff3a7dd70b655e1de05f3d883a907ca75d0a777793e2276a0a88a324547337ad5853ae027e6d34f7c2eae69cbb74bcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d805ef1b82caaece7f03cf8fcfb1718c7758dd3a9dc7edea78b9660192e1fa545d7bb809a4df4d8b1012d87274541cafa16cc3c1394329e6a9cca9c6133157a7f870c33826ff00011a9949d47539f1734915ccda9f4beacc912dcdcf7278e9b7a9fe8162c0c7badef5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11291223d7b32ded79cb790fb234caa99334bd31a26e9f21d04632751937ca897c43e6b9ab76761dbfef053ad8c61d1f61841258105fdfb7348af386409e2fbb9dacc17640d46f4f7c7ec18eb459ee752273a299da7945d572144ac9267ebe6785c5a1bd93ce53a02bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16969e35455b86980bc41373c44631ccdfc43bc7c018686674f3d7ed7d3e387c29eebde2c8540e7785ae8c200574f753cb1283c8e4313b538f7892d362655ecc2e0123de9124f2ae286058391fa3a43a99f13d5275fc2547d040846abda2c76f0b0a53b0679679979ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14713cdae08c0b9b6690371010fa008028c385e90c219a0f627547bedca741784dd75d3d42593bbcd8ebbb6a81159b37044411dee2ecdba800a7e1e77de7d4c3ff72ecf321b2d151c6de317ec66dfc681fbc614ee073b350aba626bf39daa92cc201ceee141f3648be4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3eb4606a85514f438ee242e1a6f6a57d120a07a4dd81f05e52e7ad8367a6b86a988a44ad1ffea39b70299539bcf85b788e7fd6348017ba0c8ffb29b5ee7ab9089c6da63bca15f8d8313169cb9559e68cab54f029e6df79e859df74c0fd5718fa7e0124198e02d432e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2688deabe9c3684009df070d5374c672f8730e7ea171cb8e3d7cb7be38d8927ba497724841fb74c36313a01e2bfd405622644b11fa99c5ef19ff8650e9e93b97cd9a3a709732c3c0dcff45b0605d2e2e2ce615f99fd844a1cef3c43c54ba5ea643e1c6590fdbae7e37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e2456d4c1cebbfba30bfa221bd58bcd73ab504a8b0c5b124535963326ab06163d01cc2738162a965b3b9935c0f8e8b66f401d0290867d7f4610a6492d7128e3d93e693baa01ad2e96afbed33b8a9194b70cc6ffb09a65daa1a039d84ee67d4d5a7c4ebebdb92cc467;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc268c202d48860436f156f63bf796a25090e5032f8e72f3acd012a3b84053b753b227ff59e498b5ce2a645472033d1db88240a37c9245282b96aae80e64e6d4a89b350736e26c2544cdba91d95dfb852bc7b8e8d541e6ce364cb21c9dfa68f1bd02c0f178f51a66f5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1095330e89a96bd899d642fff42c662c7d290bde36009b73278c3c9897b39c91e9f584e5f735c262f95f8fc680b4a6836db2bb0ec0f307384ac609a0924caceb5655b43764224f8fbc544863f70a7461c96c4340e073ad31ac527d87160395d79edb17cd5e7aa817b1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14970df7e75f40d5d14d988106622a1ac0357eb328dbad6d69ddb2bae81a2df878e11025470a4c9354c64d0b17f4af148ca8dab5603689057d672f9011e23df23814bef76bd2473f4a44104094e4c5bc3da6be7a305f0f0ff87ea6131d2be66a302690e74d9682944f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89503de051f8a63eef33d62ae42a781361b003f786b9271a441afb1e6e5bb11f3f18c0b74975948dce5055740d039c5aee2995927cc24bb3a553fa6dc61184aa2f4fe4f031c9d603c51ffaedd5d63a15ed23d4b9b671ce2ddf4cc749e0b244fc4fea4eed353731a44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea252d3e95bf5c96caa2e8fda696a88434893c358722bd407a1c83cae37b3eef74d35ef031801ac46fa22810808960b498b4d6958850350784f6cf0bc5af02327a957e78b0b8feecf9fbf5b81ee2aa53531c05878161edca8b747e43289345d5ce51ca88d290de7441;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f33bd23653eb30cdb6114ca64c8b321f73b1925fa95020ee7c32b8f9caef175ff30ec9a46de4eadf4b4fb280ef441cbf497d9bf1250d6846faa684b612ef21dc97bf89fb82bace9f7c63e20da23dd5190206624dc92340e91af64011e8f21333bf5da5a234e7be9672;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5dbca114e4c4cb13dfa8290d1a02607eb7ebb284fe87b7915f613e38b6706f0dcfd52d648717ca9a4470f1a137cf77ec764c68695c4a8cdc83aca72b6c4c0eab9cd968fa084a709877f1a9a7f2197a2f13b81dd836a9e8d489895afb0556b292adfcbf6d485cc6cdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6817ad09e28e65f7f5e84c5b87019333be235764a736bd60a374d2f699707e69aa6b2349de574fd5dd0b80840b4b8643121ad450a4d3bfb6691310b491c191725c496ae533f544e2842b01860a07226caee1540ee03c77a3fbd5bcd8109f8a86b762d1e12df69f634;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h49779ef81db859281be09c9e0907c40863f62fd4e9f212152c65a561c84fff1bd8b6d2b5390495bc43f3f78caa320f6929f9b0075249d3a828880dae2eaf80817ae835c48eaf5605eaa1d425b90518b26054dd33af275c4c98c90adfe91044ae2d334e00585df9b3c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e19d7ef5127bf1f384f58aadfdc3c3bff6c22e4eb9069b31f66753fdde44e5cd3cab7c55556233d0519a54618d85aac3ecf360e310e8a65fced488a144202ad1f62e55381d8ebd746255b508646f9ff5524c5deb025c377236fe8e419fbed6d3abe45608ee6f8aa651;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae4662f1df367b305177a68d7283e48b72cf9cd56c6dd5fa85fbb2875f078626ddf70b3a22d107572d40c15161fa28e739ab898e494f820acc7b944db443d0d681fd7f43cbd99e891e48832c0128bd3ffd6e125bdbb5f39b7d13289719ebee04de00c599f782b79ea8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h721c6cee379b7187410db19f6efe04910818883ccac00040ef2a2006af101dca8890994375df20ebbe03701f7dda45d7b195cdf99cc9be9ffd05573eb0325117c939534b61fce2009fa085482965e211d9ef2e1eb2460dbc98a082822ea30b98a3ca0b5e4309711de2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31ec27488ea3e6af2bc57bcc2c7fd4fbdb266e3f8585679ba52beb5875d270001ec6ec71ce63f11c0434dc23c9ae3afb3484c1c30d7bf4241d6ab42ad38c00da5fa1a7fbc1089c3c0229435205b3e4b5bc5029964f97a13865a862cd375bf5c531ad08a454eced93a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112b050348007745509574d686d07c7b63f03110b87f3f2e4d05d772449a05dd660d2a61fffd104a6c0cebf8e7ac9d84e261739998b0dff2a87425b58fc4cea0bef28402e786a74fe22186a1f4a6ba3787f9c57ef9c64fe8dac098d86f4ec6df899842f826f3022f311;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3681cc456ff6374de965e1882cc9ce2f759cd7d2772532e05c9696a4e39684884826e5bf58e37f9be9c0527381af55c9c974334988e9ebcc88da717da899c8cd19786f256311cfe484169c90b70ffa0c8f1a08ce94d5f22f53dec91582d9c605b6c8f018532828a5f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99caf92747f60cb5872881fb956eec13b9b8164dda6ffbe51aca5bce39d47491e52129cce1a3ff8649d4b21cb269eb5ad7b442273b897cb845e97be7cc2fe1043015c691b03f089b00aec4321b8efd3e52ab00e7578a7a3a9b771f056b0412d4f8720a6a650e625871;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5355ff4a1e178df180fd173bb17d2ca14b86da6fb04a48aadfac851b7537648b26d5219009ecfcd809b03e5fb13c31d60e4411d5f50cebcd1ed32a143fe6cf3095b868bf8df627ffefbd3e83af45c513e578c8c1d3f33d7b1b337533b1f1be9d2781711d00e4893e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f460b5e05d2f43e5faa59f4bfdf2800f495c6cae0a86851ab20b1d28ea6fac34d69888f13ca1406720572305470a7900e78cfce019b2f7ca827e1b9b48937c9d4614cf54d8619131b87b77cac6b09a74877f04066ce774e4f5057cf2e5739f830370c5e67b0554e605;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7f5cb97e4cfe0dc84ccb1c8489477429af0492cf9ac00d231306ff8f84c0a2536184b8c304ac40a0bfcbf01b567911a89df8e0c9b36723bec4311e1704b6971339a85de42a65118bdf35b06859f3cc3840d483f701cb0568ddb931ecc66b7eae8beffcf8c11416419;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15dc2eef2309b1503a70d0c4b4c1523227e560eaf1538ac514849bac8c72134624d736e1203f15c1e9847162c4938e90d34224cbb6d6cdcfcad6773012d26e1568e1188a2de801fc0c56a44a26e6e0f17f66011bbd6bb469eb97130dc29c69d5f51b703652789f2d7a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f455cfd88ecc74b077f75caee4f9fb954a70682488fbca05d2b8f316edefce8657d2492f024c3aec4e40cd467e1d32b9da741ddfb1853fcd590dead47bd859c620a5a0c87a525bfd51744b14d0d0395d4bdad2cf554b01c567f1233a61d6be725501ecb04a5aff903;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173c29709b86c354d9e5a066365bb8e3abe62d38657b649510c2ba8cb2257dec94e12ad50abbf0a04d43c1d1feb7271fe72a3657f6c2acff2fec7bdd76089b9e8acb21177dd4995e530ed83fc63ea35a60a4aad711791a9f7f0248560a18d5075e90ee838b20af2a0ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b2379472898f66318f5a13d877bd2161293b2bab9ce017860f3d29f247a66eee5253be32ac98fae445a51011192debc3e57bad9b94c57f8a1f8462085321105041b53f3f79e94341f9d19287a0ee95328331293a63a8c0404a2dcdd977b2326ad2e3f4136421a95ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1538682c86ec7ca0910b72ee2134a6825924b362d7307f76c05eccf29f1044b3a7dddc72ef4ca6bce758678bcfe339332e6dd4b37666fddd00d858ff58bb9f890ceccbc9a5137028b2fd60c9d98c91c6f16cac0a4f20d214e4c47e8752b2c00e9c3611d2b6946e75594;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1696c9f0df522d7ce7477bb71f029311d9a5fec5f3c293e89879b7b0297737ff75a12b9df2da4631d85fa46cb6d020666e7cf449e99640a28d1a389f7e1a431dfd9683747114f083b484d584cfd447f5dde98f7717487093bd5723db21522f09d73c237c389ba23b470;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f8d64489c959763c7d6c687f58198f0acffec1454de79648ec03774cca4ce61f414488c2f13b444f955d2cc237a5e6335106ebba0165fdaee50d1737d3aede938f4a58e00597ca9c6c46a82ac2aca163152c3c8127a1b43e3d456f2f53b942d978568dadda09ce204;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fccaa7e49a20fb218d4a26a119d0251f6b1636e891072a7c2637a48d57305a01999aacc415d154e6f16a703b08b09db193cd3f82f97db5f049c61ada8b477c5b10d065f9a1d9c7b4150e97abc01ef1885413b3a09621eae0c37af450f42a4f865291ba4130a04c842;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h371983919b7a0d38d8cb6541eb177ab1eccbcbe8bb6c4d1156425c52a6f6cc2a262e1e3e2bddb0f3621b4d25287368509b2c45e70e392afc5697d1ab0cbe223600b86dfaa0ab0c1a8c80a5902ea7283dea17fda7cbd7ee22b87df9b99d1395389e79c25473e6e8eaaf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f7e001d1c8b9bbd6b19f7800beb1ee6192ef7c7889772863794ef665bf4d768017f38536176881b4e9197b8ba336ae9ba189f54621c301dc860a580cc22ccc1fc64ec585331ca8cbebd08de75c442bdc2fc1ed1ef405e2b00d347d2ff8f4adbc9af326a5b4c152674;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107c9ceb9eb787f1aaa1523aa9d1f66c00a860668a66692dea6e2c654cb33b38b65ddb21b72111bee5b3f45ba4954383852d1e489bae4402893fd1bf402047ce0f6dd8bda716a7ebe51bb341e23024694e38911ba73b8e92154a161bf7979c9cab65a04476b8d3f9497;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a4ffd536e6a59ee21d25d052bd84063d947c040c7bf7220e03b1c3d48b6de13f20b9630b2ba00c6ca28f0ca2e3e9423ebe292e776d99f31592becf603a2e01fd8ea7f42ff58a2d70ef1bfbc76fc63989000b3d01c489672b51f28f41736b7318778d11577ca4e033;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a948ce5ee4ce4286132e9325bb571d778c524fecf3676c39c7fbf2f7613a861201bab141f4d94bd2e30598f9479bda08ce917b3c43503b0489de73bf1b4bd8371c1960c0124931efa4fac6663e355db8bcc4dbddc0a1b1527e8120f4c1607cfec40f70be3834334f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96bb37d25039bf0342fd0f17fd9ca334f72cdd0d8e200011a28481eee719e76882d364ec5a63d5210bda41b24c8a49548fc5a24612fca05f9452801dbbf9d208580e79f74810fc3b89011f9e94e7ef735cc0d2a2eb2fca010ffa2b5db1ffd4484819bcbd1811217bb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd716f6bf69e1f7b2ebf0b71ac0d8b02b87964fa7df34ec3ee23ad65c0c82a0089dbe1c606e877c3a5765145f82bc51df296e07aabb8e41c821f061f6195909267b4290cfbed9f481ec7c1de39e06cb224c01ed28248a7449eed58979aead8bb037451cc91a854076d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4408fce42256b9a14f9ba42c57833129f7cdef6e7b5f43471f553964b51635c3204c06fcbbb16912f497bbfd6da5e6f0548c2ec8ec832bdc37a3db64680a72f34fe3a6fe4f951c0f64bee9301872b4249db798401f3019ed7504c8fe52cc505e8ef1112321a0adfd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7cc14d87332b9f678aa351626213f3995d079b01246edd0ce5670d6bd5fd8ac2f5a769018b9883fa54e3b0a6ee63d1c0136b4b9f4c50dec7cbdd43416207c40265cf2ca6edc544ab5a8077c14069d3e5606f5f802cd1643804fcb0934efb06bef5b13c8a9ab3e4236;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he76761a081ca6da5b50d7b244edb68305220d36e5c8397b3156ed32e7e18c2e6ced807a94607f35cc2d62c93e84b955b871e3dd7064527a0ece9b3b0a38fac85e232b7b3bace205a139a41aacd35644503bfa1b42340594cd211b329c12a20c49b2a233d3a91547909;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cba9163c27ea3e71d165c1f4e3bb600b3f247f3264ace0df36b19fc6af46d73fba22228de801cf3f3b6649f68c45c2785aac40e7ab863f03ed03b95c553a4f6b034cefab58c061d9a68ae35b9e04ae7cca8b5e7ad06dcddffe1fd345e0d7e31a4d7ae4666928e200e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d535ff4dc8ac59fd3de91f22da7b0ba7cd22122bc91230dbc57436c4657aa238761dc3ce6ced39f5e5506ec6b3382e643ae3e11f76ec74238d7a93c1ab9230b5001d60a072997891e17701255fd27271823aa68adf609780893cef1440b7d7206a0afd21e7c3ac1cf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15bf3bb8ca9865896717de9e061df780d935fbbf85f5dc4d55364295e759b9d2c772746a995777dc515a605fbd3aa7ad1fc2c1168684097901202906a4f7c2e07ffaaa62bf699cbdf4cab02f36bc649a1ef52ef62b6c5b7386eb80aec637b2cc55a724c52fbbff8b6d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h360ed887054e51a97d30c2242cb473485b87707f5b768ea6de71df99824ddd144f59792ce22158865a243dacc653de791dc8de7bc3fce70fe62f325970a91dfeb47186e6bf390c625e13a6724473c02dacd5aa56368beb7a20510b6ea2a84b78c8a9eda9696ad472ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ce5249604d978ceba96bea1dcf549f8c8c620b0bb6dc3474b73ee4ee180ac3b8f0277282d669c4a6913d1bf81ac17ef33c260622e8c5197c647ffdab91bbd7194b87813bb1c985e3110e8f781f1bb11f9cc5da418a1b4be8286a77f92dc50f31091fdfa2e0aabc4c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1812f7a81eb393a13d7070848af19e63a62bd74a019ad89877c683b2a4ea452ec047d5b63a5c918c6d439f3378afe2bce1b04d0af1b9ab8c53ad7430f1355b9e4221ca863afb43fe11da435ae52e227fac8f1f3eece31083ba4f22b0d17592af75342c10f8cb4723d85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51095c0a2243fd8640040dcbe06706d166586ff5b9d5ea7ee9a08e2f3cbc4242fd9cb16f7e29eacd814e896f4bf24cd70c2762019a23654b1225585d206a2cd7097ad4627f8534066739790f25f269a41758f4d042cf747fb836c13da332c7c60da0d06c419c425498;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1375ef890549e944c370dd3a1e94fa4455592ad5a007192286d8eb5edf1b0458689ed1ce220ffa58ee844453cdb954ef837047765213c5a0c524d24ef0e210b7fe331c1d3c0c7a69df14ce78a3ad549793793f913d369897c9740f543bea563d3159260c83c8923416b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eba090275cf91467b409144b26f4af07181326f0ff4428448b0f02e33758e9eb518f4f936bfbbe2249d90c934bf55d7a34c580a43b087c92ed1b2b413238d9f6558ca4aa43cc94fb6c8dbbef7172d193058acda95f2bb5151f269479afa519494cbab6fa3f4a7ebc23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6e54b45d1ce81ebe2c1858fd32b2057c46c6ae5db1aa7a79accd0a268f36776054924a47d6df62e5bddc901e5fc0b6273794171f45c17763b2d24fdf8369261213ce525365dd857396ed19cb5cfd94ef18a81490ce35985e26620552712294f82ccbde663ce01e697;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce8e052ce9c11753980bb4f4c488c5e9446956913ac05ff9f7c810eb855ee6ba11bb3a3bd3d37645c8e568134ddcf106b4072f277611d7194bb28aa3b7be35c02705ce8b75caed930c9e585700189cd9fd2962487b594cf657e31bb31c862d342adbd25aaebe51a0e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8eb324a4861c587b764137c91a859b2b06a44d4f29989e4699e17eb8fcc1f004f3e3d4986bd9da4c1441e7d2654555301fa69235ae3eec8dabc17d6f7361f54a461eda9c9b955d8326ff67d90dd3d64aec9d8caa7c7c13e50c242e15e5f225c91b6b01078d398957e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19de1f1701fddfdaa9c51402f8287aa5f5d3c091a92fbb9b3d90f1e09cdcd701a5fc82625e0ff8dae1b91b42f16312cbf8ac8eef9506009b63875de64c85654f2346809f57af9a1baea59a099c733390a3234e6d1ad905f7884c048fc22bee97091eba749bf118dc1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146a61f73c718987efda1d3fb672a7b2cfb3ab8d0dd380e1800a4799e78a4ec9d05d7d310d4e2e04c1f49c365c403e2f28d62ecaf135bd228fa487df2bce84b24b05baee52faba5b315deb4b14845eb8d5bdc327c210d17b9ff45feab7424a478d25c06a712cc9e1f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9dcc0e765ee95b4c6d2a64e089e9d2415b8ddb14f5c0ff007c703669f2bc49cdbd75fce6714e252d2c6d299e5c48488f97f941a1fab40215a34d9718cd75d51c566b56f86b700b518d60ad47986d58313f1a6cea89070e04d271f456c8cb1566dd8eee22e1ea3c97cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9862951372f675d8f967b6fa10834065d9e6bde603f7c77e9ec4180920ec0b4d85f89fe8c14e1c840bc1f7ca8cc19adba483313eeac08ab2493bc9870c04970da1be2aa3bc6047bc6143e1d7d8dd50db52f15fca3cce9920ddf0db9161df7f6a418fa3a107e55a25d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6bf2e73bfad9da8b6cc7d933728b0625b84edfb97a9ea245ec534472c6408f03499982bda99f84135c4ead4a3c42057d963de266072a951f6f4d6655a4854c4986f480c745e2573ffef00f2086387222d5287082c5a914173f0403c22f4bb36451ad47c5203fa7007;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1858ea0acdc40f91e2a0ed8e15d38ebc10b9a62713ac4046fd0e2abf7b64fa18880d2eaac657e7526803b34eb1417a7ca240649be639ebfbc6de8ec47b74a5d564635fa2a7e16342acb45fdcc6f7bdf3e11581f8173879580cbb0039783ca9839a502e09ae025fd312e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56b3cd1293c94e1e3e890e6f7f69410357a8768c90e811f13d32577c7937963c02bd9985885ddf287760e00dc42a6c58d076b305501ff5976c7db8a33a54a87d4cf409648c20e7a7dc37f9cc955a8317717e5d86868136a9b1bc5561ae98191c8ea381dc815a5fc0b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b145f1fb5f7c5a78839cb47b5c10d800531b247aae9c6bfad7591cfd46766e32b6211395945bb9361b5fe713d6e1259be918e47bafff420dca58926f02e440f29650ebbd7867d93de76d29a3f5c84f42bf19c933881e2a3046044a10db2a8cb5df8b79631c597852dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea677665020db0b2ab6dbbb21d5ccd8cbe34087e02425fcdfe6809b4cffc9f35282fbe03bc19fe783f3b5da3a5d5ce7d2cda3e3f9e63f2b94bbffee49a484eedd2f95f1384c4ae486d3a7b4d30259265cb7ae4f19995773575c4d806056b30fbe40f6bde2435fabd68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60fcbbdec59e49ac4458b84ec4c3ef615dd6c608ff12c1993b464b7637e377a1163501221ca6ecfc0d4905264db4b1e3a686d0ba34c5f8b6999915764adb4bb97eea35308567e93267e24ef31ae5aeb2d41658c7fe79262246c6ef05f1881b6274145f3a69f5f38d65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b50d32e664b94cfbfb0521cd9e31dd0a87065b002928ad5d56079f9fd5b437d1847541d3ad0b5b1ab0a9f7b28314f4f4cad3601f058d7c34f9f6514af8d39964b48d214ec65570ccc99b46907203ab56a7eb24bac9155c9ded3e57366f9968dd3365c7004ec6c924;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d0544025af372ac5c8639f6b429afb4d3cf87f48a170683ebe95e1ad674588e3387ed0a6890c991aa988b8f9e85bfd31442f4e38b19d7dfac0d9a8107967453a5c36367a321669255e6eee04962fefe7cf87e928b13d6b681e05ab727ae415bb066a30cfe1da687aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a97b5e6dfa2be02f79a9da031571cc35df5ad2ab0b667fa542929f4137b75b00de67b7d0b53834cd8c0718861a9abcb94ee37c29054df1d1abd2bc9d66fb738261a5a4277eb7805ab65a287579155bdfd782f67fba82eb60126499e10902cba218e0a8a958ff139168;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1830a1d97e3df67534ffe43ff211bebc1e7a2bfd687ada33fd6cd16c973240df447d47b8bb766e1b1daefa0a8b4d27b050e9174a658d237ab1051e21c66e4e8b432f6acfdd61f6cb0cf9a46d1cdfe0c8c83d03dd2623dd7e142299b96c01dc7ddb6f7c9ab064b9d58fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e91e320fa58182ff12ae262f7fb063b4710f5e386c3585afc2c0ea254560080f84e96329f65b69217037b1191906c73e529a4ef0f21f9f0c23e93b17d63769d7380fd0424a60ed07cfe43c5495be6fa049fd01dd91639e1e090f5540f01d0e212403bc9805b855e2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h440f00a6eba4e6283e09d5706da6adc370d398453d6dbddef9dd6020c78881103963d11571ee00a08727cbb01312c3968fa2eccd15ee9bc5bd72efdd6551681aff75c5a85c9cafdb0d3aaf871df3925f759a5a141feb3ef899cb59e1e42fcb746f22fd6a60509c820c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1933d3a5c808ec59079615c95d7e89bf9420b629faf35a70d108f5f365c8d9a134f3c073b83b7ed2380d167c21bcb4486d310573f62d7af03118c8cc04a1484e9f5d0ece7df575f50e50fbe8930807909a615d0630a5504c50ad7842c92e1ae9116d7f4beb5e48d83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hded822e36ec6a5ff47f02e8e3f8862c80334897e84b27904c517723b1febf9ada14aad87666e4e606cd7dae97ea930d0fabbf6d49c2c292f0ce292d160eecf890c00948999e669a1e9f896a2a8cbe396e43a2e192e2b5657dfa47e257bda7a630bcb53cdbb43fab02b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf13ca01c634895030b1894f3b929cdc0b616f0c77ce03dc543a96231ecfe0abca6afc8d9a90d2a10ea497a4935a9c57607264eb00a8ad36a8aa87542fec3652ad0d27fdcba3ad3c513eb39e7a3614f73db2095b749e4a4518f79bde293e5ec00fae74e009b066cea95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16af9da80776238920170e0de9e5ab571931b73e02a2ff0986fbc12faf928ebb9b48d0e517c9b631c7852f979028ceda41a8f48cf0b2284395c51cdca81acc1354ccaa3c1232814cda242b2a475031360ff1ee1a0765153fb0c2c217d1d450ac9196b0599b46a522c70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eee37b716dd85f694f88e01002e2396f3321352dae9d7bba2b85a2dc61910894d4948d2b2d20ea098640cb624a83a597c2ee0b0015c0f596ae1aba3d16e4f7c64180af57dc59330345ea44cec2329d26800729164a0e91aadab022329d105d10e663d52b76ab929fc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63982f9237e87272b3beea1352b006bab8bb711c3ff249395f5128c820eb425720e001d775bec97b773425f747c9999870c9d48c92da6052442df741e778a374e9df329c2dced8c9622447af267ae1f75749dbdd0538df2f8a45d20ae3e9501807d20da72cb204143c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae9757654220dcb3f9d69d3d7eff287ff70af1e80899d9c8eb5717308a8d21a12ac52b107c58060e4e91f845e96e30be63a554c462b4c6cda2f19b4b1f9e1c9465113c1fb294efacd884df7e7bede4e45f66dea09da8789926120f41c9ba48683a3a4d36ac2b6f57df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f9748867d0c40f40eef20358f85ba488a5ee8b07e80346d2510e4d5f1754f572ef820fc406029c7f2f3c2363a26342fb731c897e9e3940d4f72e89901b15e5d5a89826e4137c593609116b0287444307e231a70a7db22ba1cb22bc633ef71dee63e79ea15f426c658;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9dba5cd822b0f4006ed673d5b65163a3386fdfeff5e62df6fd14b2efc084161b1579dc7b10c39acd6503c9dfbccc07760950eb0fb58f7cd20cc110f77349a45e129041a17de9d4fa1be113bb3acbb5046c98dbf54d3de79f548eef3d338e2c9c66b0a01dc79f037d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11cbb9469a18c104aae1a6d0752442c9dba48e1814398c1ecee671659c4555b93201cfd460e52302fe55c78a8a3d96ca693660705565380bf2de8bbf035b30ca73072be484e7155444e483e97caa26a87a623ebb8894b4384325307e761c829a854d29e2037defbb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f89695a5bb2d161c457bff6ba13c3557690f7db318017d93777b370e95c57f2806e2954e6a441bbce173fc88a931ae7919172f0d129dd5a89c4e543860408e186688ac29f14aeca695c8b3c83b4e6418c0def83f4b2716ddac1ea6ba334d7e0b9ac9055f50b75fca33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f42a6ebd341a124536f132e018d70d144aa9bb6602a474ec63be033326b4dae71f6703b3690c8f783e8fadd7dcc7d41b4818866511d95f31b19a60cea45218b0d818380aa48db3d5b44fa5b3daef39fe7ec79665421f5a877b3ccfc75417417e1da758dca480ab28c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c551d83e3c1ede7392ed49a7027a8207b33585115ff9768b0c5910231b50c730fabea1b7dd02688ab60a35bd37909769551801f5e397fdc909e2ff7ab2013b9feb1efc8c675d27c85dbc398322b5ccdfa521d3987df9ecac49f148b3ec238bd4a26d01a8232edcfcb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a59cd0794eed82fb678f4223b2c4976e9b8a20154aae1e9166d9e915dc7c3648ffa0dfbf6a85c8fdf08915bfc63b318a987e0ae7728c69a5227b53fbad6695ac93adf22abae4a535bea6c56f7da8bee687439b202ea7289027c89c2094b8c15c1c21f4dcbcaafe2e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3b3c792bc128eb05cf4b285228e6d6779094a3e0b646c0d725c0042eec5fbf339c232fbb436ef9870d94de2d24f559b055c099fc66a75d9978c500ced85155f3d8d7826ff0a8a9bae9e875c54052dfb84ed9defaa08bb639064a7a4f493f75408648e2fc4d6830e08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c2b444ff111e653e1ce26aef9774ed98a63ac41963627f824e61a9c5489b473e6d49d4dafb46889212e28760647a96d01fc522a83c0d6b941c18165d9d7ea25f1be2cfb6748574023e5c4b134ad05f287c652df8ff1728259e7fe683625e3c231fff1372086da7c84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197519053cc37fa62b408dbce30a6fdfde8bc43cd8f332022a06a3c090b12b60a5a24dc9f5f692f9cfd7f2054b407a8b5357b87425aeb0e066b7bbe2289c6e4e8ffd8780f0eb5babe0368804dd873af530f946d3f893cdf3ac4fe59c6980f08b72969a8f3fc263b0b84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4b8d59a76f011a1c81e87ca55cba5c219b5606bd0a4e8515952baa3fe9503d9bf7c46a6dd83c50dafba723f110f153ff31212d21ce0d2ba2d22cc0adabbafadfd1219b767fe10101aca32cf9ba2768ba6829048b82de1522139579406cd57318724f8f0a30e70ca54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf99847261a2a09e08f81fe594a02b12a3098e9316d075ac65d9c8fc8ea4bf4e34e081573b2e0edf4a15de6755b2b1c061f3fa2ed7f125f02be3817d890ad84704133cd7d1ee171719f785450d4bfc29342eb9b168b02a45e5f046e7698ff8afcef3366ba1145045f94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1230a60e717d3c87902898d5a88badfbb442acc7e6145866794f0ff4e8b05e98cb3b69d6dfde5e0376101643e53c2a75810e23b8488511795ebe413868ecfb65c23b4572b7df1caa20e4ed85f293947b41702078143759da96b7bbcf71519e8ff6243226f7f6c80e092;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb4f86da92bf44c1878094192b7cd8865ac6f7988b68419cbd05736c9ded7503fa10bde86ebd1902861914523ce67d3bcd5cc9a407ba3cdc67525e3c370771de238a56abf03a8e3f87448568c87f34969da2115c92e4fc0d96bfda7f3ef87b63b9b9d43193ac5a5507;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1865c3edc268ca197d35a8641764b9577e6d0c29c3015671cb1c61de400bd1c1f5b04f5e24934aa52bb22ffcc0b58a27811787e3b8e0d4b9d5f2a84c24b77c498a5e3d0a5b7dd59134ec18277110357b5612c05bcf1bd8eec16127f81e59b0192f23fff0c95daf782c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1794a50cf9b7efcaacae9b3a1accce9ae901e9e013da0a48d10af8c2437324b0b4db67724c3e57b9ff527c03b7097166940623e74fcb8795d8f59c93d3400c59c4b9f053400c1681d7da57f29157655a97b1330af30a1df63d8a88abf146c6c13ee46b7fc75a8ec849a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c5495d4e9cb97c038dcb025cdfc2f7a4cb518a30beade734b6b636769315e485302feccc5d93e9fc4aa50ca825af9bc529a0e1c69986d9b32cac8022548e8d3c0ec37a6569213b415788df009794d2ec5f12e207e2e9f730de214d6743513ae436dfba513d097a4a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f720aee97c3eece82f38fdd1a21a433172408b23261414645827bf658c495fa1bbffd676fcc437f92a28f879a469e55beafe79d4ebb47085b32e93becd298621dcb5b83b909c804a471858b4280262bd50e5c72f35099689e1e12a194ad1059759b3e324a7f1071267;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdef0528f6c3c7b102306b36f314193a646f9258a50bbf8aa01902446c9b37f193d445e4dd6ee45b5809e5ec41feb1669749570fda1a1c2f51f9dadcb64ee513df9fea991abe3465bf63192b406fb19de5d9b795c68763ad4af2da56a9a834372bd66660169cb073bde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97b4d2fa4b3e7772df73e96c2fb668d764cf3ca01da9c40f462247dd1913dac793765a35b7206ae53493cdf5594b57e2afe51208c5ba85477213e02be94223671ff8ab0f4210bf4416cd874e3ef3ded53b17690eb1234047802ad815fea6278417873f96837898c2f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a49802b832807e37c9cc7eae85c527ec23e5445d527ccd030b25390dab9ffb3a72a573dcd3ca2e87fdb50aadaab3f6587ef71fe61df01651d04f8c4aaf432e9a890adc3f53217f9f238c35a91b11fc263c20b42a1e0629374c4cbb869c2d560431245073f2b1cdb9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c639f09fcef3cc3128f86ca5c3a9c1184f571804420eb3ab3732d4153696de668d938911bb5821b0781f848c4c076e8c82584762ace2b80ca314d79287d79f80f39afc35897809f2d33e892dac1da1926b3a4407a5af541ddadfa25f7199a863a2232627849424a41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1219f5560a26cf0bd8fda27a813a4f45063ad9a8e61747ef2aa111bb45425622b087b3831e4c1ec554945fd7468ef881fdfd7bd5ccc29d5fd48564643c4b66f22677d86dbb0fb6aac21b52ab584d892b756d72f4b4d81339b1d8a564c4bc2518796c6f4b63ff10dfbca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfeb67cac19ef264938bc8f4819f296358e23f9eb33105da3db97add17f97feaea52c2efd42811b4678a5216cd28a1541d3aafc38648507d06a86acb302d3f67cd607499125763bce10c4ff3a8a737471f923b5b489993a9a3d24d5cca7ae790f256cb561c1bc92cee8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ba96f63d972826179171f0530861370c82e1d51697d63d5d1064d1e2c5de6d9bc704c17ad818bae22c5e7752aff8545c91c135ec5373655190ada78dc112630cd860c32c8b3d5a725c8a715870e5f2f2bda07e80417783c07d6a40a06e7d330e4f95ee523669c12c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed652fb24f0827384005682738cf9f612e6d6694fc4e3b2e955bc07f65a6942cab007b4da88d08f8bcecc42d71ca907f81b4582aba5cdf6333a6193f733513c016a62a1981068c3c849cef45983dacc9dd6f81f0cb3f28af6301f4f350c7b499dcdc6a3637a39349b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8a35ce77a2d433e1376939fba1debf6c21f009d7f1dbc9f3fb0a9bb08b33b85139df32aeab314aa7fcceee94a841c00f0ec6fc6dc035b62834e77254c7a417bb197a36111724403151e39371c53f081ca67784a790ba0f956d2f7ec6a96e39ded70d068d57e942fb0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e027764a6af6727d6242b963530279db275e8e09586be6b071d620f28276ff9df1138919d6fe35693e4b810adda2409d9a34bd5dbe8398ea095fdfe28ea31f928dc7dc29f28bab59915261b555cbf26bfacb10d08ccccaa276977a4683daa92ebbff13b3f3d82183a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h139ab811b834d64d1ec2ac20c6d5d6ef372766d623c442eebdb2fcf8777bbbfc48ff3ed1d85b6dc44c84b663a74e842884458d51a366c15da489b191cb589a81bf9a7613bfde590a06fcae215adfe961b594be559fc2ea962824bffdc3be75a5917732b0fb6e18501eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82cdfd58672752563f638136523e85f97c9b29e0d6a3a5cde97d5cee3aa56dcfb9ab95a69b0df7e4c7098d1e4fdb3f6afd364dcc41a666ee907971af5162158a96eddf902d1cf5c807008f4443aa33b772ac7276a0dcbaf5e88d74e4f612b3b3fdce53d5c3bf7e17b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ae5f9ded55989f2bf501bb880a089ae70b2066f22a41cb9fae27a9434ac1f847716b49e56d690efcf99acdb7195878bdbcbd2ed780b918e1e5aad944f1fcb634882b1e8f82bb68c9900ea4fa6f643481eb008266c7bc541f43ff474e4553990516f4c679abd57e5ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4959d0825f176a11c7a460250b32e54b368ad9ab5ed5d1bb2f2fb2d363fef1e8ca1ec2d48533a0a874eca9372e13fccf9302acb6676846ce8dd616ba56ac8fb2a58c5bbc957cab72e0e5e9687040da948cbb71c36dca2072c3e6240be016147964d3b9fd33b99ca86b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a7bad8ed07b6d0c9c6d9a89f832013464f4aedff5cb9de84705e99cb279187158a7de5a11fb526c8913ebe1f7dd195f779cc7b4dcd942fc84eeb1716d06d39ac5d957ed85cb80330421434be1546abc3abf5d1c7c33d100d56587ec290a84ed1b92fc0b36d8c08ed8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb2ab57dba4e206740faba959dd1cf6021fa5c4da637304da4b7545cbe4acb0ead4055310eb36ab043faedb6424ba723f7f2c048aa57f9f322f102a5271142f68fc95f1142587d2c7ec527c546bf4248f98cc8ba9c646ffc79d6486e496cf4f510ec9f3d8f0da1c420;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36deb63d5ae798b2a5d90e7d779581eb06343f4f5ee80c2851a7460a57d2445c69142bb3086e885a1a3d18fa40761efb581e340ccedafcc74307f8f8d76c1ea19b1faf479d6e2382227d7fb0de4420487064d775403e8fac694f7c109791e72092ee61f86e471bca7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e68112729963d9961cd6f5e0cfac4fa00123dbea4b7d82d5901293c746eba31f4b56b6c39b2227576eec6999252a446f2d719b1b738fcaa549bc77de3094f66dbd1a911dbe9272f8468070af06df91b6d6c7e4595794f7fb20b3e685b3d3a483b35b1a6051ad6a8c69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83d2c821bb23f1610b61304211b083108de253648a80e6aa22fabf105b1f37e10bb4961ca7cf7f18abfce1937929d61596e35258740f7f69e20446ee7ebefbd351f5a0fa6d064b53b9f418f7875515dcd7da7c42e174103a771296794fae01be3076692740817d9341;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd573f0a3e38c960d3c2052ecb9b6875a6c923d03870684cf8fd612257681daa0b701173a52f9596af983b555aafcc13c20c150607c7f1f8f686c5172f96681eb2a7aa38881e1d8f07eea2bdfc858208be6354e79cb054a098d877f4942b1c7c6aaba05244e07e92ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he567c4f61799b7eb53c7c9d9bc3cc16c1a079d82b23e5c6f855538313d6fe4ff89ecb7926d5a8bc0de1b728968cb210758e7d541e2777f7c17adf301b8516b2aa1f21237103001a348ddc894d78aa5a2a2d9d24e5191f47b8588b7bf8b25573e6482f4e929587176d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142dca6f0ca9f4ca4dbc76d9057be82d3d907c151487a0029d160aadad9e7d4bdd32c380b74346ffb54d767a04966349659c9a2c810f69416a93e54326653ccb7961868a1f2850da87605c16bd1a911232873d8d7c07b483c3ef17b158e4e291628ce6f0484665d931a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da89a78aba0d891efb32102511dbf6c270d09c1d9a9adda82a25d29dbdb55f54792335bd0459a018e8e4ee155a59edb7f88ad3a80462fc914ad58a726dd335bfe98aa9702c73e517f3a214854e7d781e840aa986e01b4fc5a0aa13cd351000a6e04e45f935e0ecc25f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h668086d48b09115d3bd7e99532ba4052435e1eaf46e65b04b2f399384dd951cd0c5bd6ad820a92ed9b8bdaa59fa6181fae24b287bdd463f15e32fe4ab4ea886f36fe5c4d1af3ef5c4d6388ac181bae391e45af4be0d6dbe3ed7cf5ee055d13388c970422457f67fffe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd8372a334934acffe5b5039d0ea27be970eef39656054c2863827887fd09d2d2e3cd874b7208280b912361c692be4cbb4e895f54ee141787c23772344cbf8cfe88f1f8cfe0c37d9853b31c2062e80b2a7ec2e9949d794c55fdf7bdfc15742f7a3998a9d3f5dd56bd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda78f7dc6e7ff5b0434d841bb823f87704121b91e1382c5b6e7e82749c6ae2ece887924eabcecfb04b7c019b7795214213eb8720eb12fd53f6f8817a8c6f3137ac1d728f2a3c09baa4acddfc83ba1e6670c5485fa7851603a13152ca76296546e2a476afc2247d65d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa5b2e9e216cff27445e446d4887bb517484157cfc2acbb845337ff579dbc041faa0682cbfec1b4d924aee319234fae5cd8111add4ce228d1ae1d77816e7216e49bae7a231cd65184d5c242c4fa3ae7e0c90b256e963770d27c1fe9bfd39c91aec458bcdae2fb0b3cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fdedf752ec49b36d1baa1c2419295aa4ccfc77a57b7f10618c92266d7d7010062cecdb97f7a3e8d82c9b3e8650eb17b677b23679998ddde00d11062b263626f42fe81da565d06ba1b52eb2f4032e6166f7261d0d34679379038a5de393f439139bd6b9027257745d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa7500dd59d2c973ec1106bdf7c955dac735b9bec2225a82de570dea24412c4d922cf54a9e62f246dbe88e561b73caa5d4a881179d13602aabf4c42b3fb03f9b2276121948203a4a465f734d39e76178468993615db440479768b1370ba2eac751bc6fb40e4a07f641;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194b1bd3fad5b5a352f926079cab6e27cc6d080f2155a0c673b4d02b156b2dd8dce274d13c5ba4c5b59dd4288ee47f79cd9d486dcd31c99e724c3f4c4b10070b379821d66134884a20637985d08e3e4ccf973b60c60359f251a3981afc9bd7e6d020605a3bc360a8e19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4050536f0e03a61b209f33f51c094b24a02451e8b43ebe8a58e9453a931af2066c9345865ad00dc86bebd453daae6507d75cf66277da7ad6da4e03570e4c7a0eda8cb6fa506a6fba96d1a908adc526bae46eca75234692b88c6552882bfa73c081069031b7c1370b2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he676b609992a2e91a6596f12fb7f8a60bf92a57748a6e1307946dc7ee427ac25bcf869f830a360dcccbda8fe2343ca6facb9cbf168debe1f5cb31b8e4c572a5edf39342d02809ddc4fe2605a8abcc78359b42e4ad6f4bbfcb23d25b76209c14e429862e3243d860d5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197e315cb0f32bf90e5e745fa9ad290325b024b8db18a35ff47099f6af6994437d89de98a4eb8f48815130aac44af33a2ee69f54b594d59ddd73712b935cef5644ee32b2c79f4a55bb156b623e98bbceb0089f35f976c4602e3d4d174fd533e8c7e1cf78634224af15b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a4415dad3cd9fc83bea0d599b2c0a62a9cb6c53e30e3a42db95567017f9b9988681a9dc52687ff072e0a7c29066e6a3eb8b6c1b0c048fa074fc34d25e2c06a521097a0f9ce97c488d8afb5b1384164f22c53125b34f6d6e4b9ae70ddd42fa39898b1d1b804b5c4a41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ecaafcbe2327f2b9da2c75eef82ceffc656e48a596f5eb53ca8d1af40dbb006fc2bb864e8c517512e555edab49ab1f9b26888d1352b42b91df340b5c0d843535d7f3a05e7c91c958a4c52b26450965c24643363e6788a30930dac1dbf679c250852f4f7415e06b3f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af6e7bd29c2b4f799b109a5dbdbaa282fa34ab255d0b56ba9ed01045a15540ff59c94e910f30f9f6b3d6ae167b12cf8333fe784c99760fdbe4fed0e60c599e191e86f94c91b4e2dd5ccfb46778a775b95b31cdf53b7ff635f50e84863c6f854c1339b5c28db4b3ba0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd3e9b44c18b825b9337cdc14a2f7183740c81d46a60937ba602fba327cbfd18750d768229c32516211b16f6e2350b29b3a78bd3d2bae292c9789589311a222d3953a50f10bd24eca5b074106a121bf9614fbc0292e10c86e4aae31ffd754d4bde130f66c383e1825;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ee6ee44d82c4a646c31d7cdd69db76bfb8af85f033a143357a4c22ec7dfee027c5e886efab073bede1f0cf5da65864d6a5fa5bf53ad4d41625c50dab79f84a41ea8b18dacedc137ae44dd6d5bdb0b9672387c3c2bf8d2c01102f8d866d7f6c079e67fe9e83fcd2438;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188c03b4fe486ec7ea8398ca0ba671c666f6891f1004ce5121a164555fd8c8089752cbcf9fc9e91950c1108324ebc00e381d3d985a218194b9bd91585ff125ba51885c1bdc9ba1018237c49702dc488f06ca6e257192ee9f0e41d605a46af0397c08f31f566bf2c6e80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19613da61a6dbde9bcdb61f222957df8d70e8c6cab49d862f04325c3d1182f89f684a4d5d76fe7218bb6822e2faa4890f4a41423a1aea468d79e3e2f51c247f28a90b614f4ebcceea0b01b4f6a162722552be0cf83f0e7d9135b4f5083a04c4b558e7447b75ee07f03b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1022bf7c09122e6545beb8fa69048bb7524e2a640fd81bf31857e5145845e4b4b6d3cd069a4441ce319322198ad2c937b4c141569e9247561f730f6e4c99e43c124382fee83d4ae13406a70c2c9bb9a40e43cfc37102167acf5d6d01bb6eabad8ecb5d96e4163481b15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dddff7bd54c937e51387ead8d723b78855d77ec4462b24d3255e31efbffb989df203d41c27b3d5909c81745f737bc205063ad2f3f80840b5a6a861e6c7a5b019e6d5a22e769e561e779c3c9d2e4e36678b38c31fecb845c20826533b9b4027b605f5447268a430bc0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b6b33f8abbc76b1433e7696fb046a20cb1bc6964a3e7f4a8f30480018f1181277dc6482e22367cb24af1fb0701950c05d4827ab7bad7c029ef6e89107c0d53e74059abadaf0392b97ceacbeee56bcd8f8cf77072de01bdbe248b8dc0334f4ee8aa5fb55c6a6ffb413;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131f1a6e07d3924d2a415d25e1944911bf9598ea3441e0be7d2c7f91b2f851b5f44c673fa7de6186864319e8012c4fb258cbe33ca476eb02bdbcf802514c6acd4f66698d5981627bd824378322519e09d1a0ffdb1d5e441e41fdd884b5b4ecd54fa2c1fb57867d85c59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1183b43b9ddf16708ace006f4f1c9b261ed12914053db74e686cd156de7397976cff424750474e893de6101be314543d357cdc9c12345d571a14f7e5efc2ced47b7a8e95ff254fea2520d874b8d0556dbcdc55eff9e8f6bb7a8ac86db89ed3fbdbe756aba9004338ab6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b3da6f3382ca1da8b34a015044c2106c17a4762acf8df04f739016cc748aafdfd3965ba0eceef496fc545d857fc00a878eddd4ef24b0c7628f8de3e93b767f16e7c3dfb6abc0f9b46eff0951d8938bf37d6379d1900df9f8fe4197af1e52b9d5ed2b00e631699606c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5415e407bd6ac793f108b751debce8d41fa9ce8ed264d66c6c1bf9b8c7dc2120a723d4048f0e2fa0aead32a67f37d3953c610d5fa8fca6096217d7f67be4664b90fe9a721b6febb28298083fe15532c67b6b651b4c51423a6b89b9e4f069682c20c21012069d8e52b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e192bfaff94dba20aa4f217c1e51fbf2f8d152caa5e2218a5822d60caff77cefbbd7bfc798c7fb6ef1d3b13d51b874931d1e11041e85541096695ff8e22da890a96ad49523b13a456a398300811e6bfe3e39fe8607425496d04f6fe70fb23542988cfeb7333e0af25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd957392eb27a18ca06dc89843ac28bfd31a07fd9bb3e5ef773e95485f6f4681e9048bd226712e890b4fa81e8820a100086f60f4f35f4d70ac737895f5b0c2a9737b4b89974e6074d42174be69b9159eb13fc2494c026e0f5a042538e5e96293c91359bfaf3b05db514;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd58022b3e19ebc9405fa2e14347457827c43ea3fadca96f614e3fcc3c14547bcd254de2602d33bfb9e604252102a378c23eedfd8c4aed598daed3e060ed79160599752d693f19cdce3fa6b11a63d22b2ae54a0021ada630711854e554857e37f03604a1897fd8e2973;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1f9951e800175e683ddd773911e86c29d06be3634bbf850c8dcf5608a956b1faa21e6e384579b29111a3e656a39f6296f09f4e6e4793df5c6f8a72a5b6a8ece7fe339bfca570eeeada9b5f6ba2faa557e996a1b9d6c9c8d294d4f94ece16699f9d83851dd638d041e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb01811df26f123bf5dcc95aba5122b223527424e52413cb722b0e406aa6ae199b9c350efc81d5b4d72b37a74cc4480241412e7770da15ea61d3c85cfc481bb6bffba7570ad574b0afee93332e7934014bd1a190c3967589be5484b4af5fab985e870306018c44f0c18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c6d7b2242ca96cf09da950919edcabc42181bb7ce8bcb4631e27fdee39271becf77ef21c66089ff5c2b4abbd77c72cb0c969ebda7ed9a0baebac52b8bd58e2fa6b6b9ca74148481bb95e630f4ac3dbf6a371cbb1c7421c8c0cf463f054fd80d5dd4819b156a958d1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1961c33dec03fc267b983e07f9a754566c00bacd1f02046aa80e207371537fafbfc83ebe6819f7f1a4ad94861f3f0decb807327756c66c99692df0f0fc6187e0ebe769f0c95de5d345984a5d79358481ca7a57641c85b15686cb5c16305dfd6140305a05aef0be15f4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a19ba2b8457143649992e0bb018c2bca89420c4a823d15e833590bcea99cf48472c1b9bd5559c7215ec345e105075ec7658eb60a5a9c40c638331b649d414fd89f248e359131eb6bbbd45f3c269b997a49767a8de0fc4505b628e35101c42ff2c8b0ef3263a433cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha622da6e090499f58f1e6e98a8ad277b0935ed964bc82ebdaa11e9b30c9960c929cedf1e5f10a27fe60c0cf06b0be12f958a94d31dff2eae6ae98513da7dfb215f1bc8f57f36c5f91ebbf3c539c0d08be211bb05d83c3adbc0e37b02e4cc41f8cdf9a416a13985e504;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e07d3dbf30e54216b192dd84e25c6e0d68cc2cb009ce06ef2a39e202855367d3afe9bb1a04974538a072297dcd6ca7cbc58cc998d9362d75e2b8182168775a9c0e26b886dae21bdd622f2e818dea90cf6c9a3d2f78afd8c25d61c2e2bce561935b10f5c3335f7a5aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0acacfd05a8b169182ae4310fb74f463fb50772ad9e64a41928d00efdbe4d8ce6f54c27bb9471402f85c54ae51273f0c6dc6d272c62799b75d86aded0ce5ad50951a474fb85349960bbc0dd7621941e9a7e04c48ef0bdcce34ceae6f03dfea4acc342498a419c0c7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bf5b65756492b0caf097f1cadec34933384963e9523db6881fa0bb568a22740fd7178f57a603e711b57602ae3ac5e821b052e87a13c9fe6b7d2d127af93f3b84e417ea8a75386aae62b1ae597b28cd19f097f993b2681852e16275d7f04bae2755bec7fa21b1cc7ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34523a33ed388bf152945fd8906b75217e8565bf999c9da2a2e6a96ab378aebadb9b1376ea3b7be7d27bd6368da980c44210bc9a04c64bc020fee93f0054d681f255bc53a8cea809fe2a7bfa1a4f19b0ae1605d739f1519e60f21f5b4c5471aeb8388ea3632e7b23fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ca05365d39a7da2f4a0e9f8c94f453281acca422b8c5d3df167fdd23dea5372392b0454ff01014abed28c7bfb2e26b978a2a0ebd3a06523540c95ea1d6c6610b301fa12936bd2fc8acea8ad777487e35f9afeb9e1c611245d9b43ef57cf783be32ac6cd97ee015001;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e1386e45a37929ee1119322e7495a55f52572076211a161e4613798389147a9757163828eace615116cb94299c460ab55de4c92ae7151d302d0c5d737b1af81327dcb55e8d3740fa4b5e409c6a6c88e3a849759f2781c051086dc87120c09d2aeb86bce7477761db7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b60d902b288aa5cb6bdfe598c96367b2026ca8c6db78da66ccfd76d8d9046d554ac3a992a9e3aafb04386f839cb81db90ab5b1e8f0960363f816c22054d3e6a062a5e4035531b27d5c2b2881293be9a7f3c7789b502c7b18a557ac5ed11a4cf321a2b78cba93b4034;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7ec45f0f2d8d16d744b1f20b3cd7b831bc9e554eb3408b594cbbf7e7f5426482f63eb8ee1259cc96502c6aeae6104eb917016008eaf59bf14161bdabcc779365f005b043972fc6815c21ba9247ec04fe62c3de14f03dd7a860e17ce20564f23fd1df453218ecfd927;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3040978c9eec5e6a0baad59f262f39e156de88daec01e64a465a5cf8d8db666a6fdd15de7069621499fe135ade6f45d87335f4f2e4a13bf074af199de05589c1ea5c9dd971a262e3db473bc3a57e1b6d8f2378feb07c370ea6bf6751b07402fd0b60d698f383e4179;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa091a1998896cffd6189b41a45cc45aa2cfebb67a73afaa47dad54fed614fae2ec9b2ba34eabfcbac9e5bfafe78aa8066174cf6dff55a9e9d969714a3469c67ca15a495d36cea8307ce7cd7559902c648e62617cbff73ffe69dc5a73216ac89b48fa7acbf9c1017e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb98b8ed2fa07eb1127763ddb613ff383ae904359a7a4cfa398681a5ff7498d28b813756a29c975e611047d87328bc19d41e95e5c1dc54530426f79732bbf6eb3f12c6ed4e475c39130d9398021772942a4a454ffc64b8f95c90cb736c4fde7ee14cd31312c451348a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e6ee3116343d08fd95d402bc26383db898ebedc1b1815e779b2b17fcfd57fbb6b9fde5f68b1745cdcbbccdbe878b774e892ca67a3bb500c3c32d31a1f3064fece3037fc61f12d6924c667efbbe1e9c8b2a1c9213d8bcdeb6411376d62a27256ef75426af677462dd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d9e7e5e63529a86125e77598858e04237a30c1642944b08183451dc9029d1b8ef717a87036ab93eb22fb1fef27f9133576eb64160d86f9247039c19c8ea1cb9736137fdfdc7ebe6d77e2af8661dd70107df38ca6db2e8652764aece705ccca928a11339ec91a3b8e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb9a5412dca3455268c021908040859b7269ee7de6ec484231143fa1ab8d478e3450f2bba7bac6291baffa0ba05c7e7cb16ea150018bba7c1f5dd515f9a81fe40bc2e8b193e9bf57c6005eee13bab516b37c6296dd0bae7885ead4f618e3df4e8f460adf870d283f5b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c3dfc67239e476cbddb8a14b17c9df4f8809a053902ad4ea010a8a7aaa4c6819ce93cfbf3ab5a3e2beaa23b07d5d2b5a7a59fa82c545ff8585272c9bec0244af9d3ed46ffb17223a60b6784b5521a7b684de2537c15c165a43e87ea93c0537da466ba1bc78a0aadd5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c937c552cc16e6b020a927bafa3f4c1248fdd7f33523ac28af3f2a376b861381530151d6129eab9aefa2146b4ffcf1259b17804c8632b2ead4e7c5a8d2d725a4e8f2fb72e49613e764afa122433631114d705ca9db1b90fa67a47c79e27846cc09b2518c1925b577f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15bf3860b38c4621df3cdde68e61693393628a728c2d29bcd70b46ab05ca4a98aaae4a6c342683ca15aeaed2063ca23c83ed3497e47eccbd0c433a60bd0ec3f375b0d4211c849779bcf1529359f2543d616d903c391e624d9dcb7c616bf4c294379c24d473f15379c0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10dff6d983237c7ee0fa4c613be081ff11f09130bdd9e2b9523fb5e36d332cd9b7d9ff20b4ce17be4cf0f8c4e5444586d7d09980c35796a00d8498ae9df9686b629473b3467aa213d089660dca03356cc48725adb680c98c2227ae52235a43e9070582e79a7219a0683;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13caecc2a0ec3c757de8b7e1111a09c27fe37341f9755a4ee4cdc54be57f45f8ad781deb8f0a980d8276fd7028981129201b502bca21ca4b278aa77064c91b61bd0faaaeff28de182156cdbb5cd9d2b0fda441c44363fa799e93ee8dab3a9d855c0407d0cea3d8eb0a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb22d58f05cfe20462ca831fed56132c63d0993793f7da80f8f515934719acf3f81e75b05c1151f15aac2770c4fdfa6cd5bedf6702ca8608522bbfa054e24883edabc1bfe536657e64de3166458fe019cf983494b427a4223de881813de560546dde5bac5fe2c804bc1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6b60e6550ac3f4e51ea1db7473bccb1c11787d120ce476a82d9a02697ce73fcb3dc35df2c3bc19de5e24cfec8e872de1e92b0ea07ff9e9b73975f58f82130005faa730d365b098fd816d84ae9b4ed35f7372201f659dea0a73cb777055f78f7d586c41ae1068fb531;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd318c870e0ed79ac6a622f5d66364f024bf47044d80b4547b66a0c75d4533df3a75105a195aa8a2df5f9f997f49dc1efd9bc995245eda26afb45a54b368e0e0987508130cc740d016ee3c075c0083352b4316e9c2c3bb7628dd2138deccfb57665cd353726fdce7d43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e38fac25092167b4d4bf628e6ff904a64cbe8e30725854e6defc03ce5c2044db4331f3cba82216e3ceb2564b582aff9ee37179eaa1bf9e23c01d34c89283f95198a57e67dfbfc0b54098a12e70c3e777d64740b78954599dc3eeedb357092480a8ae5efc2c423aa1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9fff03cf9ae1ededdf940dd50176cfbf8bdc04840c129e272571ea85c8c54430a36bfaca6b4bfe4e0f0013d0e5667099ce2e029fdea3ddcae0f8553f80755650164e6fc703ca0a3acf74ee726db2dedbfde38e0407248d39762ed7076397e68e9a406c7b019bdfdc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acc5bbf7a779c13f221a0bc5ab2d0859c796898908432504e4aab290f3aa1bf3bf618d1b42cde3decfb4c9c5f788faabf7ee90715bb836f2c645912d87938256a200592d39fe4fbc01993027c82d7d92ef9283931ecb577fed5ee9d593dcbb30889790fb742f497c92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb4820181a8c701d2bfb6f33e7ade6870ca853f965e1f3b43f0e5324db41818e8a3cb1e542d9fbdc0e38e2565aff4b5c24dec642fc878edc0bb6f00016c1fdfd6f4b491c108e210ad01389c3677c5995a591838823fab4da191c0e627c9ca5a28226d12ec9b2baf48d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3d11925526f318283241ba083e8c5a0be756b898255ae702300cde08e1bea827fcef36fb3d967c7a4c512840be7a99b6fca3447d05187c239b641ddbce9bdc43a9291eb5f68ccb643cf4fec251aac9c0476a3d8fb1c6f9c74e082c25ddd8a7ad160a1df31387bdfe9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9fa7a1864357a83b7b17a94242e169866e92c0a9d1e971b3ff6ce7dcf28e109888295be31546b96ec104071cb578f1da2a986539152efaa7eceef3530cb486af29c56fd7efb735d268ae904164bfbcd8701159e84656f4488a9378e496611c23d4b05e369bd7fcb80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1217558bf9a3fe6a6541e36078be79663312220ecc959616e8bda7034c884109d9df26f4a06ca6b836b737fbeaf3b89853944c6de35761fe98ca51a5c3b01538afe2e209ab7288f42d00d74db2d2b86a1b106f4901493813042bc4596c743edd6a86f5b1fbdb473b113;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1adae3b8c607c388e4a1b5889fa79f399beca5bdad7363180b89dc9a527b2d1973671cbe8e5cf6ce735bdf664c81fecc5ce5aed5e5704dc90f79561377e466fa2b4c2e978cbdb085f551ef3115a045f3398dfcedf72f6e0efad6ea4eb70b1f1f94f0b61992acab1a4db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6df6c15d96fe79c08b853982261816145cd9087a43c7e14073fb5f10aef2d787b3c79f3f20bdb20c8639a1b683bcc67094f18465f006ee77c4bb9ef694c1206b9ea5b2f3c5b81a07014d86297534b65ca24b3f8cd382bac2f46cd468b24b714d33a43a2ca39407cf12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170f1eb1a86e5aef31f4cbf283ee0c1cf0a28b976454e8e4e1d54781904d5e043f09d1ed4cf5cf185b6b9898595fc0dc1c3dca8bb1c9be63a61986ab2899731012403f003fd7f686e4666dd74bfd3b4396fa59142f9ffd4516a57e3ea28c26860c8f185797fb71a4311;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b6d83ea0e3a5e84ebf5d37f110d5d835c49b8ddc17b53cf2a8030bdf92059209cfe102c254d31c8ec2ab17b0ea71ef454296c7afd5ba90a4ba37de2a3ddbc95c3e21f2d1a632b3da1cde8172990b6d07bc83efffb8e413406bd6cc6a65a890ecf00f326da556dce00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d0603761e214607d8c85b5b0481e2031c30bcbf8fcc4b1c5a636dd7791c2452caf05fd462edcb7e7a406abbc82fd81736bb04be5d58d2d2ba0ff67a7400ebba531d14c5e187131748cc02768956d68dff9f55f1e27bfbe5601922c6cffc68c0cd0290c25392dc9cf9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h565b02f6592caed939715ea8642539fab4fb5319a6eb19f02d45d24744af6dea550a3c33e6803dbe6e2f1a01fc878a44c438bc25af245466a8014a60fb3b00de1e6a8cc8ed3824219d3cb2ed3618e32718915cc1af094d31d9e1ca511cd4b46384696aa03768f0a3f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac7f15276d6c2b3e89a965f34e8001a9d60438650c6cf51f4dff963dc4eae13488cca41e66c00c45063886742f1390dd3a609c90c85fcc076152a2b5bb935385d90b796533b8d7b352e8985dd945385d1dc59fbafcf1b5daa9ec1d778c471ac3e526691cceb8bccc4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fa411fa2ac319e46a1241c7ef4337fc472b2a04bc894db34cc4e295f8f538799cea40a27e0d7ac41041c50c8a9935bf590f3db58df14e2f7428c04ba8eae12e8fcb02c509758cbc896d14458dbfe1954686e0e3dd4d119e0a1e08dcffc82af18a632ad9633c467010;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10714bfd225f4eac96866266d6d3cc87510123ca1af1f061505dc035f2635fa751dd32ba248cb976c50e0074aafc39003390808360a2f1f88f44908445486a39322bd0f5a2bb7fc8cab9c4a74105e235f4116f0b42bc15dad3382399550a0781c195b5b9234407ae21d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cf3377f06dbc3f461a5e2829c4d39f238d9c03daca7e16a35cc6310e54b9f72a7c09c0ce207d149e80c33b8762a267552c4b7f8384de016f0b9e04acc684cc8499af6cab22e736cbbeb1c50d3e2616c4208b6b57ef74d17511cccb4a36713d927e70f689b5c637fd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h236d23f80fe824294d56a5b0171781bd3cb4abf98f1c8e1d038e12bd8f0e79068f49cc4631364af1986759f9c80877fb2006c4c333ecd6bb4e8f0e3e45cf51e5c5419bd1846a1efc15e856654bf18de06fbd5e8e42497fde220758e2fe0231451225d8258c6f731255;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ef2570949d6ee0be92ff194b37e97642f8c6bffc4ee3ace401c6d9ebebb18f1c25f743fdfceeaa8a9f006efa991056217f685f8d08b03bd48a51c2ebe8f73f2b7d345a343140fb3e60c3a6f85d66e35644ee7f8cca19a02cecc89fd03bb1a0594fccd8895318ab4e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a255dd42e1ac7d28ff0c818f2c40bf7d22abb5b531bc6c55b31e02a55a881a2998899ac0802d142f77a18bc4c09a9e068c7a39a085567c9c34f5ef762725a6e93757d76dd8e7bcd57bf903eac43b96e22e975e24905c0187e9e304a4ee4fe21bc282ed24fb1670cef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4a47ca8341720ae607613ddaa1851d5e345d1009b002ef0e56fcb581cb14ba7774eb47ed5d3810ba96aeb327be62c6f47c9f5c2ebfcb0c4dacfaea51849b039025f6e45816b8488948058718f93dc437c018c775faac233eebc172130d64bcf1d94742251ea541ad5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec64c115c279e826aa7198e362a615cd05a49971514dfe9aed82bda95a347e108000f24ad0a8853beacfa6b2641f27c3922959d0e3628d7d98e3e5f2930909c8396c34da3fccf20da15c12b2d6e3fe974aad9336c1f4c6b95391928bca13b314e2c21902d63819f77e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20a42fa8fa28cf63e5b0fcecdfcaa33d45df6ebcac3ef25ac55eb5e3b6594dc2e5b7804fca1712150dc4e91419b744c8ad77673465166fd714b46aa97c0257492d59b971192c5846c21379c495e8ccad70d95c622b45f78b595204bbabf5ba53654a98755f55e3d6aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fd7220a3952c88ebb248f8935c47d3055e507779047e46787e0a0725faf08f239600f5a85514f71afe7e219a06b3f39b97115851fb5ac3c112c845870bab597355fb763485746395dfe9a88afb2f1f54514315660d9c1bbe0b3c5723bb860cc7db3f44a093014c2c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1996170c677d9f2601f3962f89347325dd413554a890527eb4ac0ac1596a1c3d83a7c20839a00bbeb962a6f6f7d50a9c5926a48f7e5e8e23c11a636effd8c8f06a96057fb3a0356089c21684f5cea4cad38843363b58c4a0fa6e97b8c7f4f605b702e19c3e81a30cad9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15731453257da873590753db7b8aace25d171030ce021aa12eece9492f08586d4ddbbccf2a29c3bf988a0c647f25d0185342d91fc07dd4670d65cb54fbd727e7fda5419be5012cadc9fe803417577818161187336bfbeca9c394d9e4868643207421c7bea5015b6e96a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbc269fa2925ac2f3818753219397d35e36b5953d81301953aac6019d3d38382177c58ea2057ae3e14ac34f9f2b76943bcb50793027359bc41284501f5eebf1483dcfdf522f5ffccd7bd9953d4707f98a15d90566767cc0ed025e507c062bf1a9feff4489752f07fe9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3b613d9f625104b93259c489decf5efe8d1a02247e11a94b2f8278bcca9a85be6eb9c973c9b92abcc8fbb21e98e0f102c7637158ec86705479f43f1baf55178130abbc90a4d47088a8321d4abc905c16ac4709400193b23567c86af6d8a3727646909a26156b55df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f306af48cb2ec27b846968e8321ede84bf7f4ec98e689f884a4467d27d2d45c2dd76b7e492c13227b74febdfab195a24618f14aee390708da00686825fb648fcc42c07a59beab969a7a4b297199659feaaf9ba5c5975fcc7f1308afbb77c94cd7e462dad1bd1fa1978;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9253fcb6dcaeae26cf42e87dbeba457116084fe997ac00e3fa3170416e09fe4a281b51b608f14d40d315307fe87fa710519afdd12f48fc36fc8f67a502bc4b87025e0f37c55fef06198f49d08700193d1158ac5a74b44be29d7599d120566b80223c0524463bc65976;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha56528ac11451db5e1b7c4044efe5f1c8fb1c0321c7290f14bd2e3d5582050a0da7a4525eee4bd43bec0cdcc3227040f1d9ac837609862c8d13f806030588cdb62cc5e353dd0a38e0f5ad9a276932c6ec666a57c7e109835e7d621c4d4d52bf688f1d32bd156b6ab11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ab87cedf1b78f5b1a611f8f2213dd3dcbd49415e4807ae2a2fb75b0e4603c89c3bd8a88833a847977e376c69cc84d730e77585702f95901e678bdacc301542abf7c743fee282e7cdd657b45606c9676eb105b2f5a085198dbe53550af2cf08a3b56b2b4c36f3edbcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18eec66ca7730f2c7bfc2f27e8f3ffb7b3862dc5f075ef05663e931314e2410ca4e0801e404a9308601a843d8500226703a104650db5f72d0838baceb8b044aaf3e73ee1c52ed8a9b952630d3aea9efb96c4f0daf29df5a7cad5e060fdd21afff3fc619a4a961d0ceed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h275632587aaf14274cd445944187a7f782e97d644f43901f42671700c33fcfb365faf9dec1e50445ea13fbfd148780b812d58f6ac706b689a2f96e4b492582d2d21e026c4aac5140bdd8de7994e20d384dc9d7ec54e4e5b0feafa2f203358b0989d7943afdee800a91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51eaed1c854e9d03772d1cbec639c16e44540df6ca3e06a59d29741a23b3c8f69224fa2736e501f4d43759e601e0f6a9ea3c17c9eadb36b649ffa3cf26ce684b9af1be6d6cf1de2b895b1d69182559d929ba55fb46221049f99270e486df5b0a74a318646bd30b6017;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4826612d561293225434a82e708cf345d766deeedf49fafcdafa71e9ac35177cd66b26e670d9374ae4f94e175e9c269a5fd15085951b162ed79b0d30704bdee8436f599040be87df541f48ea2d9c6507140459b1f80c38b13cfd51f57538b333171c75b33cb582b2f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h730f7d4b8bd3018f44a9104064317a35361b1b423ce3b44a9c43e3b53fbb5f6d0a54986fac98157c47945ef0dd448a15d581a12e71de7f95cf9dd328d5b5c0295809425986e67b2d8400cdd93acb36665449df46b7ec819ebd5e34f8177411e32955b9a733d24a7c50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171c410fec1585f88628e545c8aa1452366c795045117506c2f94208a25635dbd3f361685b98c99bab1ec2583eb1c85c27eb35b92edf7f5711559bd933344f6a107afc88f9e5bcb4b2733e1386b5ed86d87f553969bacab71a3ca7da05fd4036e6a89afa4a470c9f978;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1834122923ee36edf4d53f643c3a871f44b9a144090472e44136327f0cb0160ea44f98cb7cf8259f3e4fe5d5ef9ae8b89becf25c34c603bab9864e10e8e899607e2c590ee4b11fee7293052384cc71984fc7ea9caa6754b9fec0e2aaef08f270afce824e519a7edcbd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1346be49c1ef5bcecf9a5e60f63d8c09e14b36fb42b69a9d003b31d6300c0d533c3bc190ab30c62a0915edc3f2851cfb9bc22d9aef866807a5fb558a8e9a248ea2ca1e8343cc5b982efe99be2d5ea0aae1a64355c5783cf99fe1a28a2d3a0802ebe555ad3c7eb6e5032;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f85adb29b0e77e6463482e01dc88ae91ce275aa3576dd982a25fe5190b54deb49b63cf4a735f4dfd155fb9ffdc63e1f5de2169bf15cdbfc2152951f259b50944be6d2ac7ad8ff79eb6f7ef483e1fb8c7e12371236618cd7bd2ea2ebfefb6def0c2a4970a3db6deb97d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cdb4a140c477d3a99817346628445f78068a4a6c70499885e176b90fd26699031ab83283f6c1101c890394753808d5d64b27a9a5d62fb8ae82ba928b1e89bbaffbac84eae28729a2f298cd70f1f04875b29c6cd99d58ba2c0a8dcf9343d66e0e74282d177dfbafd14c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf600001923f4a65f89c9113c35853a1de0ab385498194ff365aa121720e6a7794b7072b0c4bfb5cfc62ac71f48587e6dd285c0b71dee968f16e04ad4f15c5b6390a5916a4b770478fffb45522109b3af5c5cb500739df9e8596e7150d2f7d02756b43958572a302fc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdddba28d682b85d1d4dec9081f80de8c8e67f581c462f855d84300e92c22522ef57e64e4641855d0907f7804ddda256de42fc5e5edeff1ef5271359fdbc2822e5687dd0fd37ec0161bd708b45366e721a320278a507d7db9da12c8b7b373d4e52007f946d0eadd38bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha221256cff05f9c7fbe11d6258c82fc55a712b27f04f7a46813c95bf9c8ed36038b62905b923aa92bfc7dde4f5327df4b268150a289802bcd11bc40acb136881adacb1b7b570de06ec7680cad106c56ef333aa6a1acfd88b612dd2f9b870b1dd01e972d9b6caa17309;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1445513460e61cab331ec8b14f4b110acd34ad6f3ade7cd49ce90c3c7e68ee9e31f6d169ff059e799046a17fd214218331c821e72015e93668cda87984797355deff5643d0b25fb7fe19ba13c23e6469f3b5ec6b205f31e99341825f55240db2447ab4f0116ffd84f9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a93b99774ab5d5981167430dd13ad44ef89b224212ae11ec62c0b8a2e9eeb56f22adf6aecf959625689e1ac1f9bd24dafc63b0c5d485aa6734442d06caf845125f90565d1b04bd77e8542f95c1c91fdfb3ee1a5b50429e2dbfa2c95dab4dff73e4eba103dc7ee464d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17610673d5eeac42904f239d92783d953d08861bf75737cdd8df37e5d0927d59c316525b494dd30099e02174f0b92ecf18d31be6a0a263862e6aa7cc45dad83081b746e3b5e2f67bc8617f060ed17a0b1f1dbebf9686387cecf813ae7b5c597cead7ab7cdcddaf30c40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70e535270d80d3b0d484b1037f72dc143a271965e170a2ce053a5aa06848bef0e3db44ae447444412a894a593eeb1a4c072b367481400ed23e42b167a538400a8e4c6f28b56ee258fd11ff47c7af4fe6c7ca1298949b219e5a9b37333bbdbcc0ef970ad361b147dc78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ec129f28646cc04ba5f4ccc0285c5fd953e9c62ec3de9feb5c2d0036665274b59ce556db72def1cdf403c7e590dc3f9d704f3cdc354972048538aa67114e9f5a7b2ffc6f69a7cc1dfd77433c4d4265d5b8630f6bacf2befe0e75e81f7edcc019c04cd173a8e1456e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0e160630565901523d76153344fd6fdcc1332959b5e34a42202ffb023ee07c4360d6220fe3fdd4bfaca5e6a9dcd6087acb3a4b1bf7c1e27ddf96c0ae7e0077f2d1ac394f9118c8beba6749ac0a255fb61eaaceb4210f20ed98d154a9da60c9483e8c7ad3cf3039cb0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca364703bad3767e26a60054eb3f79bde258106df55bb2454de368a9563eef24af1ebed7d365a573420d8fbc62f1f4600958d71b3b72a282b7f40f09a9daebf5ef3383a70166897d246d8947b03ff07e3ff319a98c18e12bea05c50c00babb0c53bcfcc73fef7c3260;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8052eab8269c74488938fb5d852551cf8fb7166b31a0d2829201c8eaba94356384840e6358907ec38d88daa151c26a88fc4420b2d7a94f8042878acff17ede3ce6ca261dff5d0415d5bb7ff0e7a457a609990de499673e6ceca68b4bbcaf501f34b7934a46a67ec53b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18464440ee382f51bcac9867c38828a1314a4e12929fd79e5604b4e7a1602d6a16935a9a8fc54cf5d865b1dd707d30f9f0746e934243cd6908ad74c108c3c57a5d49c35a147b753e5879e3ae4e3116e2cd03f05baa99743c228ecad0846bee673c5cea29a81912524f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4197be84e92a331ee572f987bd1090dc6b0c13a03025c817bbfe1725eeefe75da509f5c8a6d946cd8e2c5f58a3212b37e8c4e47d8ae02b840825e43f049f644eafd9e96145cde8dc8ea5c78bf4a65f6efa90fc071a52913cd7001f823cc1f1897adfbb01bd914876d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a35a14a03e38e957aed0ee3b054d7852ccad5c67b4aa71fb34fddd9a3f6611e08cb550f02966c41fd11b5b48c9f761b93263408ca4832ce16f2f7697c1e5146c80b40d08215fbcdfad069d18f18397ababab4d4f1025cf218347bb6babafe3383c1fb013f7949d7f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167ce66e8e8743772dc20e52d572a9d274a14ace00c3b790a89fa7ae32616ce0f327cf477964c56343262320d0ea363416781d60eb05e89530adf3adafd04e30fccb416a030b10f496aeff679e36b0d2f5329aa09ce5366d240b32d9301a6c7f6520cd4fe1fdeda5e37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170eac1ea64341eab598f1f436ed307d0d14887a54ea955a57d31cb249b7143100705a0e1da698dfa4f405a6b62147e6cb7b55af2a2fc5e0e769d64fbdcd20b7694a341bd1a60e7cb5b0eeaf55be6304aeb7dcc65d3d76e224d65ae8e95917464133386ceb94ba64677;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4e3027065632b069b904c7e42464585509aae40960c9495abaad31f5e642563789a204cb21585a2c4d4047d4ec2b63b7fc3d92d0b442e848fb7755c55e3c7877985f1d2d14b9432a03ee4822df059a1d7a87d98cce4d7630b5247e5fc252c0c60b0a1b7cce80d1267;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2b95459a85d553348a738555372f68cb29df63f950220791f856b6a0901cb25afba14a3ba1c0e58c2a89f78cf1082e2298caef91864af77c7d1132f431b51a58850f4f04673988f9a98019cbf2d5363eddf34f750b9aa6dccb4650de669493aa00a60d039ac97f568;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3124079c249086dc06285b20b4f6b49b639dca1401b84abdbfb76d6303b9ef2c1611788c66f147a5b4b9e07110e14f33f8bbe0f91b41cb6d54ac88c1b1c91d31df1ebe0ff0f4ea92f04fa567db8c663a3cd2e51873a7f0cab25ace08f71b305d51e280db0abe358f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ad5187362c09e6a51ed7fe0cdea6cbb6565a52f086d05712f0da820522d5f23e4a45b5c447aa97955d1abaccc917076fac1712abf752cde3fedb4688fc61cedaa3884950be53d8633927df0a08c1e32988c930a3b54caca91b09a08325ef7dc2e79c15169428465d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e24d982e24b1b7988abc18f9de4d9415b3e4f850c59e4a71752013eb3c42d1ca28b1058cf4b45b1712d1f1054a5f466239d5f1647218b949045b3b90d792520a6588c19a45a7dc0d3abf8cdd7de9ca987483cbee53e56a4f7fcd931c0340bdaed68da8215310c22b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161401b843dd91e8ab833f97e55c7df0289d06302061183ca205a3fb227835a03425145a22a3dc52986cebb76f0e0d3aa2bd42fd8d7a548bed4f0a1dd842693380aaedb9664449e8a9f32cb4d14b10f6dfbd5afa3ec8c0fb426627a757e2f5951da5e7ed52c04f53357;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101008e5cbe5d8ce80aa23b24ddbb46d4b6d70bd3f5e80f659a8c92e6bf23ef99ad4dbbbd908da011a78e63bf05e9fca27dd4a2877247eafb6f4539ed610e67a7d782f63ed0df508280f2e830eb277f7f89f1ef657b0dd51a1faa38aed43174031b31665aca5d9ad8c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d774d2fbd5b50971334eec5192ae1b4b2fc8154ab5222dbfa6abd05e89018e1b87fa5cd2fc6748ead8fde4e814516a065bd870f668799cdf61b4c6b70ae54eb727f217564feab9f4223639e6a8adb6b6a14001e68de8be9b88cf72ba22147ae195800e80b06ba37838;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he23c297eba5e5c0161c39b8a2d08e9b5481f97cf4f0e3ab73983f77eaf44ce36ba323834f5fe7fdaee184f4e1400ec0d81090e9afcf24185f9c65ef7b89b5cac8e34aba9464e79ffc28d60bfac694d75c3c63f020a71f5b38c33195cc22f5c9585541f15db120fb37a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13be8fc1f5ab66ef16bbdeed47b15939487a00f8b393a2da72e14a9a0cbdf89e985a627a4d19e7a64f0afa8b666630dac22885c4de2bb166e46cbbfc631f61b28bc858429c3fdb583365bd7152e4fa0c700925f5ce85d65f4b441347ffc933ee9caa424186bbb4433d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd6b9bec0978d36ab43865e3cfff2234cbd73ae30650822c1034ed7858a3087c71f6634262af3f75e83d4ced0539492a0ea8f528aafc7b8429fe83bfef6b049210c305a885a43beea0c5bf3093dfab3fcbab32d0d056ffc2517dc9d8b9fac88e2a9b88c4a32cc324b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abab11e450333bf9cc3eeadbfb1f97ceb2b471f8a6740d000418209b62a63a386d5561768ec7ebb4da8ed1ab49cfe842689d2e369047542089f316daeef5c9960af0bb5f9e899c50416ab9e025c32894b3d2736b63e01c95f9ba9b509ec203801acb1e83473d18b5a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d78168b2b95c1f652958049cf42dcf356120a0f2b5b9571f6ada97665ddafbe24bcdf5de71d9859e33f3adcbbc47b80f5be38140068073002e1ea83d101f81dcb5175bc21fa392ab2859c86ca004a3d8112b0a215e30465c48c0801b5e9b67dbd640411796497d339f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38f98445f143a9ccf533c1705145dbc22618981f9db193d73abd004fbbab235ad1df5f2967cd62b16dd9e85572738cbdf6fccad72fce4386a1dfa2e612307d510ec2414e942274436d634f36fc21bec0df52daba7e4ac5aec1236c71ee85b866cc0882aa710e72f305;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed5c0271ba49f1d6b69471175afefd19b3e7f1d4cfafc307ef50a18ca7a9fe8d1226da48f82fa9e79e40d798b03fe6840465c6bc3486302f737542f24bfe6cc73de161d3ebbe41c9d86d08921f45a0c385fba01b740776169bfa1fb08756a28acc78741117c04503a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2aeee2fabe2925f11fe0f25774a8221936a76a0d3692755f2318a2e57b423589ffb1edbcd59bad95afe6ddcfe11642a80f8db2370f3bcca4d045fe4ca5d4bfdd7ae11ad3e63c6b7a79fd47d1869ce54a42e5990d60fc3dcefc019ae2490a44f2105cc100c24d7c75e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd99b3275027d43bdc972c822797aaa5cbb72c95b145c00ea4385c44bd881c734a28baa74a1394acda955678528a99fa23eb957cad17c0913c3d9a37d7ba638e1b068e441895cab7c91e71a79b072ee55325ea8768eeee8a6831cebef1236568d9c50fbb328906d1ca9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h582e0358aebbb39e10afc940e5fa7c53a696495b4e12a38ce218a1725f08565a6bbf550d07a6f5c079667878f9c6f77ba98883403e684bba00fe51c46086268a282d956ca75b9d73c1ad690bb0a293684f93747041e881041988dd3a4a1ea447ced4ce6d7af1d62a72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6bc712c49a6ea29fc6bc2dbc64f958e4a93c9f5989d8c8ccc560f03e173e1ef213c371a9924660368cde11cdb41f1a2f3e772e7fd35bb90c707430419b7e7547919ba15a657a9163b39b9063d7ae19186711e21bcb13cd9c7f4ed61e1e622aec6ab17374d444e1126;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h609afc108ab25c63a1bfbd15985b87a4a7906e753758491665ba8ca1080747d5c4ddb5293033c628a5e41c72cef394d37af3621d072fc3beaaff233a95986ffd1beb32fa453beeccb00ec7e9756209b536aa646ea8e6034e369c8cdf8b147525cc0809654ab9c77c7c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca03fecbce5a9dc98e13179e65d7fbd84a4a194b7c72c950a75eb31b6dd8bf879eb4370ba5a6dbb0e143b6764b9ba5e9bae486bfc4b103bcb4ed4076f4746ead185f1188acfcf1269ba6a5f27af128fb4239f63a517019f40638dfe21e91ddd106c86b61c6d11dfae2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb15bdaa32f4b56666082e2b1640221034018644497d843bb535e813bfeff69d2d2d12152077c2ebc1f9cf9d0bd4090d88defd3a15b8a3a4385c0d524562c56ad6bde1c3515817dde3f9e2afef074a38e4fb976b52b5228872eb45249431e017e32f345715f287e4ea8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b167a7b07a3d48e2c42c4b56d54b2b9a18afa54da90abe043f99f079621b6452dbf6e75b1bb75949abe71f869a5423335ebf33bb23b75bb978cd21628df5d615332961a436625b9e3b3647ad925950734bddb5ef3c8510a3fc1088584f1c42b54d6fe8a7a1f5da76d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dab20575438ac1b5d3b4658478af472ba6c98348ff88f5f9a309bcc8a059f63059f2c6d6a96b409cb89ee3a8add8e48fb2f26e83e89ef26341bab48c3ae08f025bfe004613addb5c438043d0848c4a4e1e8858d1e5bc694daf48fc6c8ba76b9368510eca52e404434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16694c6c24be42afccc5e733d4ab658c18e65a43d3cbf7331037a8727756d21f60f3f9fb657108731922c667cf41086f3698c50d4911780fb5b478ed93eb21d8a4a6cf9719eab5cdd030af960943654dc304e5cf4f69f780c6f0d4aeca8cb1f2a5b8e6caa09a72c293b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdd537776da8af374793d31947cf368b36ed1eca71d06e8900f73893ef769ed3948504bd6b7592fe1b40ba7ddd5abdb35606ffc513be8ce4959bbf8ea74af9228f5be1fc6d46abde40568f5f1a8b208ce2aaf6e6e780866a58fed5525d40c124c5ae7b667991df78c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182b06c9275786dfc337e4f192476bfae2a8000ae9e469f89c89e8df5edfaeb8467d99ffa656957c850018241f8b32a72f91670f1985ab47fddd8ce3d01d82958878f8cf24b32a9da31c3f7f0c7c0fec4cd80d3f90a12fbb866a7dcf1d0c033e22d41166fd552b00903;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf02b7fe90b2950b21e61acf9dc644173210457c912478ce1ac17d4f5f6b3581cc60915dc78a6cd480f4b973ae40a4964ad98215b2dc0ad212961e338c3fca9403cd39ed09dd0f0bae938a07137565dca99f42e1cdc0682341997e6a695f5b539bce54f03bf9551992;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1437c4bd494a6f52ac5534f97dc4c60db210189e012fd78b6af27e89f2f17562f223686b349ae6ee79ae21d7ed11fee85a79338819e203b5ce7a71aa364205dfb7e3cc2990a33574c4a0dfc3d21202096714aa8e640a32edfd99fe3cb7cca4bda657271d6ded9f49c02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1fb681ca870ceb88b69ee5124ac0a03adee84f8c81bae078438fe112246781ce42c2478db1ef9a83f989c87eed567014450a645865afa5bc527a6ff54865325e8ccc17c474c15c5ea3eb608f6925f0770cfc857df28ce0da170ef62cf5426599a22b9dca0e8f729c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6f73e7afd3d5258c1b5589f4ae87ccc965ad2596ada1da32c2823cfd96f0486386c4b4245c5c0d53d1edef325854b4830873a4bb5bb5253441fef3d9f044cb977b9f967d494bc02f29140ef6653651bd87169212b3750cca0ca20875ba289407c9fd578c34bcef401;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h629917e113e2362f6d88d0ef58c658ca6dcb38094c96015781bad6616a12d8c6a2f3a4fd3b0d4637d94bb8a988fa7840e4da1ee8954140dd25e426ab715f4c1744cb37f8143f4bc1ccabc0dd75748316bd0a690d08d6680d3e298b3fee2fde4e6b793ba78466cc20b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1388e2c721d813e044a93b987cd01ac0538c1f963e7381c944f14231d3fde111fca31f10cf619a22f3a97d94a6cfc6da4551b2c15a3fee2fcfeee73b2a20954f8303c677082e26a4172c09e740636eb42d46bd917d4dffdeaa0d93fdb2c884989b17f0fa160c5b63ba0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1146fcc4ba462a6ba70110d2ec2a6f504f22d6e114d31b9edf3062d8218ff761ee09bf1f0ef90312c077fea8adb08f29ae123f2894ef08528d1278731f8f0062798a3a03e7366d44328a7d0200dcce133e1e7eed352ac137fd187f73a9e11d1946afca5482235b05247;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d5081b2801d9b30a326b9ca2f413ffa595ec4bb3229e9c3652524270f972475623a502fb2b31498ba2cd712fd197d6e30317b150c07562480855bdb1bde28f4a75463373a0e097158ae84f6f663c2169013dc389e7267bec18c807ef12b8d3225c8328d67a27db174;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134e40fcee8f1d43c505f9766fd91e36d9689878299496ac9a86da30d4449092fa07cf677923b44bc67b92271265df2193183904c5892eb01a631e8e1580948760e894729e31aa9cef1ea1663a3eb855b31f009fb06b3422b22cefc07c98d35ff47234606b22d5cf9e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186ccc10b350380c10face916665dc593262343e5daabf5cc0bf73244ce3532dbddbf4ffee52e26dca309d786b7377fca74999e6e70c9eb55a57229743bf06dc357cbf99ce0fa7a2f2f8dc6253b641855d5c72cd5f73c4a8c5d0dd98e477a8cc343f37b73259d410522;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125b168b6b03d94b5bacba9915f8a0e0ca493f197ab0aec872a72d19a2f50d0fc4ba2655c250509f938f10a4c417b109d53f9a8a56370bec5459b9f759a9015da5fe7aaeb5614ea1bde20a1eb52a0179e85fc0f473ff8264ef79b33cb5bf9246a1230812f895fefe724;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h255103acc79a4a57259af3a91f82096047dcc1ba1510d9b0fa6cbbc2f11d559f9dc6eb91bf38f5d9111649fceff8c34bbb70eca0d685bcfd676f979bf97c67233b66132ccf12ea6acc659d2a49c8b68794c733ed84078366f7d786d0445c4bd8e9943f937f8d54628f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47faafd36fdcd5bee631969b697826104109c9a41537359fa602e00dafdbf583941c4fe7c6fc15fcddd3229f731eb1c71772077e1e4a95e0792b031928a872373c0941f75f2da87f343518d2483ec3c7e98edbb21ca6c82c0accd812828c75d308f20676c8685c73e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133f07b5996011777b357fc9479be464d103a728339879141ca44fde3ff74fdb2e6135178d3ec21588b6ff7ab4a85367a86ac078d56e4745e6d80b08c1fdf66fa65bd3b2d0c27a5d2641d6a9d4cb4f0dcbb08e063bd2a9c08c11a3f01884c728b2c0d671591dcd04511;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160e8215de4451fc4459f13ac23279b79ef930350ef44bdb78a74a36bede6c4acf28c43d968aee94ee115fa809952742b987cd3af05857def506a53aa323cff419fb1bed12b6bfa69a7831cc6637f8069072562ababbb901cad9de9c4f74a1392d0e378596965b07984;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b87d5dd3966550b3568ad410534d90f3f46ea9b30d000c6bef19f5e33065471dd581dfd77204c386a56d87b5ccd165961c5377a844032e34e5b5d4e117724494958b7a4dc9eabaffcf894aa21070cc717c6ad8cd51bc7028fdb6c525ba2fb8f38daf9220810662493;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58ce46e84ade96a15759805c280cd36d2048ac61f8bb622a57b474c439fdfdbed98c7b6c8719625c60624b72c12aafa698bb91341f982303bf8890f185e6189ce829d8c9b0cc7868f1dc88b1e230fbe61768a79370b0a7e2d78e14d9e8d32959d64ccf956785a1c769;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20690d01c1b4b9b957a40c46f8757904e32d3443f83e1d701b6a390eca55202b9b3db5dc3a041e39ac1fb129d347d675c3562f35f73a558498d86c4bb333b475dd4561a4204f16db731ffbede6e29289c6c877b442502f9ea63c650c023167fe65146a906126f15266;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b62101cac7de06cd3209076f0fe6ec169c03705451e4f6ae877e83e55ea31b979f3072523ed9d5bc5e4d4b0573460415dd26f17cb0a89fc6c2b2fdcfc0e9b0f9b20e65cfda6948bda779ac845cc15e5d719076e01865e2bf7afa20ef3a1d32d3c6711cad8fd55e64c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1274662588e83df43b18950dfe4c11f7713cf7689d3b8c8fd6d5556e7aff38e57fd77327c9092cbc007648a312a49ee6784e9f61e8b811dd342b739819bb03d70f96dd4b811a1b7a12dfa19570974e2e258bbe4452c0dcc5f55deb3b559e2f75177c1d3c1491fbf171a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167499e21c4a37ea68c5a990997a82e073249fda2f61d85d255b8fadd0f3e7c6a25a718dcbb1f3a8c21acef1fe39c1aec08cf067cece6a0692000666beaa0c1f05612487267fcd02951b53917ab05b3865f60e4bb7a2b7f3d832990effdd664b99994de423ef5e65016;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b7ab3c6979432f5e8fcac9c4e7ebe8f18d8f7911e83e20200c6ae2b963a8e27171f5993f1c26a508cd0c146efa4d44ce20f43e41fd8060893ebd21a336a9c692cb49fd1a9c2a459f975c2efa4d8c9a8144a0a31fe67c6c1091963b39c21a09b112214d5472448617a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h973f92153585f040cf82a7473670c380e052eceaeb56689d04267ecdce9f04c3f8d3d906d463546d3fd1ecb733a290d195ab487756756944d0b767c3835fe25c35ac6df12970de8640fcfe0ce3dffc7ac074368f9d148bed53385afa057b4240eda69fad838b780734;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1368951add7c02e7a2c751cbbc97aa3953ef9c116ad1df47fdad7af278f077bb5d7759458c4b0842e38ad9cb35beac8158bf1e621802c2156167d9c3a090854fc09960297d86c877d42a9ed779ef14715d9032fc71f37df03e271dffbe9f1de3f508b97713dea57b578;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3cfb4391d81dc166729ed0d2b5cac95511f2aa73ca3064b7890c938728420e98ea682aa07e43a8d8d825384c3f7f71a5ba1f7a75b7687ba1e4d57c453161d12fb732fd741e976a28aa663f50c8079f66283b6bac1326216eff11f35096feb76ad2a42cbbd066c11d47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eadfe4613449b49baa25efd83801d51dd229aa0f2378a71035d33e407a207357324ba3140bd416a33d43720c71beba9733d053f0dbf74329cb523ad904ddfbe9856ab9aec020a4630b11db9ec8e7463ad41768307ce62992447df00259074394e27144d1649054ff6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ad175fdae5a9150e762f6c038c727fbc8bab1d798c84dc67425ba1a3f99071898419b43dfef8c56d449a151879dd771e2b59c83663694393243580b2b251b84a3e81d31b6b6dd26fb9ba4fb47170f190233be7ee6abe4bcc8d07aa5662e8f3043a6a498b9749dea33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6ebb0837dd7b104ccd95e923d582683fb7545523067a24e9e1b7d7693a6c65b253a37d7b3cd9e1c2c4a4f93671c583a8d9a978656977947d5ca77c9fc624c09ada7bb72080d184dff8859867da358d45e4fa21459b81237c28e0330244429b8495c2464e88e32af8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140744d4495f66d22f6d43c436620d73c6bd34ccf54bb922ab74f3111a6f4dfeae922358c50af10a846907a1429b796253b4c31edf2f45e0d625b45aaff70c62b91a57402d74b8d178eb48d949dd2f618af7753c02353b11e11d738a6cbf409eb2f785cf1b6e2592326;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d3f17b50f12c252a840f58cf1530470d04e2be2feabc52b6d45059f6fa81b5393ee68f25f52ae76854a749d996b405ce9c16c7742e5504dec75cc51bf09801d09919a9882396424245f0d969cad8abae717b7477e27933e163620d8da65ff3187319bf333ea87287e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce61764cc71a9e5527372410f68bd09e9be6b33dc9ae676e72d804b621ac7548e11f2e2d905d72a61f1a4c7de4a1be3b910d2a32bad218372ecb5e7d452b1b100bb067d547f85c428706285b7263d9ec6f208c7627769d35bf63f6d9bb3e33aab6a57cc9eb8f0778d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdffa45f3a646d1b65a698a4c1a0a0ec4d03cc890f8149f5592fe40cb7f20b7c6892887c7729e04a3984bb9f3635215150cdfc5efedbec80a71401d8744ec299829ddab13bb21b2ab347489d97f4348f65913eae5e804f5989c5e2110256d7fc7727cefe8ba26edbb0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfdd964a47d82b88ee8d57eb4d2404578bd43b2e0907c44f364a287eb23ac416074f860b14b1e85260fda4633325276b537f32a1ea2128a680c99fb33036b84cdd3ada04d8d8fa0eed87bc650991e914819e6a3b9fa37aa2ff9fcd8680fce12510860f1e0b9b9e773d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59ad29d0ab72cf4bfcccebbf49240aa1055b06e7dcdb66841692f76f8bdefb4007017e077044f5c45970c99547a601fa503445efafcad45bf639e2f7690dc8ffb07a1d2b5943b2d92b1dc79c2749fe06c531c853ce80d3af9897dd5f85c8fb765b9b337fa54d49b896;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1ac9651d9891ea599f4ac0db5279b53cbeaf4d5248ad1af734286488658f7d4c40cbe4c4e4b2d88a8744f0f2bde1635c182f53a53e6593895dd4a2252ef42c385481967cf4fc65211a61bf541b292d855c7749cc3bc0b069360644aa9a6502c0794066cf9fe5e589a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha996d9490380d8e8eb43aa705bbab12da4953f2eff30e4a0f05972eb42880dadd4d9d2b829465f6cded91bcbac15e26dfe899b038057f0a37bc0c55661716f43bd56546d2890201ae16b5fe30574168c75d0746e2c790aa07efa5d7d59456a3d1a841dadaa90464357;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf5ceecbb88e9711554729d576f33c846925b3a1c53d7edb00c0855b3f0cd52f999593226ac3e06050943f8c0eb9b2e14395c7d720b162cc0290754734022bee1377aa0ddbbe017897b7be64065174d1e64ba91eff72bf5ffafa79cbb55023693e81f3b7ef99c37d6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2841656f3d41808c358537fb6dfc06104c440bbfd48b619e413a928ecd359b2a5ef25f27da07a54c9ff3eac20b12dd59dd8b2e0f7271952b33c72991b3e240f79a202eb33172c7472a837abd4fda2437d987c920925e6a946bfa3da8b2861d8419903f214d48cfd293;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17802fd51a68f6dffd0d6b75135aeb883b295ae083538a398b967a0988082a6faf2b1fe1205b5284207cefb7ace582b4402966ed52039f27235f717dd979888114d6675b10623930808458d45eb87bbda84f2ca26e2c3768fe3689fc5d9b3251cc52c06e573110e62a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5484ef1fa4814007254240b518db2b753a7a7d318830a53be470056a37f3ae143e7c9adef2dd88a3750e1aeb79fb53a326f74c2b82bc5e8378365af4e59be32798a1091702c68bc8c1a7002f2ab7a6cff40c14975f8194af84b9f968bbf2ea9f6cc1aab5e7d6448fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb585db63d3652ea00acad9cbe5534894f477e4af4da62eb72cbb7cf4283dfcb7dd0067457c094559596b682b2ff7ea9c489415021e7a224bf29d5ce07e3c1382ccadb9d189313287fa4e6cfe2567a6a396983aa696b52ef720f7072dd58c4eaf93b0b35fabfe9de65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118218a2ace9f9270babfab219b22a10d7a489ab15e046aff5294847ed4028814ac1d1e4f2374d03b3464dd1b490ad31dbf348eededba95ff64aa38074a5698ac1d1ec638221197bc8f04476be3d1185a7915d858b867e121535679d2dddcd19dc3b55ee9720761f806;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a03b77e3881b381a226f2c371424f4f3f6983245471417e9e014a396a4e1ff759372c8aecf68b4d12eee141d79b341e093a12dcd7e0960366b4641a3f9c6546ccb9777c2ee7b68f6d6d8ea8b3a930519a79f11d90b93a0b8f430632de31e51b8e539a4804fe22e3c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26937e41afb4964b1b4ba3751f8fc58b7f2bdd38f13eed0ef2655d7418ddf868dde533518acb1f0cf34355dd4f4e5e3ef9b63d9be71a80b8c8225f62df9a2c439be2e0a15cfd9d9b7630ce9584b16d8ae4a36d62f09fc3eb7d43dc99d7b8d837c1fdf6156cf3a86713;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1494607f79331818b80af6d7adadbbdaa99d49a9640d05f0980d3aacb6a7cc406639a68575466f4c1e346d80cc5ee4fa038d3f542eb586d127e80802c27c515aa261be9aaf4e685da80e1438520d9f863c871203c11c639320073cbbf4895bb8fd4a5ed9b272edbf96c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3cfa213c0a35aaff978fe2eaffb4c54c7fcab557d69114d1b86021bf9ea902f49ef49e4a251eb38ca213bb2ae38a0fa8a9b57b4d7cb3b0b883845661da0dac3f32d9459a8c1aa65e83687c75dd9fc362264e830d32c831c38cc195eb4e1ad06b2fde56da6097f67aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5f5799858b076bc43750243e3d5940d7755fdd7ca78d18ab07f7fe6a22cac51ac2aa831534dda53c77687521b850f9aaeca093b584e7bc93b083ac4d47987289b2beec6e0efd1db6694c8861cca643ae172bd4a0550e461b019d4a0dd0b46a592fdc6e2a60902f9d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0618ed3c84313461e5494096483c7725a74145d743195be7685645d70c7c5f6006b91f4e52a5c9960e2734f99a88ac9357d79d6e26d93d6c40116100c7ef8e027b2107e68bf30feef804b3e1f0232c9572e49b7f1897f503a263543958de7967218e8bb952c6ec78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e07f2494a7db8d0314e75b10f01d09c798ae2eb6f22cd6f2f89f433ba206308e417863f28321aecdc9e6387dcb5b890c26d6ff4f4fb9309667edb6280386b522e6110c76342df71acdea37023df5f5c3fac9ce9cba82f0cada83f739340cbca8edc54747539cde88d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ddc8442a9f1ba8722a5a1c7bcb82a8c6e9ad09e76e27f5fcb4b081d1ef814adcb2c57dfea7a974669b5ea984819776016a8b30f6418d4cc69c0883a0814b23f45a744c707326780e609023a7b78b2268ed1cd85128aaccee3d43e8213254a5fee2c91c849e489e207;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b4f6cb685b07dc4e538b9a5503a121308892d924704795601f4e85edea564a9bcc5405b1c56e009e30752bc153a3673510dc18cda7cad5da8bedbf5ab7d5d7970e65100a10b04e941a0f4d9e9469be27127fb4f779a103ab590b91fbe15189a35f1659f5223f2b4b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1795afd82476c4dc2aec4e8cb3d1ea4c5db2bcb9f012ecd182251524f01596b9851c4de8b0e73d1b5b72db0e6fbb5e21259a59e6330aa6c9c1c525bf46d8286031fb68242821a032dd7fc05c6c5753ff08392b2a25945567c0644701c2194beaa03c3f5a4a35184e80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab4b76a713840eb095190f901d5fa62bc4bb11724bee56575dea33120b1bed5ef6ad0ecdab1681ff0800403d7e9eb8e37af9758785734c980a35f91b3cdd8c82ac0ea8263e6cd892a5ccae366f2ca4d84f9c1d5f4cfcf7dd565c13102b2a3b1943167ff74a868bebf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45abc748c5b7f2b76ce72dbefcd9cf3e62bffa8796fd0c8d54a7d8feb0cb347fe71524dd4a334c2cc9dd011d59a38e57217ef34112515e802b9ffbbb94a326e3ae81a38a283d47c81a76a5c4f7459fa0d27991d70de4f4f990ea30bb058d3a8dbc809d650d76265b02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b4dbdc726d607a4b4528c96ead4bd482dbb1ae4e0069de8f2a7d870508a9492a87ecd9b86b5320b248da06e008a1bbac9f0202fa8f52f2a96758f188e055af08d452edf6722c74105c75e7659a4b0e10a2bc1b0acaac93c9e09575b4225f53f78b760124c2adaa903;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb68f93f5133f610351309ca5f9659933763d208ce2c577529d17768e2f59ff34ffd30a1003335e4100752c8fb02a2f51733f9eccf9d982a631cfe5a1d27b141b5419cd5f8a8dd5afa6bee2a3f32a5f9a43a7cca10845430b01457b8c0bf23b85b405ea8530cd74868e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15377d5cddabbd11278e1f5f720f49d5b85a66051f745e9a33707fa30ff31911be56cf3e361aa1ecf7f8beea4f3c303c4204fc51e95b07b24c4e32c756aa34346ce4427081e6a3b9387d325e01cb860fcd77de0ae0ab6cee78765e47bf4dc146bcda4fbf2d3dd6b0926;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8cea788d5c32650e17206168413da16c27f5e0b8c0ca1e77fed207e7e4fb0e8b4ef22de786c919483ca83d484783209844e5f5d56dfb7e22566f627e15112d263dd114a0e9c07616bf492268bf99bbf5c4aac102d6409a1a8cb867e07b7689fd2646bf82695a3f4d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bffe6927f77e323d1fac3b8ee5d1a29ba8fb84f69e119261598da0f4bb04739889960f86bbb951bfaafaef704ed2eca0746c2387251e6f20d6341218e17159093d432439790d1891b428be34c6e4acb1d69101aa0e3736b476f46c78ac72377454dbe8e1734a45ce14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122dbf8824a58882f2e2e3821935f6a5a87fad6b5d3248f0e17a1ef5fe8b982814ecf05e037125f41702f0759a4c266a031901ba0c4918d9e398a50f354cce5a3d4db9962e1854f61b27b220fb86e4a336954c108590df2e402babf0c7a020b6e8ced20d54b9bbc3bab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb496d4133f1371418a80de91450d197d047ef0034c7cebeb031c52aceb65cd50c064e608a6759b2ff1c7173955e2b92a0d068585b52a38f417e619905857a75c60f787a93b60320f778163179e6e2ea62d847fef360e4f98572fabbc599fed8bb6968550f029cfeb25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h500646a89f18a0ccb6fa042a627efe2c28cfad1f9e7ddf8edab00ff14c58e36c61c02e30b27ec3dc24f776bb421ea312bdf4f680046ff483f94d35dcb5f94200a8d6a2e86d7a418e379b279fd9be836b5ad10ab5e5e213b9b00338808a36cb5515c2f21fe590e34e4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h541e36bb07ed49f28043e8111a37f19c53ed27801faf0d31af8db09c24f06b23f44e498935baebb3eb48e0bf9d77f0b8f5aadb145c5d60af5e2f2ba74c7bd0819fed48a061caa343b8bdca25a80dbea381ef7a88690d1fd2a5c7114519ae1cf18e3511b1de6c88faaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108a8496aaa47c8645c7a3df38e5ef98727011cd8ca56fa6584ddd297df2ef5a0a7d30a53cbcc3d9c645d89c919d937e21df858a1af2d0e18d96e97d68697242bc32a53c2ddebfafad90dc62457fbd09eea280bc5c1b9b2d77614c319c7a4cbbeb3173932d3dd4f3023;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2cf329a1c80e281343cb61b385e98485bb297bc2a8601e0ff3b697b04ceab8992a4c9c3c7f9f59a5bc18e00267a689c42bb6972078347335cfe13bc52ce27be92887fb5c4b6df21240468cff2a58394946c9f6fabdb713e6b58b87d23c1430ee89fd2373bfb9b1375;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1ab830c070fbd8de1a1b99581bc73d989aadae94acbca04783234e4d2bbe4541052494d4f5fb8863c6735025c168addf097fca048917abd789ee6defe996b92fcfae4a6cd90cdd06bd39bd8dd0862e28b82d31ba46922ddd4da013c9af911ecf250ada916ded4ed5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a7eb443b73b5379c7f7d93d6bb79502d36957b5973f0b78a1c6a84b7badb375159c1f1f52ceed42058323a36a77aa504c984ac3496d2ad926fa56d440dd9ba52d6f6ec378dd84fb68cf00190678f3b87b4610b2e83ce092e16993abd282bbcd8ade331ebd9a7c6e22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb1ac8946c740579221cc388bee39e44b1de7b11602b98f552bb0edefda007397cf16e97766514c3ee06a4279a5e8c52243010b4a943e15745cb61c96fe12d97d3da0a35b824fe1be74f1a574d4a3a71ebfbad6ff46d6f5faff1caaceadecfd6fea04ef9d9ccfcbae4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11438d51a6e0ac2358fdd63256b74b91d8421b4f28b0f13671720101d8df9d0d1eae84a8fbb8471210f7e1c357249610fb37c63db0efa969121ece2749f83dd5d8cde1fbb0b5f4561a6a2ccac763cc1c02b48c6a080d0030835f32fe064c1a3fd79bb61d8720b660b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102d45b31d5f56df623a8e70d6e03f9fc2c1d3a7653c34263cd5f540d2418e7727a9eba2628334af0e9d0671defeeafc5f4b5824f9863219fc8d9630327f1fbd064452ef4f235545e7563ea35ea4b3268ecaf715148309a93b08bd88bb48bf826edc2015dd90ac5b6db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h29f3c0a3059a45edbe789657bd6d2b0a6be606f5e7500c47f71c84ef5e9e8f102d61a26eb6dd451b78f0c3241ef05553ab12226de74fdb1c44981815a6571457f66bbd4c15b91422a7ceb5f6c887401637a6cb5c726329c7d1538fd58b34913522be7a9b34fd64e8bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8e04a3535e2be508e6d2f4c774b999a8de366da8c86b1486fec4948bfe3e28a6d7749f5a3a853e6ca2a120cc9841442bb7e58876b18d25db6e12a33e80640a9818e89eee6e07ac3107b61ebcfdfc3ec13067fb1ae0300fbee61bf0a69fb793136b8088d3b760e0276;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7cb445e3fcc98b5ebec0feadd2dcef43c02036ce939bb56563182f7d3ca53c5d4f52028fac773c11a18d8195cb49cfffecc4055bed3bc253f2a39dcdcf74ca2aedce0c410ba9538b3609b8b2cef55517c70d9bb5d01405a326ae9588085b0966425e74b2aa0b63b3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23e1acf19726f3e7369de443f8a2941ae561c5073de65881a3481e3359748cfcbb10e59feb49cdc10fd0ac38ab270d3835bcd44355022af6fede668d778d8f46272c62d92cb27fac0464d259bfb887b29aa9b3b728dc9ac14131f452a76de671c463494d76985f31fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2ce807a9678f22aee11184569e99d6b328ea1e17cbbe01f946d9f98e43d85cd61e9ef2a628187fc6876b2d5fa8365aac71f2a7ec6ced879038801107c38b38688e8b3adcf963d250c1a7058514e3cb984d4b95bea53fbe663b016f4a5607f9b517272840b7c79b8ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180aeb68c7a1b87182b2cf9f5e99856f57152996b41129d5831a281bb6d29fa206e529476a3e6c120c99f9ae8b9b14914b8fbbfac7946c31863ff2d13295d698118078af5abc07a5e30371ed1beadddc62cfbe8176511807c81f17474722681cccc5619ba7e49ec2c59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48324c33f93ad8988da462de57f73ed7b6bb066ccd7a44634df439684f0af6eaa8db0cdfa2ec1d9250ccd1546bf0a9454c3cde6b3c8a3ed669f3ced3031157e328835fca25a4af2f97e488aaa7dedfd6fe90e482718fea67c6858bcba8b3aa069ef05101e98df2b30f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4032b2d093ddee5f64041b9c12b73dbbad141d2ee684e545727c1c425d97f2b463dfdc9b76fedaf6abd12e56127b1ada84ceece82e69fa208725be39043ac6eeaa9a513a29175754545350fabaa22ff2fa35c36672b1665592cf22cc42805809a0109b4f644553fe7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba71c32d76dc6590908936aeaff0f5676e932aa38becc4f8a76f130e6ae25e0d53ad9f77fbff05286a5b80cc1df079a48b6decb4c814ace8def81498c98867b16833da73557e43cbefaa8a93d3b6942bda3e2ce5f4974b43c11712a4fbbe1201ce2beb79d57521da51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6248bd11952b86feefb5aa9dc3597e1f82b30919c9750ed053899ccda0c7a995b0a7c30fa86f0aea845258265ef737c7189ef3002ec062cabadf9a813a6cdb8d08c52ca7806d188048f3417fa9ba47ec003e6c7aa3d091b1e3264ed8190c6e9daf8d6e65f7c9341b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfdd34634954ade7a6fc8a67308c1f17f7ec947c9deabbac0dcff002e4ed37848438138afe433f7f28993d2197ee54bf2b137e4d6d2daa0b0b29daec0d0179b8c68094749dfdfddc8c890eabede6052d278453bce44bde034bc750b4eeeb858937d982d5863da0a14d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c88b8bb49f15244ce75f13a65e5a3addefd8dab7babf1bd49b27d5841450639c60aa20cfd450b95355892ea308aad1e319072a668c5d7e0373ba22ca9fe089ef1a0549a937aea7364c21d6dad4af817081252556fc9467fb9d7fb786263f0c85b6bbde0f863b376c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b101f987f18defe7d2002b2c28bed70ca8be2f8ef9c0994e819c1c272e9adae5229e6b9bd5facff6cab1a74eb911f708853ee5aee19a1e599fd5d5b54a8b8f33a2d4c18b05763814ed1d2fe95f26a34f8dc51cb8757bbc2a2d5db1097699bbd613b189db64390703c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8f5e6578f943d76e7c04a4f8308525950a21cf8d46968d33769f4ccb0171e61fb3aa3954623bcfc09bed518f930c05e4a7d3040f7352822e6dfe66ba0dccca7836fb305b5a6407debf9f4ba7ed3c8d4c4bd0389d7a992946598685e19aaeff715237446d2505a5948;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h139cb7c148690687c69660163452b2853947c5b689f27700864135cea3ae67d1c6420eb5ab0660981da0c5ddd024c00612d80160c2860bcad7ac18aac76c28bb3cef5b2b72e74b8218aae459ef31d9104378274ddbb51079bceb6249105c2df1169efe9f4353acb4d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6a8ca70a99119bf9ddc1ba3019c99f154c2262f933ebb19af942e24b2c175affbf05e117c1482652d7e6b1d17089242594bcba99c862885eb33e238a405f7bc9f42621a9f2164945010d758dc597e0a75e74e7c57a520e5b3b8b8e8d1b3afe7a3bd1981dc6f80635d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb03d512b25631681d8ec571916bec442bdd88b6df7c69ec7bfc91ffb630e6491d6fd68252f2aeacd986dccfcc03f3598111e0b1c7f2aa24809cc8ec44564fe63484bfa22ba00a12702f036aa28a782a82541d2123b86205f5758febff68c05ebfb448889cb28cf91e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4d0348a69c8eb99d42d09dbc93674e25586f1600ea4372be66770bdc9a63bc6da85403b5d7810932b4726ff07d954c39d4277196b3753904c2f6af42fabfbdd7e4a99d9bdb84501af206a7e0c56ce707cb8eb62bc47803de3ef6fe4f9ffba00f89d04281c9c396358;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa9236548000fea940c73cb6dc68dd6557777bc6dc5970843786177ccf3cc8b8a6bbcda3010bc3a7b39675f2f673bd90c5f367e83f6375aa773065c0571b42ed57f2c532c6d3c8e292a6d654ce1911e9491518ff25d7fa3ae5904fb1520c5457a9d670996c0a199ebe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d4a965612067dd028db0a54bb80166e15b2fe2d5aea0b7634d842c9510a24fa400158dc55203d1c59a1d44d93f478e41d5785d8cb49b8a2921ba8c5f061ca842ba26c746d1433aab6c71ef62567fd6919cb6892ad9386183f92e1f418675388c146b12810c1f55252;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f042719bbc0f77ba05e01bb1759c76968200148a0882d1a9226b0f114197cd4d9b890ad92916c5e32886bab145729ed80d81a693e04e64b63faba9eb10129b8ae632d7c4333902417322f64fec2cfd20da9c9a016257899c28d9c3d32f07b1dc0dc78be278cdc14c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h364641d81c6bcc9e5149e5dacbc82eb8cb1bf392d8b17294f4ad85c0cd058920f63551973cb5674551f9f24912d3daa2d6f7dad0bc375a34741af80f7134d4404277339c69b53d6dcaf4835626009d9ee0b4d92b029878f8dcdba98fdfb119c34719930ed233c433c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e866b5e60ee4dff805b725f3b319f1f703d633def758c6ac98f6577f92828dd6e95491fadc84ed6cfaf5e470e75d96abe315883c6813d1c714c7113a624913f3efa377db54cb15828a3b8fd52968c093f348cd0afc7cea9e62ca2ba52cf9a0f7173a126774f037d41a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ff066ddd2779d4c5959f43955b3a6949b6d4dc71cf8b8034ce4a2c7aa39c4d3c05a1fffdcd16e759f4415c91db88316d9fdbaf9138f8c73d0cd482b1295156238eec1610c9fb482c3586e12114b83677b5a72ccdcf082b3cc84ca85b63c9a7c7460d934164409d95f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc3ddf099e96b296e915732954fda338a9d8489ddfe2b5c900fdd1b7742ae2c4acf6aba1d2d41e5baabd9e7386da6ceca568f23c901955d8371eee2e383905fd8625cc2e3d43e4951de72d59017a4d3924c9317abe21077c6eb99b716b8e2b78d7ddc8b5c247581abb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13117971703ce532496a00cb9ed012def1f158febcebe014858128f3b79f0e2b1e3bb3c1bcac1c7956b88ddcc49666545109678e11765478f00d07c247fd9e9122e697d3131c508eddb00281df085263d0e9ad093002cb8fe544dd6af735d87daab869d75bbf09daa75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15eb37d8b462953bceaa931e9842e49886b64f7164724e23ed221d4d11c0300fb3fa0a3ef1a5302bcf41520cc05ea17f411402d23a77f27010123abb38ccacf6dcedbee4021cc6daa02ed23c9bb01801f02927285473a4431600d902487256b5822fccb45af5a12101;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5881089526caa0e2a4c6828c8eeab8e9feb16cce00d575f5f5081264dd26d02dc9175c406d9fa75490e9f1163fa7e4317a6fb2b50e108aa029ae5b3018627cc57162afce947dfeb43f09c93c2952684bf700c9203d5b547e1c4d0ceb04cda90d11991ba9243c8c24d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79fb1029d6cd4d2b2bbdaa5699fd16b98be141eb1eadc5f8549febbf485e8dbb64d3ca2cf59ed5b0c9f906883cff57bf1a2ce84bd30507f041c9c3879d27a535bcd8f857adbdf20bcfcdba628abd65a30f4e9c0127982d55ca500472ac7a73b62429046578260f8e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba3f29ff9a2d7f1ca201e35022f28b611b2192ab235f700cee47625e3f190b563f07c9602ec32aa15b6cf8fd007a9f939ed4f407657a5272f5395d22926e61456b926a97fc2910c1495c774708bd3767863fbb791e3765aac669a9c82acd96f5c5bdd883dbc19224d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54bea4c6925b358971b0885e548f3eba71139f044e3f249b568d6c7511d2e60446dcdd38df7b50887c67cb7489d5d46a6950c8dc665f3329bff47e8246d808c8d4a1055d0c1636b020b7755c10635026ef87d8c7e1224130b0b2acd60c3f8d270972f2305d88cb873e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0bd06e6b6912049b0396ed4f21781da66e77c3e787033d6de7ed1b4b37fe672489aaedd7012056fcec2915c6b4e69aa46895f09ef9701cef5904d475a4f4b2ef09fec88b0a483819372c96f4c6d06144e1ff06db92c6cec97d6f1a183292264f24fbdf7807b00d950;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd4b9a310024d77e0093752f385ba7d32d40e05e7b14d1a3eee314df5a08d83d584d3ee302343051b49d1784674e6f91d51ce2058c2b97b559c505d8e475f297f078823ced300fd1f81a7c7897f02c7bbe7cff5bc109fbd42b214e37d8fb8875884c0e524f94452fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf85276b913b03e67b1765944a58a5abfa57722feff4721e8dfc6515fa9f500b8a805331360c296a302f058ebb46c9f1c53979fc802ae023fb9d229cc4069a9f011a8f853135a9f57a30405dd1ac33667e4f9a979f585738c313cf2ea2a0b2add4e75bf4b7886f1752a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161b0b4bc846e795ca699955c5f13e98922d7a8f7cfd604a6646b9204ddcb56d6c4de88c8173a69ee33aa7aaba4e7614a80aa89b925716a3ec50c8a9e049c485cf962bc1c94ce46f1fc0924d285f438fbcafeffbf51097af0ac54c815626205b0d70c95dbe6118052f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129773554bd7908e3757c7b00849e95620790cbe9631338bafcc0a0a75e23503176c2bfd55278c337af87cb786f0f28bd999d9248c6362885e1e27c1220205158e60a30a77b016e97f79ba2a812c53e758b9223070a40e5ea3bf188e6758f6e1af609edf4bd4924718d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a66d56b9557bff2640c964c788113eb486895e68d514e5475de6cf9319c8c2b9cd1e80f788f8e8f33eb5fb9e432cc34faae2ddb3c3f1363f32374f31f4c884a463581fd71662de676c2bfb6ed9ed27f49db75cf6c972fbd2b547e197b0aef9b4a46b74dfedff6e15f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66e1820828251bc9c0fa62eb250b1072ff5ec74081e03c405ac1a0b9790dc2deecd26ae0769ef352c29158b1e03ede7aa6e2878f01b22304ea1b61409c56936d750b1b143232c7e3bc18baf65d1506ba9fa8790c836339e3e8ff1b296eebd5af410c9fe030ee33cd91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87cce267a990dfd6e41d665c6e2341a4b4485cd3caf2c1b4461b8bb0f96e18c33d350c789be768d9931574ba16dad67698fff52fe76d5afcf3a194dc58c8a57efb019e7c019cae7e543a8bef226e27691568a24a60d931b3d98130a74dbc7b6ef3ccd26916a1c1d0ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12290048cca7c77b66df064fbdd23ad4ed6dc49afce5c95e226320b6bd5f35c43d51b06ee1da657877ebbcdf5f19513be09419221badae26c3fc42d2b8067679541a51337445ef09894e8cf25186b4cc123d9ea2ab684d622cbc299aa5459d6e3a9287d5d61ba922f00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65d2b4ade3362682c8d08cc68c7566f8d4adadf309b85810b5bea4e64f067695dd586bbfaedbdb3329c8474f2eea8fe11c7a66bbb183d598d6ec8ba2a603f5c701cf9104ae151ec37ec7415a5a07a53971b7873c96f89755cd4cbffb67d9949c616e7735687021dc9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d1a3ef8d6a91195d9f6a2f87577f2d69edbebdb6862567c0dceee40f7d086ef6d70e0b526265e69fcd1501b3ff4363f2573f828c6b012ad6b3889fdaa50dc1dc284e3b1d643878475e90ab05e4b76ac7ff4511b16aabeb98412a3ac0d8f0b29f8af2a9144415ce843;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1277475db5801f3d93755bfb5a8b214098ac458ff6ce09e6140379ad392066f2ebe3a92052c0c3c1fc8356597e158972f6acc561d38b0a95b2f2ffeef146c5eec6c6d394784198a5bae660e145d8df902b647932fd5d54990d4b172cd5e088c0a9d7c8ba206c4cf53eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135562cbcce2e2d7eb8e1b3f5d9bd731c89ccd2dd44b9ee1633489b0e1fc89c722d691b9f32d3cff42000967d3fcda74236b74792c7671c3450c56718e7087b654b9ec3b1eecdf2119c3478a50733d07afc1e25519389494bdc9d9bab97641faa50fd8a244df51ef80f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fa829a7e811d0a76648c9582d942a5b756da90a7d24a46a3138738419d98f59b615a035bc16b2b72d55387abb27a8acf8b8b001df293c3c3dc8c2f0bc65ce7bdce6841eea7f22449317c907d454eda2008762c1751aaafd32968e2a4aa81df3f3357846e17ad2d2e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f19fd78e0c597e534673a69053e83c27072be58df475d70a9e35df824248bcffc63f9baf57b2d2ea3879e71d34af0a433c07dae19feb7ef21d233d7f90fb60844f545846788ca4f8d9a2b7d1a10ba9a9cd0ddf15fb87e5a2d026480f479a9f95cd006291046153059;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8dc9f4b7ed13199222a0950b4a5d202c210a1a17fa8d2a65118426cc006be947819d1a0c9bf12aa8f603f1d349da881b3da400eed42821c4012e5646c46d22324bffb4a5741f299793340097438a7d8f8ade88097d3eb431684bcd6def1e40a8c2130925881f454a4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1be12f2ea2a60208e2704abc22770bc50255d963368ff3541bca381347219f09c75fead6a77b20c60113285002f676ad23c7de5317799f94d4997c6d88cd29a11b95a57e86138c475b573c3e88d8d8321ac95216d031f0306e51f169219d03043a5412d540cd97ba8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174505f64da2d4b6ac157ef8191b87c3f57e14fcae1930cab7b11de7e7d17b440b4a742ecef887f75fbcb02624161474e153ba75144dace72acf1692f99152ceef0c15345e830c5e933e79c15b4d1b17a17b4de6f81f900561c4f18ce55bf30f1c9bf3f6a402017b633;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0b5431d503e3bef4f0b90d471466affa45d605f73ef41a94f3d17cfbba7556b9757b258fb6c88f2d90f8ba1bea625c9bb5c654cfa9f44fe8752512a3b7af75654df76db116b0c26f74a7ae70fa7e69da696e53d4060fd0c88ef280262baec62b614071f76f8681d6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h244fcbb79fbd31ea5da413d5affd8e931edce12fb3a4b1ef1b02ce2c624eca8797ed2e08f8f4ef44b553d5d8e1f8ee92d5b44a92e89eb40db9a98951f746ad345f150bbabc66e77e1a1218a4b6febc3dafd1b3d482f8c252c6fe8f96d088e8f17412531f12dee07e78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b30250eee36e865728f6366b350c60b775801dd8b0920669469a7fa3a290cd46d17d111d126182791647a67dba94bc9804d53ef0a8d8043de5c0b7c039f76bd5580b59d733ff70bcfd05eb3bfac969ff3db53381967e71d77eb6d49993b31d41a30aa1ec03d791c5f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2152b0f042d5e3d0ead781779affa57b6a15026fb165d59f5d43640a0e1d9cc1356a221fc3f61605cbdbaf79627ff3653715e6a1d585d4ca627980919c5e41649eca9beb68dfd0dd7ae1c28da86c1d72d0168244bd75cf2c7b3ba4bdd51adad99bd66625079d8d024;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18dad8a342594236a40228afcee3d39b00d5792bbf3d3cc5c18a1365a1e69ca5e64c3bc301b237181ebb8b87dc8763e9b75c40139ed9ffa7a9d0ce30f990d0a5ba7b3c232f5b4d8a1305681c638968adbab15fa135ff957768d7a7769190d035b8664cf8b3e84dc548a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4be89af4c5ba091171c5dc61f70084ccc6192987c29e61ea77656ffbbb61b59456be91392d86e6973c54618e0b47c0b07c2b6e990f78b82258f3b92ec37623b6d8a313e23ef7fecce11896da96a8a59de48698cdeb9f04d671db4a3674abc3f2414356c5d6a23a7901;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa0649168e151be28c9e9c36b485d4a2b3ed009f5d4eec582570841e713deea5d9042017a7710c584ff34807442fd1a5f6837d4efb416b08234910ca55b6ba0c54bc25846edb0dd8b8616d9568b9f63dd759fc3306c7148b60b9dc457fdbc8e4629468c9d2e563977;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cedaa47e29afa455730567c4cca3397eb0f864c108a62dce69683c345a501d92a2a5af3e4feab7e1739562da8281eb1aaceade1331862efce6d6775ae5f00bbcdcfea9a34e3780402625b461f9d50a1b2604a4eb0d8a0698c602d6089d5e70e6bfb7a8b4b278432d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8f9ff8042d89e8483de3db18bad978f6800bdf881bdf25b6cad3bc842022db570c33baa1a7f29c3350512382da17729a31047c9aca9bd11f38587c1fb803ebdb437ae27fa50a6b62b59d839de40a36a98a28ecce117e3dd0dfd676c83c2c94c7ed3e486105299a7b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8b3f3b0bda06120731b852a3ccb74c18a95d422ecab1d89c40bbb0e8e2ac7e2431e93fef22c2878d8042a2378563170ffcb85d09e6fff826b85b2dcb7fd297a148af74255eeb94560ee87a30cddcb688703b55922139de90edf7e6e1c5213c749aaf1dc580c8f0230;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b159efee52008a112cfc2d0950859621e029d9f0cf81d41ef56ef008009c2dd5731188552fb97b20599a1bf4554b09e304b8d05ae4c47765fa28c7746a691c65176cfc8e4673eadd21fe4243cb219eee2ba02b7ddb7f567e621c6629fc020ed4aa3aff9cd6a551bdb2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h387886098bdac21296c9825b72ff7537d8a1b1906ff072d012c0ca10fdbd5f94762f7d3e096068730b900e3f13c8a271a3b43a515829cbb6c7b92bf246cfa88f2ac18d171cbeec9f9178f8a684acc9c0120661618994a4cbf08e4f4e71b91c95592e64724bd1673853;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf518de197274306fccd6d0e618c88198d9e73384e791318290e9bc91f281498d1cb1cf72922271a25b8094b24a4363b37510188bf13a6b47e15ccca544cd0c79eb462bf33a9e66fd0d9333397d1300eb676da71f326ba0e79522afda20aa10d543c246f760f0fec2b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2dc51a9430a8e6dc42c5309c62023f2a2aea57a069e84b37c731e4d3316f2788ee219b63709df5137ac0ae14498bf38bb3649f82f512a956d8c8440513f7d05a569003579b9f54849d95811554b01c58c0773945dc9cdfef922ab5ba03c39d8c0b5cc0b7dc71b8a043;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154d8a0636ef45d4fb5d24257d3dafdd74e1ca014eefcf3b1c9ea7eebab573063c63073921132c387aa0399c2b8e59fdf733351f0a13def0e61c17dae4a0fd022b2316ab6dcd4a9f204b21ebd31aa338d1ed42af23ba1634987c95d7acc94b6d00f902faef3a64c1712;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159f4b738d4a4d5cffdd6643cdd9abf64b0ccf3e46d6cdd3d425e3facd1eab09fcb9c8a4583918efc107d8d13436e2038ef40d844945faa9728aafb14446f638d7d3cd11cdc03847e003879a8790e1a51d1a077a670e136d4c22a24a9ce2c8a61aba65a8b327f7a6db6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he31525b12381c98fb6164a4d1b11308af4c38770048def93f2c90c45c9921a4c0ff1520f8b366d051091ec28bda5848c7aa204caa2fd4c985b59d75e1c1508871afc9f88a1a50e9d1c4ff48c6cb85cc18082ded9158d2240fabf86a55fc1e45d3c78fd41aee06ab0ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc88ab42478f1b0efcbf672db22b6161997e19a4b47c0a9e9f6e4d8b1426e732c4ddbbabe7ad4b78e9d0f5c74630f92d695a6ed6b7b21289eae4b4928b4792666b2609ab5e1d4ad0f02ffe44a960c21a48195b142e4f96fd567fe0a97fbb60d8af2e2bbbd5dcb0dc05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160c9e820e31728bce8547851829dc11972929402d462c923fae25c8864738b33503f51af583e1d93289510c3c75f87468d3c1a6107bc203911185eb8780e9ee9fc07b1f97b94bec67693e691854b97871f7772ed981d3d6c9e5d17bf5ca5ba6a589f2e97d11686772a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bef540206073542f0fe3cabe711abed56121250c7922519932078233d51d9228e425739d7d50da4d8b7fb91bda9d97a82eb8c97260abda3f1aefb7ed98df3257dc501b3d5468b17c301821bd0d90d2c1037e70ea9250b0bfc0058f6afe8c641011ee16fd24e9a7918;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190f2808d31c65cf5e0683282fba1da4f388e49618bfeaf2fefbc5d572c4d6ac9ddc74964c2051ad6f20ddb4513074a199156832d492966e88c73b2ea0707363308b2c655cd0270c43a027cb4613114f1b2462fc9ceef860e9e4477f583b4d16e77302e02666a765019;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90148b72121ab1caebe0430fbba0dde799755221a2dd3b88225d6bbc9ae119ef30a01327c5f898376ec4a6c62c1017ce0163f811ed2de24c088b6b418733903f00e8446b79142d5662f89e51a58ffb5cc55ce35227f276a5f974cb0afe923b0bb4bbc516d8b0a32cfb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6b7830b4fa63e9d69004baf1f592c4c7f126433dad7568c132116ac977415804b4494f6a5cf7abacdd4cd5f2ce2756ac60bd3a6e864c087820eb4d2dab1be1596913721b65294c07f315955725ebae88febe15f388136711a3704546ed96f98d54fc6a4a2d2bc5837;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf81c7102a47777aef76c182a5c09b7f54dc8aed13bae395982a0770f8fc94887cf8238c0ee64f01c84f4d305fa95abdfc35ca0f96e129ae49ba5580cb12d0b3709e97e4310cf7de94a3656296517facaa34dde2968fd28ccf9c633e16ca85a49645c1e6603f31691f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h603a07faade92c2441a782c338e89cf3cf93851a5459338e42207d042d344b3cef5f811edbb2d3bdf56e608eabc0754b1e93035db9ede8e500ee8a721f94f9bab2935baa658f08600a578574e66c432cb8810e64aec4030573122f6c4ef36d9372c36bda14f76e2ea4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141343814a6e28e1db4078f315976f95bd1a06dd79a66e20f4f794e4d4f3b199d3edfc8c5e5711637a65a6bfa29374b036db5105dae1854d3cd14b1c1cb13f268a2bff98dd7e78cf71881dfd0e1ec4c638def864694ab8ecb42e2b70ea8ff4156141a8ee6bf8c3109bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8ea57e4722676f8fbe45539acc147281046a7860cc675add4876543de64f496c66aef776fcf5ca22c92068273adcf9b0e2e1283a6f5e6444439f0fb5723d59247abf404ff1f79afb978a4e9e5d65cdf550395bd239ae1e0c80258c1448ab39e593d924ae7534c6b27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17df126ee5431a87dd82945cdb3ae300ecdf0fe315ede333bea91fdc59b57df1aca5083e3660dbaab05231784d39177757a9124e94231a65955cf838469842b2711806f73161a4a11c0fcc612e54082079a39c59b3ef87b467ef4281a596fc20ac7e79e3546465d453a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ab54c2aaa2cd6feaf6e151adf6bcf65fe83d94469b889d5e39069c9d0a17021815ae9b2c2043fd9f5373a5e48fc96c322b273f4a6c6699192a1e4b515393c9c919d6d7cafe5508ac61a6bb63a613995039cdbd8a3898bdae0efe7663b6a1e130e3eddf5de8aa7c920;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17cdaf060323e9fa140c96ad8b97708a8cd2bb73fcf93308f31b151e5783fdaf41b90e066e263166c80ec2757d866e0b83a67a592b2967c615cf38e68cc3183c16189d113b5cf491217528a7902c58a25e35c2c17384a21cac71be81421fa10ac4c7b7e7e4dc98565ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbfac7eee16b067d0d33ff46fa2008af4d7a8f524c74ac55ef73823cf6b96491e67c2b8518dce693b131c8093f2e1cdbb052ea14b54ea7d3cd906c79b90eeecca5b7a641fa6ac94926a4a99d97b9a644f2e163726d8fea702094e87414b28f20faed57004538215dfc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b4a2d2d49a0244681c36dcdb08677b4d726524130f53e45995912350e8a2fb7a55c4b6d11073241037a8d35ef39caf479e858e1248ce24f7d08868aa94cce1e5a408d4bf3d09670c05e47228e1d18eb149bad286c7074ef1c10760d81852fccebbf973d50dec9ade1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c39014ccd79f01fa621d531638c00382070cdb19e79a14403fde8a3bbda10035c00a9c9060d1e4445deb62fee78ac80ed6e7cb1496aba65c4fbad34b3e46770015d57f9993750424528fe36334d4c583a009811a0f19a0dcdaa91270e5308e9e0c264eda067f079628;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faaac4c54c2e8e1e35b8fbeb0198f50083da207cc958fe6a5ec13e860a7b384c7c6b594ffca74857d867b8b85583ec08dc00520afbfd141cb2dbad62c9a1c7af2c0832b73685173d66683408c2844df8c74ca5a021a2e5808cc0d696b737d365871bd071f9d0c20d3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2f8389c27e0b2f1b0fc78e5bcb7e6f406574071f56bfbc9d51bf5c2cd4a796062c9093b34e436b10220034f800d7714fdfb9072aee1569a96a59dcfd2250cae874b9a6c68cbc1f92c3679ee19e1014b89498d4507e171079f9cd268d1602dfb2b73606a884d2abe4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf71d00fb7c266e83d8ed954b2f10a47718cadd3df22beb965572e781a1eb39e8cee4e9c5f09a5f01033dd7f415c5742583be9212b41782db3607ebca180e6bf358698f2d35584f011d1382eee28cefefa20810957349cdc816387b6b879270c7ae4d3310cffa519294;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd2996205d38797864ec6fbb0f8c72156931c76d509d8e3d94a63012766332d9edb3a855f0eba613cd279d665569e8ea2a90be72eeb5284b649daa0b7ec06fc3341c886fa1f58055fc4ed9299207e78101f5868f23a8725c9e277d4b884c9212a30f885f6d82767cda;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3fc8756a15f74d257a05dc3d093d6c3e43e2e418494ba2e760852c5329632c4fb731c26b2463893128c09293603ebf367134f2d909861f8ece09a43d673667d158425a77ad8223baa283381e000b14c22bee25950c1d41308ead9754361259d003b4415fca335af71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had3dbf674c1e94659f5ebdf434814e537663893e5a6f739ff7fd392c11ac1fb524ac9ea8287af06a8df7253a7892a155c5ae680a159c197bb45b7bea584946a5dc08aaac7942bec4035e8f6d0cdd75fff7a6d2aef200564fe6b575f1d966dcecac0ce2c989a768cd47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36b34b37fc2170d0704a56705e97059ffd4b3c66bb59ae89fc6c04f430e530645feb452189603b95be7866ec76b98d81c8faeaf6422abce7502e3bac17e9ca3a01424a32abf2315803446ec856dacb12466730dd23f47436e5214c11bc91334c7bc8ff468340929e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec06252207f0b9059291d7955bbe789e89505c38b3dd4bbf6a35f436e04e64e80b627a1b25ab0b70b1bb7cb13f48406bee7a2aebba14bc6c0bf273c3509791fdb8af87e07f13e236fe358f2f8190e802eafd0919675793429576429cb18d560afd6b5fb618c22acf54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7f938afb3688fe991d6100ab88844f77ad9bf3dba61cc533ec321add7e7b76a4a8ebc4475e50128469bef216c31697da5ad16df675daa9da25bfb7ff1642fd60e96d863fc6ae39570c394d8efa55cc9deefa64277d796f4fca7bdbd9636b286a71eea1556e9ec4453;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha25639d1b11788a62c2e308bb2237c97075edcace2e700b3957cfdf2f301bdbb428e852af2f008f88592c66cba1375e4939cb9173080d09bf91641a3ac321686d1fb22a71845db631a51a745245ed92c6649a0574f688880b72e81dcbb406491a3fe7ef8ce11976505;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10823ce142f860aee03600296a3987b076fb7dd37eca1dca29215a2c429c21a94025347ab1a79f2a97b98f2d8a25fa42c85f3451f54258145113b37f7b966f31a56070214b83029f9b614a3b42ed33945212400f519bb4b7dabd099fa45c05b35cef55e0978bbc68ae1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7ddc1962e583784fa59406d069da2822786ad8c324f8c2781efe07ef8e5555375d01ddafdc15da654b81861bacb389568103054bc4abb3a429a691e182d6ff51ede5a04ba644f15517dbc494a66f16bd566b17ee5f80af5d8f8b42370a0851cbf61db9d8dc0e14ece;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cadb601131b93e94b8c3e69dd8ce8630cc34d2625712e7553eeb5ef3107128e88694ac8af07d7a29d4552eaa0f4e06187817280eaac53ce774fd903ac07acd8e2206576b5abadf3ad8f0418fed5610b96c30977db254b7ec748e5b54242f114de50abfb9ae3aa3f3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34f1da33078580abc6fd279c11612be9e014e7dddada3296087ced4d58946ccb954ba55a461d2594e9d2f89f7b31bb215c1df6268abf183138fc11a5ac7c207d58332686cc29ca1a75de8c053fd7fa242e7fdde2751d95ce56b5a8e2b52df955a47efa5fbcdf12034d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2defaa34e9ddf1e75d6b511193c95fcd42e5ba4da73bf6d4d13cee18d51d26a7a6d8a8e1f348764abbb05a680dfab2791a202574af722e519113e3b425244f0a168d629f4cd5e318f5b4e840ab8c2903402ccb32ecfa0f5c36c3db30b6a6185b02c3ea99b5501b4167;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc333fa888af9416796130d8ae2084283df72f521c11ffd0b68f60d31bddaeda53b2d8544efca9da2f6c951e83d28e42fff353495a3c6e2e4cd75905fc4a9748e6145d831cc6059415444dcecd39465a8db37cd2dce7ae4d19d0d0960220239380700d436382f753b89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18282e3cc0783a6614bbf245d40153c708e48705397cf4feb90f5f3cb220d43ab9b2c5b56f82af9368381b18b156886883c666f36bee8c6fd181c8d21bd54fca816376695d4cdd4ff6f1a20c9ca253e99a2e25bec19c52b1741c76955dfcaabb3aa1e3fa425b2ad0954;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d849ea4482b973f3cbd9b7aab67d26174a58b03af1e816c9be32a802ecfae6deef62857b869262c9e99c5ac9774bf1299bcffafd6ea49bd9f13ef85b0dfdd9f83fc9bda90cceef45610004eaf86bf2f0974e1c5f8fcc9ad2a141c5b8dc21032c6485a48b14f741d805;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92a677df63329923d4f51167abd8f0a34e273802740d08cdcf000ee1ff7f77fc848870bc7bb73f2cf77b41067297064008db4911bca7358154cb3228ac77140b0189c2809b89fc79bb29b22c44736119b4d0765963de81e7a2f0c5f46139e6514908c4714ad7f47b7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85ace4b233dbc55b87326c79b8e2a00903bef9daef5e5ce291e13abcece1cd3c490ced94d48828edc150f955c0eaf6ab7632161624901de642404ed6112394194da13a4d52cd30568ab71ec3b64a009e76f79f56e4ff5aa1f9972ac6b152a45f9b0ade74e2a8be1009;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10710b026b15353687a3d51d2c50457c2f9021b7721801f6ce7c5e507f40868cc365a4db03c327920f33015e2b0aedcb2e1a74ba4fc02d35505442a4d615d45734541627649bf4b6156707252613151f5b55f4cba77344f5f4af3c0007a6a8b97afd6804d609ea5f74f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e61befc5072613a7364c20a1a086c6a3a729cc6d528540ac61924c2a12635a23a8055855ce837319048211b3cfbbff307b86c44eb357a31846a9b41a5d62b0a60252f858350173ee9b0fc7f967909a9a3f641a754c73b6168069eb839d3fbea089a02f527c4281e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb29b9181d668fb3b613a93241f5361f2169c6b0a1a46cb542f684f57be9b64bc0aacd62775dee0364226b1e30545cc1ddcfcda62b43f7a6369d1d16bf1f2cad2428359cf9f0ae59db763b8f557664038f9b003a027ff95a85749fd7e4a094b28f41d7f2a3bc93d304;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h850a5afd8725e0c2ee911af05b57df53a57ffacc9348c916d24395c404afb237875d489db86438e58f7495c8ec3f035de8685d31d450459e1f7bf106c20b7caa1a3b4e58ec2141886f0dab1786ef701208fca7ec9f976cad03ff5469ba7df0b4b7075e46c97c022442;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c6301e12063a9f46550da91b664c8dd81cae394d99982fe6c2678a7a502c805027423db2090cda02a4bf95dc062c456bc2c7529a7265d64e9c68d8e5a0876d05875373ca8c4e99f3c0dde4f35483b9611767d6dcbfba09ae3a5b883e6b2f7985662b9b82c13f8ebe1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f95322f4597ccf8b30b81bcd8b22de2a2862a303441a24c410da1c1d6e4df85646072c5e14fb7851a6090f03fff14ff50fc672c7827b76887e434b44f94620abc8fa649c645e43fbd2fd8b7332a24a0034faabe3fe0dbf8f229694830334d72a68d4f4e25dd0ea25d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3de7878dc35fd9d21416634936fd968d2db8076e2ffdd09aee64d177a141f0741ba9dee0d023d63c3edb573d964d0051ebc865c21e293f739077c5cc013a32dec3ce9661289bc5ea17eee35b118c2ed62b700915f0abc24245e845cc3f5fa535d6cee7d43c5a655da9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1858f46aa5b987e9eed938b06567a8737ab4929e39a4cbe1b55db24c010c4ecfd2d7fa01470461662cccedd9504235e64663f0d41dbff324e8a26b0614ee3682d63d6c4f65d95560c4536f214cbad8e3d086b5d94340fb802878273cd919d0a830167db5fae1b33f86c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94d0a85b0d58ea7b03113043161acddd5cf8f09e0e6965720b43a98140c391ac3c51d296a69156cf13e3d10b2cd7e62835841c8d8b030f4083c8ee862ea3131529ad18a6df24b4421e5b17fefea16dd213be08b986a973e3b72e0c2f4c43a00b3a296386af466a5158;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ceb56a06ffcb3f75ae099c38a6ba39dcf0a1bfde085f42823e30df13c89e7ca0223212d91bfc3fb05c32d805ab35224deecbb439bb950f03c6a292d87e5176f08dfb08253b56817211293c94bb81c4c1f87f71ceba2bbfcb78038a7dbee0726b5a3de22d40c2f368;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ccf3760aa9f52936b83d443cdd492f986b446bcd171d37087244431368b396dc6b5e15f5cc446e38dd07212817141ccd9614e5b297006941daed6572cd0c04e467aed8416195e301b2306bd19eec6ea439fd30d21d932a01b4a5bcaa80549dc8984c99876e8e8c27eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ada0a329ea4b1f03639a9818d32c4af2b81a5ad08c573a2f8740ae582c26c8c1a3a3684385cf366c7a85d0a985d361ecacbd3e1de598ed024eaa1109c6c93eff724a41d7bd5a8592b8702b9753db8e69c5aebc915ede3a62002d0ab21b1dd2606de3c63ff58229588e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11402b2e34d1c9fbf2b94ade38ec7d1eb0cf9cea05f8e2ed4a27e02645448bd6eb2d6c54530750f101fe05be26e1dfe4ff66d9317a419ae01ccda0b88ec676af9b3e520d8b4a9027306519a54f0a1076392823c40dee9b05171bd8f30223664fc3f27ac9dcd8347b8be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a03858b952f8b60a5728f3b86fc4431b7531577ef7e917d9ca3f444b3c2caf992f0fe7d6e2d709baedca3d7473634e0fcd3f7702faf24bd226685f4d9d2510ad0f066093e332919c66f56b0a5e30a74318a6a06b5252954fb39e1cad45c6c0d8795f352430ed653064;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10cf09095fadb34cdce7b6bb894598c860979ae6feb14f4ff9892619905a68c068e4ae56ee78a622a7a87f12b227f7fed28ac4d5a2dad724ddad679f42dcb2ee823748d4f34c7fdac663d3475577922ab6b4c48240be330789598506f89664a0945490fd4995114332b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e0b42d9cc118100961144b7d7ed9c2a2cd366845db94abe3858d00f59adb8443773caf4f4745a27a2a04afde3e42338a5f241fc8383e62d2132d7b7e9ce1faed4c472ed73e06a23358c6a238e38fa29e91058f2e4162a5a167388900edbacdda366349e55c9b837fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f8cea4b8eb85c12604eeabd09720909484fc3b57e4b14b6ae3c3911bf1bfee43d53e56fd63564adb52497a7e6004b77312e549494df9e18f4573c4ac784c21ad861499d8cb68f210c37a49a5ebbe651244a259e52909cd62ba3efe0692be1ee0d957a0022d718582a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118819c1347eb32cd01deca65f78b2f7686acf4aa0459aaa97c06744d474134a60075767b1fce4dbffe46a66ecde7227a689a7b67d8dd7801d9e308d5b8813f6505823932162177c985e337fd982c9f365523258b68f29a3c2d83465d3a4300bc3d745804efdb002128;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1168bc58f0b4a7daa69ca5b11767586cbec1114409f5364d9d8ed0bd44653f211818de4c2e58ce492f6bb60ab28d966b4b13398397f166cfc7d5cd6273dc7f38bf8878e48add8fa25d5c7d1c0dc6a9ee5cea49680d3b2e9eea147ed5b2623fbab0a19d2093f5f509d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1344930a1b425f7af5da53c20faef18fad58afe0a2face78ab675c1d5bdc82be853feab118b491e4546e8bb5cab6fa33ec2d81359c7f31cd9daeed488e7bdeb0c9db21340342b3f15ae8ff15469eebd8c650daf942e671a01e2a7cb61bda9e931ce1f43447488df962c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118682807328c8bc1d20c7eb096b1db6d5896baacb9db482dafc5b2d8b5a9f57cb448937782b3f3597e2d08f0282d4f28f3dea1d7aa578e7f94bfab6148d087e9a7735b8933eee343202c012e14ab8ed119ffcc0f227ef4f8671d81c8daa5f8cf4424ac6f1236da2f01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183d9f461fcf0dc79040526f1f9dbe114f4d3d902e78bff482bfea77870472da4332b097c7b07570bf096ff61ffabea6aab2af2539d609e63113326cda92fd3469036ab198971dcd8c577d0c7449cd44050851c2029a3dc21584ded376ea8b0fdb77422aa3afcfd63b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab6eb882643923ae86721f52f3d732e7f2031c8a192f67eeeca905617cde1772cfe9e4baaa17ee3d13ffc1a00a20d165e95746f996ec63888a4df9b83e46d6934838137baf0b74d94779ab6f8808f1e01de13a577c250686f4bfb169bd2f5dc7efa5ebc2136d3fb7fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6cf31b05d989eeff50d7edf8a0632de571179aaea5323385a4ebf3d43a61ae88a9905f3d77848850b38574ce48b0a0b4e248ff14d084a31762459ea557e1a0d9aff62c18b98b23baeac42efbe11e3c93e7079533f6bcd24fa31936150aba856017a7efbd867dec4b96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18dcc429eb853ef5254ce48752f24998e1e2b7492a7a85f1110a6d2404d4020eb2b1f3c430ed5946bf18b0baebc43ac05d79eab2a4ce678ad0d6fcba2e8dcbb2b319f745516f2dbeae7d9468118f65b5554320645e6ab84b0d80d36a631d395c714c951a26cffb37268;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd261941966100f585101abdaec624a05bc62cd5a7f3976aecf5b789dcdb53d84166d70cf853ff376852f49b4963c73e27fd0a798f75669383b2ccfaa11c61a8d29dbfd4ccada23744c558efdf9f1a4ad49622905d002d59d370def636e4bf09c16bc89ac992f81b3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h674d4eab18e79c050ea1a39e3462639f0f757c5b7bd29bb0e9560032825f584dd487837e03e038f4214aefcedee0f8951cc26b8e8e08298fc9737703a0c2e4f71e30324b5d1f662110e01db06bd2387a436cd979f17cca2fa9ceff8670d5bc4273717b0b2d11096b20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1305ed41a529481fd7ce11f91144694c5e2c27911f0ce7e00b0fbb9a328705294a23b287ef91e951079df921f9dd64e2935d0d5d46b1c3be5a641d1867753ef70e48c55bbf0f529c4b8dd23914f290a0ae929e25c579d0a1bff2b3900faef21c12abdd522bdce0e48a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22f1b74df87a7161ae4557e3bc96d79bac822a4beeac35b77d7e9a1b3b5cbf8843f0d9b88522000985ff17513345a078edc46eadfac927addd4a294bb9483fda1acb976f5afb79f0990a927e2b095def2944368b997fc657d6803eb093a4c04801cc430b1f083e0db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9327fa7873a805ff347c67ea06772f5a7fc44eb032fda9b1d6135ef93eef5784e56b44685ec6b892c408e6f176baeffd8515ee9f1dc2008c9925e7eff14332d4b4279d1623fa3f30100787732933e855a5363cc6bd8f531f6ee185b8c66ffc0a477f967cb7a31627;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17129cb1fbe89b8ee0f21ed14960485acac345d1b7354329a6b59eb45e25963e99480ca3e3741c7107e7668c9962d387e3d32243ef2a83a12a590838f3b49de620ac1a730515a076d1d7c79d5ee69426726d371e1284fea39b72596f41e5180dc7c6a62901a45927c33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c4dba44273a6ae3c7500705866ddcd6e8cb00c933dea3d5d95c84b3da2ce682e022d8ca3bf66dae4284d7f8c3a7b9243eaf2961a1a241467e17c7875efe35fe2bb2273bbe3d7e44d531511b1cbace2da6c6cfe2b333b5f6927a971ac67263ebb30212a633804bf022;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c413a630c0b7388496e32a338b2e2b83d24a4f0015932d5e63b428e027ba8e483574b90a2f8473ff233e3e11d98ee1d69e04ccd323f0577d0d0b978796ce809ed218293c5bb9c0c2782c13e54416261fe8d7befcfbd195e08661f2a90e6af7ae778468ba7a4288ced;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d155ee5d23c0c27bbe156b0dd4b4b95952003fd8630a6a2d4bbff2bd6b75a8c63724430589be9613b2acb15fed54c8a17139c7c99431a422f5f310b67b07634e8af20a3287b89186fdb06573508a38574846cf81f69f1f89fb3a5ec69d99b1a8b52278a327f9b0e0c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0ee7a9d64ade00e22ba0ec1f1cf1871c15dca98b8ce50f32b04dc4bb9bb6d47e8c7d38c82f33eb83d97dd1ed51c2be507506eacd3a81d4a8df2c19e6380dfeb29f8e4e58dd866e5a3a33aa889a5b1431f4c5cbf355d13b36ae8a54f42a06bcf61a0cddcf52ec0c82a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3eabcec7630b75dc5533a0f52e315c41be5882464cada1b08d19c1c3b99b7a7689a43a3507e421559a827bc01235fdb1844ee4c80f438bbe4cbcf407867ba047ce7e0b67934c882ca9acaa190247356b76c516e9bee9fe1e4596f7faf1305fbf655b571c229cda62f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h249fec81f57f6fcd13eb44cd3674354ca1618c6c51f1746f438ad13e815f8b0566dc9bf21afda778afd0da79317d179064d381002049698254122ef828abb0265ccad4994a9770a79c8664aeb9bd7979b42918c53ade6cf3174777c4dbf5cd90b2847ee39db784195b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76cfff8cf8e47f34f34e73ca7c6c29a290e483a8bae657f0b71074a838d5299500a25a943e375d450404777d1d726747f44b8c6cfa889edbbd75ab2b347ccbc9cf73b6c46e387bec6aa7059ad9829a2b842c756c44da61bdaa78cbc06c188b045daabc1160cf656b8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd83a7bf9d6d4e7a901b740109ffa516869b40c44c5623bed027f215ae09c9283c7ed9fb5e113c900243d153397f5548bfee631e7f6276947e32ba5cbe1c7575c2b40cf666ddfb63d18dfd7e76e2fab7a90653e8cf417cd0dfbbe938d87db085d4554c8bf1e3d085bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db7c5b30924c12449f5377e7333598c8ebb4b2a4c059449c791478a7be9fd6b120111c52a35e0c7f35934f851e6b00d494c85500f0d848baa1850be28279f3ca062f458b6104cda7690d4f995d7a42a839505ed296f2cc3a7820a9014b3855ee29dae0b89fca6b5e95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f22fd4e9d903033c3312868349744c14355b657607329a7992f923cebadc9ecb77b4a0c0a47fa2c6a15ba5c173aa380108678918162b2863477d51a5ddf2becfdd0a52b91d95905c4e8c4cb7e56470f8f282ebb443c94ba4e487f072235516627f92d7fe1189323fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h221b993bf7e152e1e318c1a0b90e637a5d2fdb6098051c6724dfe9b5ed64b98ce8092dddd5278c43b4366b53512989a88889e50b97340057eecf2f718fff884b1f9d17de37196c539d8f8094e7198aacd9b2c5b709e554edb60860168ef7f109f551fd6da11865cf72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e985a6f7c54b38cbf91837f9c62a1cde977a72ecd4ea8afe40b503b77afd6e80159d71c35291e4aaa215ad127d5c8082854a2b53f7576bf256a0a220da009db5d7084ddc1ca666d7af8dc64ab903a4994319172995f3ed9ff4eb3e8ecc4296a52b82b09791e1b34b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6afca691d99e26952858f2575f2a8d1a0715f26eafd55a23dc9239d39673fc510489eec9c697f0e2333d26f3df40db931d831a49fda4c4e61642c78eb0e8195f9b19a08d460b84dc83e9339733d4f82b248a3fbc5f6a951ff015576c167bf28d640f34e38fb5a5e194;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b8fe5c45954f39384ea6dc69df599410a27935f37a2cc09aa163e0794c9891d1666e560f588a6f9494b4e86524077e3201d537e7fa216b3546fdc15ce91e971cb0134d19ce607443c6c043c380ba67f04f57579a7c4367d8fac0d2a948faff667328766e3a395a77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21655777630d5acf20122ced962976f374bb9309471090fcc9f50fdf21a9c6bdf6cd06bcab2b8c9a89dbcbbbfe26aee066c658601d99767ac1abb541169700d50d788a715c1edbb7c7595d85853e5b0376eaa7a4e93d57b71f557453cfdba75842325bbaaba25a15c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5d4dbdf3be5616877139f66e6e2d938fe9336c304b2ca11bb0ea40e840aa7f9a9c069778e15337cb98075fcfa78159e7eb56f41bd8191c38ce7a32c418cc739c97d3e9fd2889508214441c4f38c657d55be33b562b05d2d6be467a948e32ebbfe31ae0ee4e2e5708;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba6b91890d5401a21dd446481793dab1765269637172d8793d05e726928b7bc0edf6146d681507c3cc66cc569811d1e9dfbe200e447417f2e302a9596a89935c69e80e2560c911426f28601571e7a8a5023e682e4f881f75359fe68c51e211acee958c9d967230b0ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbab6dd3ed4da22751ca37f0bdde4225770ab2f3197fc3c19c93a5544f461faa6cb3ac6fe710d5244818fcfb91b9038c6292df8967ceda1b10f748b953e340eb20ec996c1f01425f8e092a10f284de9cb411c400f1ba2efc2e7a998fd1b130e472508997a29f7eca43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdddbf1dd1937d7af2109d4571877c22fe7ff4f8e29ca5dcd32ea3d560ddeb08ff7c643e48eddd6c4cb791c790f0884c5defc72c048cb17b8cee757f2a8dc9a400263bcb9eeb5c24ae32fd1e7039de5a62f34132f19d717effd18661df081d55fbcfbe5423fc3fefe15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h754403a03dc62ce646cd5196a6876d0b3874f303bbf48675689401d274d6933e89ce44338af29a1a6c41ddd0965837a5d84e5a136cb6ca7a1544d2fb81062d85a738dd51591a3f37cf116ecf141a4355fc2b2781d218504bc8457b8d2f1a12a6391326787f8548127b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27d0114f7076e161a22ef3cbeaf30aa5b5cb9974b80711664701146607f88b2bf397bfa6a2bf4a8bbde319b456c1467bf2e7066ccabad6aa7f59b853456f18bef680bf8871bee21faabb0661e224178b8c59e13934d4245b55838d7cc3e0192226d87e1615af5f43d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaf2d95ed5447de043fd9072e105116beeeb03b3ec5f8c0de2668aab506c5f95a3903d94739563ad23fa811bded153d6f8aa6ba02d40bdc3f4712d2e82d72dfa66ac1572122ed2c199770513a0b6a441a0128282765613cd38bcb4d16912f909b97d0c1d9f247bf13f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c10a68d0923d2929d8024f7d4a9d4880786121ecf47b7863f074b89f7db3364a59fb43c8bd730c7d6972c952d0074852ba318292ab8f73f84544f24890b988b704d7726d0e2abb54aceb588954b12223e9296be0550f9efcaf7a4e065b7523873f28b1cf5b7b23e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f5917cd0a5f4de8b73499c2aed2c13263a557ec50f2edcca7f82ee909ba67086d848d41069d44f840c86d10feff6b4f790b870435291a686b70714edebc6b0abdd7acb4e8084884c6177dfbe0f7546d5ca7eb3b38c834c21461f00e4669b66d8275a34ae652796379;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13918f4ef5c2a0d7e1f5816498bcd471c459ac9d441a52a83aa71c645bc2b304571b7b29b1392ccd8ebb3d81db6e3b9dea2756f13b42d2c0fb5cb35735fbe4f337b906d3e597e16c3c512d85a2ce3ad30ab200507aea8eb4fbf06eb966f3bc92ba883f5a86ef34351f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d4e0d372559b8b03cdc65e21c140c6d2924f79e8559d18e07efeef3379005882bff8160acb506436384fadb85aea5a096c251851dac7f71641cfc35565357b8543a5c1b389ebf828e858417866f2673a22f557f59cc91dc40275353a42169f05c27ee24ca7fc9784a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcfe562ca3aa9e56153e39c302d43e9924c78523808e1a8be37738be9baaca375fcedead0f518d1700d3ed06a44df3f178c58c227433595669f547e524816192df893e3e2e55ae901996b9dd0d83a435b42364f4c041fa70ab6018c907f20e6a3cafc66893bbaba9025;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a4f3e47c53193b0314083ff052d5910ee67b562d40b2c2a4b780217eb7ea5ae153b59f4be1a3f1baf83f828efb3ae04e5ff138bfaf7a825b16ea73d9e39d352ae45b42a219a2a576d0405669a00f4a35cd3a9f604097b5086ff223c6788b88e1bdadcd9ef2b173825;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f7714aa496ace95141d422881db41a745fd95f19bdc059fab99d2acc98a0e926a5569f6fd235094fe675d2e46636dbff4953b0eceb93ceb93fc872d67c3b6f76c93b7dec2fbf3452e1d84eeff3b46b3efa69ffececc1ba4ce942235f9b5168f3a7a8282ec2550026c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6da46b87f3b64de61c55441e876d838dd2b4363b6b2ff6729ac42c826ed5a930a5ca3c940f36ea52d8bbc15b36622265313e4854019e7efecc72c6ea65d14e5fd32a927f031e0ed1db943c398484774d04ef1b68b849d6ded5cedb4b072c0fcc3662130577ba85e83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1becb52876ed65307b07657bd161000f3008533ab653b437c7f865d879106f64b786d3b70aa08123394736553f6669a6bb61b526e395729efcb933aac615e1941ad5417a077ad0148430af402ca8554360d9324eda721df2a4719a87847cfd86b9dbe57d44815bf1605;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h381871d863cadc34df9302ca9805e9ffd353b4b55d01be1cdbed20546a03b8161ceb7cc3c881c90a46646a951f1916248d3ba6e3ed4e8af878b9716aa1fcf7a142a0717c6bec28819de917a3bbff48bdfcd7840700917bdc9749d792e12181264d4651304b02aceae1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e28f9aa3619f2c7505c30fd638de03ca7b42d6c327d0b1c2515b11d49256b863e58b65f86c427cf103aab4dff89cd3594d53807244eb80a4d69e746ac335096c0aad75c1774e9b7622f2f855753d903c47801f7cf0889f796deaeaecdb3baedd374dcbbadfcacd734;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1665262ec8a29bcc2f5a2b9f8bf05109d84cb2d3eabca53b253b9630b782ffbd05696a8aeda0260ec6e52190c86cb95d2b4bd65d902e68d1e4a87e41cbe4c9b70c55dbc0235f520fc9b7c0c4ca7d33d74f6039a7f8bf332ad2bfb3ef562ff9d10ddc132634a95a34a51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha060f4d3fa18d3bbd2c6f2653b46b245fb03ca63c624ca85741a18615353f2c838e60758bf2cfce49813e33e75fda5064ac7c28c313b6debece454dcc867d111c89af645c17ddc277ac9251896dc2809538411afc6844f7bc1c9586e567ba9fc422874a71ad9bc8060;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100a2c367d61e37df4fee39da9e4d45c605215c014b7f2968faab374f7fbf422b4ca8bf8d119f2170ae2cc08dc31ba796a24953e61c6b0e26946a46b6a22120f5de8946446999a37c73d5957aab2f8c16cf8cb01a4ae76fb10bbdcec524b4e97f28452830d5552de6ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf616f5827e99c17dc7e2ca425cfec03d7feb31fd49993bee4090fdd71579db5c7ab0fb0232265e47d4ebcc939e292760c20421c12a88adcc83b424df170215762b2037d1e4d9d9cd53880775b8c340477c0a9f71c3d5944be68a87528d626a391251fd1cf71a539185;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd4a0390618285248b80abce1a12067d706eae2b32f6e20c4c8acea4e7b8ca8c0ce4ed6743c1b18237295580ac3853c26333041048a414f887e8f8c3e898b26d1bf8e0fd0fb51e0f599e9c93081446fa7c93f463c45e403d4321cf226883b16028214d87cb0d06cc991;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde4075be0b25412d81c52a265344e3410f0fcb1db75284be2cb934a921725c251fc046edc1a17fb514006e0f4b4942334b87f41fc7af301bf785d7d3ed0489aa118d645dd55cb19769c1cec1429dbb1e7a234a0208ab3c3acc960dfd2f33117cb3d78c6bf47fde0b83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1aa114836dac9ce348f8bb0f35756716b30d2dd45fbcc3939f79590a28663816451b93ee1768337c01e0077a335ef463bf332151341fcd36c1bd4c1bf41c2af3f45c9ebd34dedd7146b32519baaf4cd86d31a899e179478a1ae95a1146b3b1eba139e8eaed6a700e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f532a0df4bbe6983111c8be18a5f1647232d46bed99ac900bef5d10a35905f2d4c8d9134890577826c5648688237c22500c563fbe9c5633347c51516639ea028868171fad43e97a15cd58a2758e7b80314d37743d1c02305f8d36dd961755c880f01bbc5139bb3e3ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bc334d7e63e756d72f73d48d19c8b2f4a4f6d09ffec058957d99cf5fb823ece4ee3bcc0930626ac79b36a183d6a9e8a99a7837351cac9cb21d7e1dc16834966b5c041e47e16c5286f39cfcbc637ec99d1519897af24378dfa6b1dfd8b239087d5e16efff692bd0631;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35813e049c75cc18c92b1bd7a9bf10b8826651b56d56ac5f054f875f5687e47949bddd0d7d4e932476702e213e60bb1dc250d8fc9f51571cde32399ec3e17b43baf8162de82c6bc353c6c23ac0559b8228fc35a0cc7d1101b84656dc7a2cbf39fed49136dc8377aed7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63be35ec72da154e0db2974dcd9fe3f6a9f353465351511e432968bd45fb6027c8d628679ba0af2213a41ff0ba60d7dcb3802a1c04c6477d9722a6831ac7361232046a3b4a3c379fff040e21304fabca314fc6f1bde2bfcc402b623bcc42346cb9076dfe1e6b0ab1d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a321b7f59584348e7caa1414300c0b9cc5a63829efa45a09703a6c24d8205b45f529c132752647cedffee87273eba98c41d8f6db4c4d31d7c0f538719d42e00432e3335b8803ef010f2e5ff45dfc3612b6b410a2765eba30964418648116cd8630b39c6d9d53e0ac3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e9a3045c77d05c6f11ffefc6b00be16011ec8c49a579e66ed7cf5a33c4f178b5bfe5d48b8adf3dd4b76d8ebcd5bb3242a284e3aebc03d41f7c3827ac9744ed42ad0dfd014250930d775eb34cccf593c7846aa5d4495d0a1c17c7812c01fead18297677cf50c8daed3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf597ac4d6275677fbf8bd351d3292001e2fe4dd5e14405e6bc5b535a14fb1eb68ac76ac0fec1e3211edb551dbb4ef3cd69a834d45711a02df012c10d6d84c1b141ccf3e883e4dd652e78d7f750889de7011c4f0abc4cf69a748ce354514afabc6b7f3e7fca0599036;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b4b57fc08df5f0e3dc5cdb5fb9dab3de9aa2429eb0da8a49bfe54caacb035578125ddaedef8683d9c254a908057b6cdc1b3e08ce4b4cc6a45ca7c59871c39653172a4f45ebeb362834a8ea20cff86cf92357d6f9caf60d41235fd9cbf5a68e99712e12bcb14524cae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40ea24dadcda08d949624979ed69e4ac0902b9365fcff2723c4c513b67fadb1ec4c2c7394b0091621429584887035613551dd601ea9cdcd9e07b32c604ff92bf79f3eaa28a90b5fa824f0cdf4bbc2bc1151e16e75b7ecda1705eae3a7efe2dbcc07b336e1266e9ccc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8790a4e825ed45c10b91d2fc5f4a040f0b9d7788ce183a6806ead7fe3f1bc611544c0380a85422adb755bb9f7b8aabb02fa5420dcff480ed125bfc02f803e363b13f7929e7b041598b15f381762696fcf9bbd594f3b40ebf18d57815f058352d5d7e92328bd08fcab4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba9bef060cee696392cac858d79e1be65723c303dc6c62f70e781a06107361208dae436b6f3efe24f32ee780a6ca684209a57df2b7d4879ac412a713998684434874dd6a53babcf8ac37dbf5b428cb7fe1cce84d8258f0862ef3c441c29fde9777e2bd28c520cd4ddd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5dd822f01fc89953cd070cac9e1579d6250b1b30d166ee28c25bfdfad31f9507e7c57f56b80bd6e4ce10638181576ddec4ea026cbb171f9c3b1cb4e7c081759d394a1b66db4182c2e79f272fed0a0352c3ec93ecdef74f676b9b2425ca647e465c4f7cde767623378;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30c2cc32331f18c201b217c70a3a031bba5750577692ffb4b74cb68af4b575eb6bc13a79c91a97ad1e060ee3519668685b0956e5601884a25789f7f86411a79e5d7badd77a4eefc81c686fedffa23e06b47518fdc1622fbd66eb38b4f3a4e7948d4418339d7812fc4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b955e1cd35648d446343ec65a5e8abb2f34dacbfbf361853b10f1b39d50d7518d925f99b4ca7c10d51fdbbfbfcf59d9c216f8ce25ce6885e4856b4ca90b85d03cd9cfc18c22127b20eb4b900f71308351aa2d96d9f8c62f23b3f3a11f5e74fdaa05c6bd539d3c8e0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca1d3713cd39cc256a8c5675aff629ebde00cf4642154903ba21b423988ad130973693b9cad95cff5b51b0930a4b84023f67cf2eb8ce60b6969865196b6c2b79d931ec47122337e84765683523407840fa03edf1418632a606830b910a93bcef0ea019ab7fa3613831;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a6edf5461f33b427ec348948adf3841240d67fca840d624f38338fdb3803925097f490b07f7c3a1f24401d1b3be23dc26191b967997224307ebac54067cbe9bb6b7c99d8d254c8e3b4fe3bd287f0d26ba989820ca310417e38c2c6abc2842633a426406345f9a7110;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42d7d1a67488fa9832e9423ec9e771683e9350c38c1d2e08e026ed14a87f688f044a771e52b2728169a195c6fc37ac937aacac58fd9339ee45948841e18b1bb2c234dc28271b7c17b86f09ee6a72c6be0f0dfd13b8a5ec5b80dca88e90f732f1558e2cf579a7c5b287;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8013baafb15e2112b7b4d9b66bd26066064f29d49842e786f96c28877f3247d3dc0a90d10646a976cfffeae0badcea90baa8830592173fba249d7158bcb9534089b62f6775ef8533320b19bb7180228991c46dbba8a9879772b69030c1d8cac7097c2be209f24c55a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbec65d1d7d5fde35114493a4da395605ecf4f68497e2934c9131925d033d9232d46fbbfc04916b7e0e6eaef46e611016703ae2d5384358391348786d43623f4e7f246c2f45c9b66de17c277beef0ed212b520de5edbda9fdf20726659042c479eb15cc01903651efcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7432a3765cae91a3b4b29fc730beb70694c9a35e13e802df691ceb0f0ff9748dd500f0b1fd9fc0b6527bad2e591471ce923e17a1aaccf5682ff99f4325b421732f4a2f75451473b676a27f4bff35e2e2c83eb9db89c5055f4d166df5242a877f2c098a550848721a07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h591c705418db84d48aa672ac0298a610c0eb546ca84d19a2a5705f2af9e7e7e51ab8bcec41219c2cc68943caaf675b7dc5204777b296a7e414166ca9bfefc54ddeb18aaf51e20f08c3783c791877fea88c10cd598555ba99aca2356671cf036e6518f111e253f72c0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1013de3f0a75669a0516af9d9e473c0657eaa517775918c3aa1a28d898ee51380b8ca9200ba39f3681b48e27e199587d3608cf8f3a23ac7cd108492cf9373123b300bd7437a172e2d61003ecff3d7a9a68e6c51b690e6b9fc9597a7d5f9587f134c6ad905870f3e4ed2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha232c1d7d4b1460031f39ec09a216df128aec6334f52e8bda81939d63caf969c69d422e395102a20273e2f408a5eab74e35fcc8847445dba532ad771d8bcea91b057815311fb467a74ea5e7e14c21db2e15ae2fa46a0daef0dc14f729b4cac8eecfc44a140014229ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ac899692bba60d41d78885212ac13183de187ba2ec861685ea943fa8c224edffc2894e2c7ce5d65a1683d04839d31855cf13d0301db5f68d5d14ca743b2961148db72858390f5cce61e9f2a0ef092cefba3110732e3b043d3216a52f149a363ae6de6bb75064656bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h574c107359a688cb71c60ab74253acb1ee4a8528cd4a9653f211848f9cf6ab235cfa1cba16af29e22cbd45f3330e2abb5961ee9194ba70e67fd55248b1510319e76357b55902e44f4f230c1aaaaeab8f640c6d97f18bcb63508a9f5f67e894eb5af5af15042dc1b428;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1b82ecc8bbffaa9554bcd7218a3ba9ff6c33e8d61fbdeb3e8464b2c6edc0bb8147397e53f55814f17fa28cb8bf0d2adf343907c8b9c9a5245cf2d0dc69b3ebd63ee7ccbd9dda1314cfb74ace4c7e30fc3692b0e0676d69d1ad8870bb67e64458762bbd843e53d1a40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c78cffbe676a0b1904ab2907544768a79d515b44d78f4ea3141bd5ea7060f9370dde4e3e9e280947c54678c17fbb3c65b6d1c30cf87d8fcac60f955005cf8ebe6b6c41dfa942f49774af25695c53773dad91854a84333c138599ab4d70553db855097c974015016ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b970dffc2b66378ae15bd4a62b4a6f74ea7578273feca91e632d475c83965edd639816c9cf1d0e1120da93c1b6b2fdb02c9acfa9ebe2ace9a942123070a8e123a0bf358a00c32728f4077410549e39aa4b51158fc2cc8f1ab6b44e7eca448879231d193fce71d755e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91bd8a6333460428605de10da86827d20e1b52ea9180ea6084787c06e63abf2a9449e0d9aa722b3a626a79c716e160fd88536cacc4327cea760425f7d01bbfc50e567862163b6f0182d62181a45707ffbd061988e78ca05b2cb87e1fbead7d9c0954ffafb558d1c10a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9f7aa85d361ba23f0590e55059303f27d1f70bbf2bdca3c4d48fd92bcf6c3b6706e7e31413fb3862c6df42ca81d929ecb8a36506f687479406c03fb33ca8867548752aaf696682eea50c7a3cb96ef7e410b7614f9e552c27754e3e1d0f1c106204dc82c538da7f60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd32acb98643d788f97dac2d2591191e9a014907c4d4a2009e066b1a1265ea2b061565424f7819f7e6737bd027d7a47c2f993d39101d5739bc223249ac3b4d92b8189a8d0ad7e6b90d750f4c651cf85b6357f83e45c00f15637bdb8a092d426784b825edb690f45e18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8caf8679affdf900298138df41732ddd1662c1eb0f2697663dfcd84dee3ff981c68721b394cafaf9ba8812ece00204458b8a2ba610907fbd7911e77c77f79a521b1f86bf23b985ba8bd1edfec23b890b6991def977c4d4387e8b1a69aa39abb020461d89bcbca9005;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80c53e5704b8677796d823efd9d2c3a7cb6edfbfb353dc7f9043879cca944af049521caba3c43e3f7bdf6c35a915a3b662ff8b892e4a8a5a89e12577cc7429cda71447f5e58d83ef2db361fd36a9ebe31c7639670280d98c3c5f9a6d8dc006139654fe9715c4b6ada4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c472da7c150b2b4bea592e7906e0e32a1ad26312dd412c328ce3ee48498bac4e3952b78bb0808143b411fdc1c5090ed1e98877abc881a40f499384431c19a47e90c1eb629e50a786cdcaf77c9a5914592dfe2835dd3f606c7df9efa2a28f4b8d2cc95429166023941;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61c7f27fe7c3e49c96cfe06c78582e1a76a1968e5eecdaff931c050d0678fcd280db8fb06e144837a3130c36434359fa567cbec4b919a24b9a5273a5214608706945d9a6e22b934292adee547e49a4349b700774e0f9dcf79568694c114f1f535dfb6899c51a2b92e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68245cbce6324a736f40ed0a3b61529e1a076dd44c52aeca14a3b1aed470d058539cfe00881830672ff8936d9e22388d905c4241a6988129576b07d3c59293a72132bb742ceec4deb126e80d3159a4bc9c24c28f1b256a87773b3987ec6787fc565f11aff3bed45d1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3ab90a609566ab6a1a3d493646f3575ddd91c79efb5bb2e1da31c53fbfbe728c05dd3c9380aff1751a002225a2c07a3590eeb80a1effa527938400273e77dae7bd9730e43adfc5d92160a81b32f95f692b269ef84868b9c3e2eee991ca30aa0d1eaef005a1a9801a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf680523f787eaa3d6281875d75937c90bd073b1151a1b03a4fb04448710c7e310f0b8304076ab0175480682f5f7b885dec8278b7f14ed09b675462ff909e9f04e1f1b1e525c7897d038afb96e6f8e17d0d2a3a70c764fb20e4eb243649b9eb46f2e08338743cb2e571;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e787559207057622d8b180596a93023a76e56751b823ef75f7d4fd0757811e7bd0d9bea7929278dcc3949d5603d44f4448bcc3e31fcb05fe3a4c42559bca9a3fa5bb11f262b6ee73c130fd9dad2ba65ac6700c2a730ebec9a4a8a59da885a942d1b103463de182a55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7aca1d3a4fa13130f376431a4eb817adbd59733e193b1b3fbe6bae88f7819fa4084a01836cf640dc838781bd964fbfb828ded1de9fb0f9542ad2cae27ed65582f16e4e83c9db0f148e86055269d73b72d9ea4012971e983435a3bf495d9d1388a5bfab28b13857e705;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59d2989459d0501f61cb23bd04127baaef7e65b0b0009ce94f7e845a0e0f0c0b0288be2564f1d8aa0be54a7ea121e71dea808bc0a112a41df4c8e9ece0c3cd8ca12d025fa2ccae82f18177634020d544cbcddae4172d3f03d31ffe2dd84a3697f179f5e85be7d00efd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172cf9d5ec24ac6b9e98988269c00b60e77d6c4782cde5ce3d3c0ad1a5397fe286435217c4fff3a8d3788fccc2675301770704a37bec599b550fca4afb689e4fb0d3b6245ee7f1fff8b7a3c36a2e46c337d37df421416aff542f9e623715892e0621f55caa4470fe2b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdef23e88a654a3f3ee73b727b6b8bd19db17dfa01445df2305939512e9eb63b625fc927346b37d004b9883ee8fc19add74927763c3d2a50f16fb457eaa43a6d640b73be1fd874ada3d51cf1886e327322073b752a3d76ee67b4c6ce02604a9ec7084ce3094c35b34f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff6c16e282a215ec14953908f5c1c0a9f7f81955443abe8b8cb721a322d192a8437f0f522a450ebb3031d7632522b9ee044e35bc2f7ab8e805f9d43002d34218c27b5d3b737dcc104b27a897fbd96e8fd095a13464360ba2570c44ee4f4d3ab2f93a9fae07414ec62e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3762c1099592769b18ce681a71d583033c8935c4776aad54bdf93267df104e7eafa62d3e30a1f880405b2c9b1711471a77f57d102290274e193b3154f8d5a8dd2e8b380c31c15b61bcac202c9861b834890b36fd0669f22cc8ca88a3d88eb028962bb4f211089755d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1861bd61f5eaae9ee0f8669d7c55351b18dc54015585386ee14a79eb6b3095a1e509e97c95fe1af6547a159b7e04e0e8fd57f3938d344b81a029e2bb9a606a784eaa12043b84bf915984c3c6cec7f483f926a3ed8d06833ad17b0f1169ff8539a221c9a89e6a5559182;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7513db365bc7436455717ef1eb11f1dcb6753d48c8fb54dcd3e4d077ba01abb4821d4ce1888c0f9366b0a6d83860f4feb0e57ef49c0641ead534cd8e471c4c99508da2a2a1e610023b919a3f6c04895d789ac40d4362dfa65589876bf624fafa354bbe4608e32cc0c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101252c00e82103324b80c555f67572a3a5478c7f0da537813eda986806fd885de803cf8c924c4348b5cbb8f38da59a7a9aba7ff3779464d097894ff0d9db0e4549c69d1fece05761f790a86244b9510cccfe700d8620a83212d3de4bc6ac57536fb49a7acd5865039a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15588f05656ac448387e0ae095e9d253eda1b540d8643d40d46b84f612be14cfb5de6435fbaff81617914169b2300aedc3fb106e74af614c8d89e703a6556983b3a51d9aa43c876bdafadae9d1664b0e57247c1b4179f951b6d30033705e8389151e3d8beaf78ed845f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6385b10ad050a0258a074db251b75611e9823348cbf8f3575264d28e3d5b6d48e8a7003aea298e29dd930eceb6984edece6bae1237cff94c1d32179d046036e8da832e3b3d2c24c374d797de6133aa733a077aa3f425ae4e78990904e55f5c44ce68b6f747b4b1e2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8007528f837ddd0bd51cf130261c066b2b14ddb178edff6be92898f74719d3be8e7ca0d7000b57e7675ce8f8030e5362874534cc34e978af035e2d137d55bbbce5ebdfa61a4f995f862fb03f1f515b9f645eeba3538fbd5eed837d7610cbe69deea494647a7302d90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2bbc2f524791d27b3fee0870a78d168af441de744af8aa83fd351c97ed6d70e601b4dbc6e32ecca282ead0c2100c1f6991d167ad82086dfe2b9172ede9fd9a03a5a1c784f7948b82aa03563a3f24cb523d2c809d8ee90dd92f740d03ca149611050b5149c25d0ffb0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce19a46c9b951ad07c488b8de2119be0628fab666172ea63e61c662e878877e21ed27e62b188419cb71508c94b504656faa89d8fdc945869e69c1b7ada2a702ade4712dca99299501b88884415325a13212a3f8dfbac899cef11847d1bb5783410c00b6529b27fc35e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4da24c8543f1011b886f0b61250fa05dec1820e887f153e0b39d9d01cc36bd59122ce4675708bd10692c74509b1258bcb47d59d1052962e0c2aa63fc63543f85dd9c10f1bc0bc18f371ebb27b138df19bbd330906332dd7425ed30a968e048c5f4ce48918795d0bbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18768e0c944a7af4b8f5a2fd0a6785e92a85698013823833e107bf549c34ded6e370518bd2be24a749ca18ad0d43495e91fbd58d95a490205812f43c5551034a568212d0a065edcb3f7ddbdb4628bbfadee5af1e0448f69b43ba807140a51660db64283c18ad3d72b90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bc3e4d7cb4bb41418d4d70bcfe007f3eab0021c6d6dccb55ae54a0575517a492f75f6775b717d4416514aae60a0983c0d85bcde6a92aa66c5267a984487801ad5b00cb5861e156b7a964f36d944d83f3732c70895dd0a974e7cdc57270f70cc3ac45856d94985cb27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e908b2525ffbace9a67bb00b2ed2a1b8ce7fba8a2ffee0dcf3fea5e8e6beae720cba867acee87333427ec778608dd2f7432876dd6b34f8d369b0dbc0ca1ff0a8e722d133f8820c59fbf6f7704dc6a097c5634c3ca49baf70247fdffedb555d2aa677c60cc5cc8b7259;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h404c13a1f0a00e68ede78db602bcf4cb6ab4552c7dd53fff710a4d83a07d1af99a604eb1de2b0e9cee445af9745070496d1732a80c97e9d819498ce99c4a1dfe6e73e71586edd3c8acca4d2a2b6633714f392fa7e318fa15102db2a0a36fc699eddd328785bb8b4497;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3901fa803f2093f95d167bfe489d8cad9ad8fc4c2d674f7731c14b845f15b68bebd3e47eaf94837c4849fb56d2d44ebf406510b859037160e83c986cb90f2bef3cbbd2504bf4c5fc740b4142e163479bf796eb44eee6f31bc17064ffc9301bf4cbf98a834343cf93f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1728ab637299a81902112c9b26d0db074e9130ead8169fbe6b68f1af159e31fb149faaf87639029a1f4c6cae4c7a62a14bde63b03d1982316fdd278b15999171ba7459d395b6476c73f85d120ba339e31d2b63c60810b2db5969fbc6e1a4f5c1ef84ec02a902dad1f04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18afb2dd309935994569a8a7f614a08ab6431ac0b1e1fa7fbd8efbda6eb0f2465341244ff88555802bdb19b3a0d1c0a766a4ad0c2146e41991774c75057c41c3518244fea57671c706c008e4b9b825912b448287b092a83c984967d85bc1cfb8eab74c37c6c34189d00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fa9dd2a07c4040d783408420a0af10c4eca4fb1ad06be3e75fca7c66dc79e7c390560ccb027b5997ea73e9ba7fc3118073218a0cfa21a7192ba6526ffe292b5ff4e1eef661e1e4bd79ac9b58b5975b472b9fd7e82dce979dc8972e8cdcb026962707f2f1250b175fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6223e1665866bd2ef8b66fccc45c088bac085d0d45e91090f79c4a464b4a03ce4611bb0fe75aef8a26f8d39f64a6753c9dbcc620423a1163890ddf0f258405f49e3ac7e8f906a8795542abebcee3a0f347ca0f3aee30df4d43b3c1867c48eb7f7c4f55362e183b26b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151c674089130721ef6c77f63095e6b5c9f2d520ec651a73f83068806cb0664d2bd1a85b3ba152d1bb701a995ab46ed5249771a5ab6d067666aa2a044379b2c40d7e7f29485064b0fac8446189891cb50dbe2d21ae54bf4c768fc85ab6217a8eb6e3d1cf80d1720d4cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179e42d48eee2a9cf247641323ba77d727a94cb7d05e995ccfe0b8c7c6bd21ed8d8e56a8474f8dce3f28e500ce453bcaf02367a292bdf70d5140f0a3527073e8c2a944f1cbf8e7764b375e85aad3d6c052183188e6f306d41f37e26f226fd926ffbcd2fef1cda7a47c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9478d6ba85d2cb115408a0349b4ba4e94dc77410ee92c07b16893b5c26d1b9080365041b2beb0765f298dcd9d1621be3ce2578ff5bb7a0935196fc3a93a9f56a08d53308d5622aaddc45f9dd209bfbd517759e0b9a5ee57d78e4f30697beb1a6dbb0fe0f50445e93bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102ac4e48145909324553d22d5061b9f8858ed69d5965f9dd7f2579697b274bd8bf9ffdcf9927f583730aec119ef14aeaa70b93320e71f5e5e443a6abde92b7d48434052f78fdf6a5b82b59c67b08ea740554ec5014f2e3210d34784443eb8770c21d6f92bf0736f303;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28dbfd4da0589eeb528f5916b47639a12967aa9476a009dafce873bc3479e7e6c354a229f5edea3c2f500d131001e86501f2c196eecb12a56fa1e76120eb67231650467f74650e4df6f112252dd2e3eb8bdb5469e55fc95c6e2d75115d5b4724a6fe700f0567344363;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c84fb064c2f39ca7e82d4fe238a628fd2582e7757fe0a2f0a52e1d52b8afdfac5b378b402918f014dd801d347a76f047153d43e36c531651ca2515b2354f1ff909d67590dbc5f67a6d0ba347ee25bd994fd020ba867152ce6397de004f100d92be42577386d0184e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fad3488563386fbff52d1db803510b36b85faffbc794a48b977186ac91ec504055382491510c379241a0ee641ad85daf8d81bf5c6e2a75128f3ae5a0230ef44b5458b0471f2abb97a2018cc24747719e74c01d7a01a0f3eac111f07e61e3d97d3ebb4bf16391fd0cb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadf0d4dbb920e627d58fe6fd941c49d015325abb7583cd9348c4380f04cfa3c9f00b5c56d187b1908865bccf8935c824a75410e49ac643d4b114f1b089cb276006274b5aea3918cc709637b63d52df96891d782e33a953d934543c8947569b5fd3808b9b6d210c6643;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h199a6306b9703a0a883803176f49b5234375b38773c941681e7cd6b9653f3a4febcec94f3fa279f3b80923122bda561e94fe6d1c8b6727078bc76cbcb673cfb219c746c972369c694ded983b14c2b0dcdc3bcdc0e58cc637bf83611df3cdbffa8fb13ae1582d10346d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1954675216fd3e06d8aa3219b69ef90472663960ac79b1f59ca70284d833edf4befaefbc2aa7d8835d0559397c9d80659d63361b623678734d65afc4b9a277cc31f6712776a0ac287d89d8aadb569921fbcca60ab15d1f0a57eb58adc16509085ddad920efb0e98b3af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19204e2ca9511c873a309ef839cb24e2751c0a8030b51067d2c1e7e72b93058bc9105f163ff0a230d298d8959595e482b8b67d964a54bd33f0991737fba46a66b28cfa28019cb0be2f7e841c0d2c7e70d40187663a28964f488ea52d3b7da83cf3dd2b272d6f6b8ee7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8083a607b0070df79f231c4942c4464d768913a231d1249657b1d3f0c10cbbc128bc756efddc4d5fc6c267e2d21e30a11b4b402ab5e3a5ff6964da5b3f4d8958ee6fe4db16f39923fe521ce68be8e32e175f4b3fe0e628e1e9e139dfd2b6cc84c5e280647ba6ff047;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3daf76c6211c6fd1b46c8a7b81e526950022785a87fb1918c8899f10917c6da9e9d170a3b37c2612a7ad8d2a70af868c14ce953a7009c2cec841ad29d5ca5e6241cc18a42c8eb20214600353f5639f195769d3c0df4417fa30ea060f78a03024ceb57c4a6c0c21491;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120400df98654fc660d0e33e7ad633309e9d74874cb24abf74b79b6f5598fe4d3ff58220631b4aec788a37aec505153369dcb8ad478f6a79373625797d45e8447bf3b454c48e376804e6c258b86a2aaf0480e24152a4442812189c95f1bcd9b5c4f7796783226f453fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd688cf332df52a21c65e548a0d657dcd377a0c79f27f6f68223a993418f0850fef0e558298b3cadb2508f35c6188497642759ecaed014cf86aa7309a44157eb48824b840d03f897119fcc22d0805760c88e06d2601c1548b92833ad126b3889c30620c3bff3762b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf3324b0e65678a4fcfc099e910422c6f8b1c60b8be09384732c23738324873cad4c9dac319221660421725c7c64358deedb616bb2f8bbd81f3e0b4161afd0c9ebd11597faaefd26f3412de066413532f8fec8c1945bcaad7bf245ea2f4142d07934486e16800535d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19364f079c0705c3e7587c81618811310bd0389e238e725fa73e4f4254806a4e49c1539a7bddef1e4d463c5e588407e822f16f441f79a8629ee0fec10a087dfdd27559fc52e73784634a8f7f5401d5e20aa20bc9d1b02ed40d9514962c0897db433060ec975253b4392;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5725005ee9dbc0f20c8065dc9be87a5da4833c79106299cd0a7c63654fc4920ffae380ab1cff07ebf90e0ba91a72ab69fae7b68fb6a6829ab9a63f5ede18c6d829ce01e4e71389cc545f56a357d9274a3e292e38c741063ae053da4195eebc0e02e84d6c7726ffaee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6203f25dbb20f2a758d98f18870c37b18c503239221cecf37a332f4db58a087e3abcabfe5e93fd2089134c343b0a65429c5c3e048c407907b3d6a187a932e34fe44e7b97feaa0f4c5ad94f3f87edc8281897a1963f664d04ce8655d318b36fc96bff9426d330bb58f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68d686d59a36b4a69b4fbd37822cd001b8e65be4a66487bfebc69f5edbc29ada42c2e28ca20f71602ed718ec4ddc1d8c4b17308f76a3f11c6dcc2b5ec5fd421c9afc8a22b650d2561300deb79b2161e690e7a738cabc20e0ca6d224f7b0df6eceb347c2509679c09ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15aaa80c43a6dcad5169e7210c7b66e9e08105fc4dc8244ace497fa2e9f7af6b97553baa63236af449146f86e2d819c9dda3aa620a01e6e728aa2d4f60b80ba38d11479e400b1c5f8df244f0f5fe7c4e4a5ecbd38ad5ba276a12199dba297be1a24667e571007a7701;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9add790158cffe2a8cf96ce49f5b08badbe4c99e6207fed1252bf2df4fecc8fe059cb59f3eadd50c28444fcaf4a0fc9073cf7b7388e62d7c10db3809512b67b2b1f90546159c01977e8d91bed8e62aa312e7dd123598648964107927d613e5dd6679a375c459b5df4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8b99486df194f8e3d4cd04ff2e7167de4ff6f476fe68156e9322681f7a5a1db0dbb76381f01258f29525a045ffbc3d048e5e97e7c321eca31ea161d1ef48fe2479e6951befb8ce8f0f3120282edfb27c27b5a5aa0f4f40e4fa7acf45e57074daa745e38e7f3d80fb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10aaf177e801d1d45558289e5522069106a5cc8c722d720499e5d01b3ebe5f844acf756db71021382cd9445be8723718281efaff8e9351ccdc1f2326b0f4f5dd5b3bcf885d4d4ae960c7ab626e466f261cd458c2582bc5d038ff1f37a7f406600d3c0edfe5c04ff630c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcefe966f5c3764605ee102cd66adb8a33183469bc54419328077a4655bfff5c5810c12e56ef68962499138098bfe8669e6bdc62b49764515369cd1d55ca3ef72ede5205df7ee81ac8f439c2fce40826fa0f8980164fe9a091aae8e01d88fe7cade18c9a8001303138;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haafb3b8a9b3cafb10a6d596b0b8ddc89c847b9dff74e96a2fb45c0a2426ccc0447231da5c8f0316942eebe76e9c1a787b77af893814b6b1743169d65ef97f6dcf763c5f142c26b2561b543cc1156d722157bd59f92d83f62b0ca498740a50f0451475fbec2be95d278;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138d7b39df947a81409002d7b00d07070852255740e2d43bc18ae1171ae815dd2c18c18ff1598128fb6d46800bc712a87e354fe471a76c4c7880f5a09ad6d56c795a99369bfd220d1b16d925d060dd36a0c208c666b57723f8e087e45b2c38609ffca80bff77ff31cc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90f889c3ceb6087328d51e703543785fe77a3dc927001868b15960c2e6bb2249ac03f77a948b7e4258c39b623c284aa261724b717b87c886448306a4f4ce6b790e68974b8262495e1d8e908eb9f6e88c7fe160006d581df4ee05180ceb544543e302f01ebb39af5eb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45a899fca2c2732fb39d4185c46a9f21634c99a8a475bff9e892644d40f8c597cb66324df550efde120b55112a650fb8274d85f144111b41c4b2b218ed99933d095146887f3386d6523fc279d02ffa2b592b5ecb71640d328609205779687afaf128ca448620a9898;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed2dcdb7241d16e3db81c0e66afc73d82133af5789f9a4c12ebc786baa99a6098eb0504aef679b16a663c36011fcf313ceed1e651d9c0fd79201fab12f7360596bfb1c99d9ae4b8781b4e813218c8a93bf632c7382a0c0db31643c1aa69afcc4595857c35bf82e22cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5e133ece7e9d53376717c09623fdc37ab01041f78632d3bebdebbefec8d94a6d9fe8c5fb630d91d002582ba33eed9f80318ad56542ca1bb1cb665dd691e58a3bfeeaa2112d1ebd9559b6b3612186afb67aafcdac7f441bc57ceb22ddca5c5cab8dda5d42dc95af737;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1380fb623d66ffb3500c8bdd8e07b05fb7915652dcc04bfeae8f9fbe63686e44f253a626f0121fb4608b15e2e68bd2ee28842d3009d1090c97647f4ed85bb2bf36c0e9574ceec4b6054925b24e758af1a7e2d1f556e1654cd7dc428f518cb364c23bf943f5e17645de9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d00947868ecb4f0d11ded8e8656889c27112fb4ca8820fc3e9d1ebecdf9e818952134fde38ddb72ed2c716f86ebddbdb5830bbfb0e47f6844ed714d454bd81fbd17d8081a63c3728265bc11e170d9cc55c6fd7cb33082b7a0c8fea9765ffc25e84651700f041e26d8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a964cc9e09fa1ead3fcb46270a92dfebae3214fe62a1998385342175f06d2a97f63cf15bf21c25a934005c4809af48c37c1f92d87863099a6fd8dc7e52aaac3c97969e7aa87e51342fde6d0c5d54ab0debb52b0a2cc3502a0f54bb8b9357366aeb69fbf6d47187f9ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h772797be7a7665fd60e1d72ee7572daca261342b6f3ec3b5f4789f3ddefa5753733ec77c53dc3ace1d1335e1c5dd44f034ac0840edfeab2405116343dfea5613bb73c329dfe72e0322fb698d648b8ce2f5147cbc7a9f2e926eebacae7fb2badbd72dc402bc96689d05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ec5daad9e31b02ae572dc66b66824243b4797aaf39efefbf9c0bd81d749e69c7a615121951edb0cbaef36eb903a1031da3ac4ffc658199cc97b2eaf5115e4b356c33bbe4f2733ff7f2b54f1d74b21e294ed6db3a9ff0f07863a015bbf10e6d7d1dbd5c00fadd5392f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143a3046c2927696bbf284795a25ecfb726e69117521e947f95ee679816f2a4da36045bb970e842291f03a3a8e2974a07cde65ac83efb85ea6e4166340ab02a780bd5e4420ccc5e53581a772388fc4ef8f82e08f55f5b889ccd88c926a629ebf61fe43609c930a5162b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f1712cce063f7460eb17c86b4339fe11292eeb6463a8d530a5ee35e449b3aeda1b9e51ea946187e6576a5738abf648de8c4315d31ca5315efd3d32e245984525d567e2096f10ec1f00529462c30703d8ad2b6952292ab2c18203a6a3e54c86b6e141a0b6ce9dd146a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123089b8ef2e532c29b6864b8f75133ad291b9ef55c48ceb83c830c4078494f85c09f6e9acfe56ca519df012364c8fc32212d5b972e39cc28c572d91c95500185c2d9308fdae80554ef757b14b8f1412775d2e8f45f6bd8b967e364cade5e62260bfc348a17eb03b0ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1685f8bba8efc4fb1c0ad5f9116c09480fc32077b92d928ba8c68e84b44663435fa7d1cd9b5b12273e5dd931884667c3808665509453aade8a52cd8b8e1a6532ef1fccd0bd5f857ad1022997787c7a129f4211357f596cd417759197c0e18ca2e6ec1b65c950ea7f411;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b86197da01f7768e01a048493348ac5a3cfd7202bfae4237e76b82ddc3eaece7428f08573574c56be9617411e25703393974263a6ac334ecb211ff356e77f86b1bf55ea1d2e5890ded4b75b45868dc08dbf02e4ed38a635563971ae2f78a43dc8c3a4096e3e5770c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c666a67fbda5caf9fd991bf7ee1bfd31c513adae498b398193293f8ff351357da915597b71753d940fc3a08fc9dcc449ca3e778e31f15e40fda218a7810f019c7cedd41fd5e443d338361ce6cb5fcb5642bbed56c538824dd4a67cf98ed3d4a1c227057b9b605b978;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0f3e74002c61cd20ca25f89be5a541572b5c34163720a19941aaef47d3cc738f45feff281828f408e337908937be56e29c21c0ed46bb3bb19816f489392f08f4614b4394b0bd425b4079d62e835faeaec393ab856c4b48ad6137f55fde0f1ee08096bdd267de13966;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d24c2c322f85515bb61c40ae33b8ff5dec4b00f5f1c1b976ca999c1e12fb3fcfdbc26b364844c6a34dc785da1c8bbce21e2348726f189ca6fd98119a7764b8f42d1b8e13ebee4a63f6828a2b9642c5110b6047a973014df878f703cc1c6a312c0b500ff0d570b31eef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15161ad1475b2307f5888e917990810a2160d751e558b09429c0bdd6d07d03d06d85e2904cec35cd7769c9cd773472b74392347093255b4969b16f122afe02de325dc00394817a51f6b6ee6d56ed23f0107059f1191a92af08650605171a1b10851e640cef9b6bd3cee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cea14d20eb5b92bf1034683a80538e5c60cce9eb46ad703a15f55a690804c34f97485a4b5dace61ae7cc625c02ee21eaff7cf849bb72b74f18c89f99c898b54a037c368fc121722d1a0506035994cf77fcf9a376f573bab53e41002eaa2bc4a57cf3c476f23b54966;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95daf431c9521a5a61dda0ed5bc8412ae79a77ba17188d99870ab7c3707d354d58b88d974769a60d2ab47d0db2d03fa4499764841bc713af227cbd3acb8b0373a5ffd1120cd704fbb0730da1197ca509c1d5d476fc7ec50a0e6dc9c8115b840d521ae5d602dc60db1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b0ef2dca50eb0990b7661ed7c09ada6815c1b7140e5eb1f266557ff65926e5fdd445844007cb1b3c6c85c3092645e596ba626c8f78783a38b39d9db3f08ea5c1d637f2de5264449b073b96cf202daeed08ffeebcefe3e25f552ba9c91a21f6abf61dbe2d342d0be80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0c6f53ee861b1d0e161265560c96e8df569d01a749039003adcf87c1f8db0db10911e533a7aac11ea21cb9795287b0ada669fd306ece78c7840c6c4c36d480548bb6f0b406bca56d3dde8229c0630694f5441e5630555364f2174b9448f2600dcfbb96d97a989d440;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbb15766189662eadbb676835e1012c905cb080b0ca6cc6ad27fad499aa6d12b248b67fa12df2ec4d9f824c1f8c8ad9b6221cb0fcdcfcb4b0617e2b55138956f9e0e278c52ce6adc12662932f4877482ff08c28ebe2d643841e0606bffa7926a0f78328e8f4b62a724;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82068938aeae5c04eeb57a0cb4092d1cb217641966660809ea63fd7a5ff52a2139902d466acf1cbf2055af14be150639d19eeb358dac9e61636f6b6227ce048d99075b9de2a5353d1cd802efa5be66aa1c633fe390bde1d030c1a043c0f712632f4615eef99f67bffe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd061cee71ac07f1968219457103524d19657a0140f3d581d42a9f2ac82d9ed4862356ead0dd9dd84dd99c95281e4cdf51c0591c9de8b5d7c75d6eca913d1199d7fd3664b8634178927f0fd6515f19382e75a9380233cc8f08bc283934549d4ff0ae23b694b9c6b88dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86d6351d06af0c6f4fe6908ed2fcda4bf18710437eda8b59d8135c5f7cd96d18e607fc9982815a38a1f435f54b0121b6ac0f23e9218d1cb4cad31fa3b87114eef7b07e5052a20d99f6d6289052dff3cab207743cd6c8c27e8ae2d546a5b0e9954d3ccdc01b92a6f5c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c50f92cd316d9833bb2bf91ee3701aed14afeacd308220c68609fdeb6df5d91ee1f4380e3f0854c10bf4ba4a0e2537b0a8198da11d6019c0b909679f429529fae60b410e493f0e21cbbc1e8c591e203f0d812202fbd0908300022ec44812e19980b04229ee16b67da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e46195f302f1968bf8df5ce3d8685b128eaf42d9d5cd08d083ebad4d5b746353aa50bfbda6db8a7a3e5593aa09b4410a6df1910c707bef524e748c47388ba6bfa1c1d773049163b2365c583a2a36a9732c1ba8f6ac2d72528482dbca5cced6c5eddb1d3625ee51405d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1528d5257aff94d7b9324e5101b8b24f96aa51c19dc943345b80783feb697ac30de37360028b64d377c1f98d3b603d72eaa645ea545f582909168e56705e331d264f40660ad1439d5dc9b7fa19fe7e104ef703a53230a6f48b3e3d30076c793807bef16269561f18d16;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2adff7b3fee811c7cd170af90333f2e6bc52847dd719789e54633f9370f07866655b73b068fd4371d5b40993c53ca0e69dbaffd15978929672a7c382c685f4b4707ffb6041f3f3fb493fc95bd67db9a8c0c5c586d08ded629513504ff41d7c86d8e27d705e37d01de3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47c582cacd89cb9cacd6853dcfeee3a1dc144279315c9bd9bff5b8f1824e3c41b140dccd553de89d04e62493bfbd7e4e47c212b40af6e166eb6e4bfff501bf2be2c5060ea2d72f9baa11549aecf52c46108ce3458d02fd9b68d0aefccc1e0b0dbff6e7461f11ed9bd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137dd38e3158163e517316b2598a7241dc36e1cf9b83f99a941508412f62bd958ba974f86e2940c0414a268d7ff1b3cc62a388660aa28007a6fb300f77734aee4b4165ad87ee3be7b740f1abd61d8508f5069b93adf0d608dbc8037fa2529c1c21f17c7522fe4987647;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8e43be739d67c9b71aa432bb4de16388b034ae0fe3be7993e344e3bfac8b150ef9120536f7850c29778fb2e06c589043abceef91d91a3dc3447f4bc83e8c9b7878cb65ca4274dc084a656bf0efebe478780e9318d168109f1d2dab475a984d08ab980942321de0f51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d60c2497d7067ff4b06f6b17b903a89c6779bb6372308a91c0076f249882370068ccc27c2e235655de462fbc364b0dd6142ec5b3d8214325a89dfe3f690e09c70b776810f156f4101ce2fc58354fc32441bd0f390b9bad14f95edebba216fc8c495408de01ccd540be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aac8fe696afb9e0b60ae38074b7a7f263b2695f8f190fd068460fb560cb5d6bc1d369040f17d48d886a07d23721ac1a7332d74f62f6203b3f5fdff0425f8a756947baebafa7dca7a8f761eab391c5ea9715fb5a60326a20c92d3dcc8bbe482d7810cbab466828f8ed0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9ab7664fd69f8ad817043196a8d10fa6e2bbc7308f84dc6c73ae515c8d578a994ef16731b0b5ecacf5701940c1411bbab7cef8737032569cd7ce21a3fa4ec37c1b1230d3f2f06fbebda10cf4a8dc2c212488460b75104b8ae17979fd388f55101307f9739bef0c92a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd4d247d6c839aa80baea5d5ff3278bdfc786d0c0fe9c6b3fdfef713a1699e8cebc584abd4019aec4731ca7867ebfcb1d9370c13d52e8cdf56e6accbf804e0c771f7605913ffadd4355d59186a9c33ffd75c4296fcd1b4ddc1e0bfd26565b137dea06db61d2dbcd07c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f3cf16aae762b10a06ae1ad4001d4733c340e1adc6bfa0c7ca26dc79d66533b9d49a6c227b316ea8d46635e0b260c2a3ebfef32c4b72047d45d2ffeee7890d5da2084bf19a16b6f1312eb779ce7752498e6e5db8a95c39224c31dc65ac4151d935db0d8d95c4ba169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170bcb9a3fbefd0a93e9e024c91ea43c1816e72e6b5e033154a3f7c0d54fc2445835d58e3adbd2c98df882fb0813de9ae304a735c9709e8d4560d6502cf9530c2297c4552328a2fb652d1575096d59254799baefc28b361b127a518b5ba1f398e07643b06f2f887916b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c13e90a5f2683ee955b1f070e69da128e4b717c5feda16c18928ac8584df3587a629b6b7185b7891fbe5247d9dc941532bc3658060b6d065004aed4ec497ad04c18a597b5e55c775d22bbaaadd1bc386aaca2bd24ab83a3c0efb22bc1110df1f9100f9735dd554447;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bd87d7ae3a2e05e5bc1ae31eeabd2327918bca329d6742d389d6ea04c421e3c7316dfc0363f798633419e85e016210f3c35a619ea6b558b05b0ddfbd3ce03b819286c00edd2475dc181f3a46f6effb0e49eb21742ca99e692acd042870ba9da56ead37df6d2553942;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b91e05ef919a7305caa06885c773c01e68d151813ed7f0cfdc45f73726f94622bf9cd07580afafebec2b6467115203a37167a8a13a1492c8f5ffbd062659bb6f9ce60d422b4eacc6a19bc3b98c1e4fa937861606edd5ec97f7bb4646fed9f78287fdd494a252ba29e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2486b7f5a78803a4dd5c343d4145affd54115acf1e4c58bb78f24a3269e885994ff8e6209563696a366b96f13e71daa7b813399e1ed7dd825bfbd45a161b945e7a80be1b874c82ab733c8e72b99fd05a926aea36ca3578160a3a3659cff7f89f62326fe7bdde7fc1de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19322f314dd2ae3a565da660cc8ea039e2f1831fb2ecdf1c05229b50d2558fee16858cabbf975aca98d25d6fa7e9a5a3d08b168925c238d152da08aeb4aa6605cbef94ab4935dd3e5a9d1f397cad94ff60fb0433f4d4f9aa887212392264710218a864cba27e8589ceb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d4b2b7ee2d208f99db99e0257f201ae9c9e1a4c2d19845619daf37a11684783b02a83890427768be384a65859ec756c9fbc3b9dec8b8f8742a8bfa8464aa56d315d35fc7fdcc94b0e65316c6ae10df04de45895d00145ca5d7a85eaeb60e3a1049b782915addf55f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h497efca9be81e1530255e038641f8150355f10d1dcb1bcfccb0856654cf57058799e4142645c4f3c175634613473c41e405255761bd55f7cc27895f99e22c9784f0584efaf432a7e0d00f3c4e80e06bb5f0aad788b1363fa99b653fdbd2940126b46859dd30f31fc44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47e6e5e3c21d4047fdeaa592bc94b54382a8be6ba66200ec1085c46cdae7b00e7275c5b2c2cc8b89290c45c37d50c3cdd8d8376ceaf24df5d25aad1a775399092a9a143811b453862d198c15d9c676c0744860e9bca7f63a4ab21fecff8835882aa9d2fe9d1ec4c19c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c577aa28aefd307162c0dd832e0686577e67d17a7fcd8ef9b15fa3d528b59476068209eeaaa4b9ea5059b7f6ce9b4585f394e0eccde92b448f15aaa09fa2b4190fd90a5798af3e10fcf9ba5745fc578d19ef118dc4e96c01c7f6b70da2a9e0374f5412e77929d99d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h671f411f606319efb8ae4049fb7bc3397fa1ab7bd7625a78a0de5d47c983c894d32faec8726d7ad41f48992fdf6de28e53edf27cf71d3d5a3fd44bb6ad4293be2991f4b10bc7d04a9630453c8626843123d214b1047ff7a16187b3730a4ed71d9b2e0a34f608ca2847;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198b6e392579aaae91808f3ad3843041e48597f3e889af14e82a44f38beaa023d5cd51bfefa3f571286abd02a45c10e068416afe8f23eb1d47544b041a8af5bae9705825ce054a7fc0a838702ec739096b2360e150d02aa644e15903049c615d8921e3b76afa5f69be4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c8f631c7fbd654dc8ac9d3b28256cca6d07d3f1b467fea7a7e4bde37d7bc3ad138341e5ba4603df511ff18d2fd94455cd3ae420b19d631909078d32e480631eae370c005fe34ec5a683a8270d3a04ed90082d5f5ece27377758f19d002e33f35e06942a8390988130;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33e26eacdb97f587ec6ffb4b8f49270ede5bdcd681554baa22642b4368054c902e2db6b914c1dba1689f31c8e3ba3950ee091ce9fa97aae7152742be0e51c4b35af5bfd113e8d87d1eff4c050f5047020abde857a11531042cbe4127ffc5d9377a8e462405a8721881;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6331758b3bd9719c0a5c1cbbab5d0a1e0a8722e4e64e7a3cb63a327d09cb94dfbadf7fced11f86d25122d1617c54bde7ec6629ed571a164569ac013fea818166e3c34ad5707019b487ea089fbee6b76f8effb46c1ba81036745183b9de009ddc9b8a1bd6e36c9d3b74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5204c2259e8c2bfd2a75d0c3f4e79cc8dcf0f6bdcc95fbe530308df46eb595e4fbdf55684d27a20a9b7008b2bd80cb84785395c6d0a15e6f04130d1f67b85d8c41de9da909114abfe1bc8da507af3cfc72f04c3d15f1ef9ae9ffe41f37894aed419358b121a9126bba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150baba74782926796a793c3a0fc70450ae786c6d3c2e1559587ba594cf3b7e2fe1476f622fc978bbafa803368ddbaab5da2b852e74c1d6d60b8d6ba35e2dbd692c91c7032ef12bd9774e8a63c83d6bc622fde0c4bf825df93ad202db7341718df732afb00376c362a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0be1a043b6417360709835a16aa25fe60edc44cf1aa746b86b8f304443f82132eccd6b78acefa13d9ad9aa339a5b8f25c23978eaf6a17d72a286e7d1a9e301b4680f92666c1325ddeda6357f61e4d04b7f381f0acbad2a5ed346a86ddf4c63c962f0a89ab3f191f5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f91f3e253913b7720c6083aa8d01b7541ee70388dfa44f9d2fab4710899f124330daa1ac1f03f817da2e2c9f4c7be1984cace268e1599770cbd0e29b187befaf6efaeea150308921dcdc195b07da3c8032e78c614caee9937a513555a4359a9d3597a77ef27ecf7869;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e087c0a19472eaf12d65914ac505bf5db64063056fc4b4a4194fc75c7be96f91682c8cd793fc48184d9bbd71bb6f5eec821f68b8f3350353d49b9fbae2487ae2463b52bc804200cdbbc7e7c3a28f256abda8f2021b6fa7bc7f0039163d1f3a8da1e34c4b8eedc8d78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cfbae6beb17b66d4f17b1223bd496a5800dcdcf30eea70e01c3ee10515232636d99b8ddac9e3067376b98dd8ed27755fa3923723502a76ab8302767bd00d1a37bf7500aa6304553ba7fb872d957838dfac4910836c013e3ffc9d4e68d42d7b7bcc2af2f6e3dc8a182;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a571d8ceb18d00a2441f772eec2d01949309dc465bdb2d42c3b671658279ebbdbd34b019fdf080d239434c2dc67c7db32943b9481fec57ba33b611ff6ed68ece469562374ce41676e721362e8d4bff5c9749c324ed1ab5dae7f7b8203bd21be88b32b799082eff59ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb3b3f6495293e02b0c9252a1d82977b2d5a08a3f5fb72b0b523bc1309c6a2d2d788183563c8a9edb5fa3f471dc4ba6b18ad1b3614db9c26e4994917b3aaf8a4ef6cfb5cc7db87c5e2ea77a5f7fadcb4ff7a4d0913f9221b3f244536d0bffac34fa7c3078b2f2b0a7c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbbbf94d899af3eddc9dfabe6c2b73ad07e1bb0519416b104b104fdb807dfc1ccca1f2cdafa774ee08083e67b9c57f910035576cdb41b1c6d68b7fbf23b7a159e2392d5d82a7213ebd8224c921292e964c8d0976e5e2dbf6d331e770c470542afad3b4a8b36b15f3f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd8f8578a44d1e522fe80b60a87437c2971a2ae55d5ff4ce84ad678d4cb59b01aa836a5a2c950dbc3cb4e97a4ba509d464bfcdd7613ab8f3dff3f1534c1cff9e3d5de7bc7f7c3b5114f44148aa64cfd94ae01f277b3b0a72b033c59b0e9e8e5d123eb7d4e0c5bb8ae8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee9c8847c01af24a0df3231bdba9358a1f2d51ccda17cb980483ff070410293a583c02acf9b1d250d1642adfd1cc50fb6f93a4efbaf181532ecf0b735f7f206251f609b3e2c5758c0ec3f2ddbb6cef7f0cf608c07c64283b5d15681529ba5269294ad146ad64c3bbe4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df14c6eefeafb1830266e012def650c0fd6c66a280592a6ee88a2a5d78516df02ad9fcfb48b0cc61ff880467aa2b4f47956d22439ae7e13c0bd1e071cb5f51501ef59364509dca75140d7db237d269769cdfdaa45bc611b99cfe3e03159a95ca838b08c7222aecf6b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d27894624f93f178c1740c097ef116304866f54593c82878185caa609ac0b240140d8bc5470eb18765f67ea3c119188cbf2e88e17b17fb43ebd71bd3f93be666fa48a587eb80ce134253b743be37151f776fd191789edf83d107fe6076462bae0efa3ce0a2c887e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e28cc90e025e45acb31a5b93e187e44c1e5cda0718a8545b20bcb374e4fd2bdd2bee90a07e5df2e65a2858d6816f70c3bd8d5d46765252871a5306b872f40448d0edd47ecee7ae345772f8732d5b33cc892e151fefb1cb8dedca18a5c76df359d93df9a68bfe648358;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76d5251f1ecd6956e3edc4dd27b820487f5e36c3e018fcb8dad63a677b2ce3e2a0bd9c86e84df26b51ac91b13bb3d7ad44084403fe20f755aa7b806db00e041773d2dde9541b0cadb188c60a4c13abfb4fe2e4818e88266f9c246766bd920c5f9f90dd0288f3f85c33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaa2afe984328fb31fa5552770d3e2ba0c297a63bb2e96e25cb64bb6e4feb07dd8cc000f84c45f50139907396face27ffffd84fc3c4fbc207dc697b6ea9d3cf6eb16513f86058c1afa5595c678239ee2895116f90628fab834e824da4cb63c1373f986bed1ba5af169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db93fac63d67ff08f9cc7a567e6fc8b365200a9f096ebeee7df7282b3bfbb02b992e605cfa22df78cc3ecebb149f1a39db4f1b4a0af520ab58353434ae802234ad57dbcbac94431d16c8e5d710bf7481f6fb9f4b4ee1a54172d53eb51606c0e4922444507a67af60cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19eb531c0b334239e27967bab8aa27c00e03b756d2ad44dae19fc34f775c58d4da36c95b64da751a10b6476558acef6c7c33113a6f0665c87f0c349701e11f2587684b9f18d0d9f691e56e71b528bebc8d3d6cfb5cad6f9982b7668197476a85bb5f729f68746b56f6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18dd83b7db44ad11f653709a391a1fb3816db2bb01d91e814fcb587077b87de6eaac1cbbb74c3282fc0f2a160a8f09c904cde6c57ceacc1c1f17b14656cd67457a2db5f2da2d78c2f9dfaa28e9ab7341aadde39992e4b08e176ae16c89cb4ff9bbd313a0db859241be7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175a1d5e5a72ea5c7825311bb616214c1e825a169e9fefe3b6acb8e3e2a745a4a2d405237f82bf9461b0bfa400b32669eb5021f6e622608891c04a64b11d43e8d464410ab01f809d004464d6f24e13fef9ae8dae5b86837112081130538a6d4f3c63b1a228bab03a491;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6026091f9603f10b5460226d638515bceefedb801af4de7b3d4cf9d8589edd217dae190fbf8dd5b333c7ef99a78c35b1c0d07fb78a24cceadd530994406dbe60624cb7ced6a2e3f8c781a8cd5c55b390a3ee36e176a84a1415a8613f88b31df76901ceb52a3b444765;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ee1c5eefa9394ba1d48ac825bdb7dd25f711e4de697a5502818ec51127e435295ec94fbfae7fbf8ab71f7816031cfd43fdf6bdada54ffad7c79bdc09738a4bc941dc68ffef08869c778c8e3eac16aa7c113e5cca28cc568f9292fdae6b9e08c16b74ede495d66ab59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8b0e2f16297d736fbec3d4c328b150ecf12847590fbf9a91b30aa9e27188c38bf4059843a977358f42b1fb31dd2428db7cef08531292a1f2f0bbffe4dfae165977b751c69b3c38de5cdc75f794c6c24d6d63c99b91703a165fde917290c478d8d0621bc6305d991ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9fbd2d45c8c21f954d67ce70e652786a856411ec429fd0503cfe2d64cc3e319eb1340a6726cca7165aea28d2930a76bc4177689d44cd49613f60200dbb894c52245db62d76628252c9ae1cee5f604af89b925ab6067ebaef3289d2d3091603518a0f8b8516ef7d08e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbab7dc68b0fb44cae7493c8e3e01cef2b23e6d2115d0cae6a45c396668084a0d9d66c41498b97ca464faaa5e91ee6e78eee2dcbd0e20df8415f699afc49c24671342a39d003e3744d329077fb90ace1085c1da561025a0d112627d31e14a66b237333855c19f42b68d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a83f98b707b66fb6076c81fd780b871fe971911f91b15b6028a8257297b2fa8524e582dbdd5a4fac82e89fc07e06d9eab1a3e78c26692dca03946fe93b63a06440d7e1eed3848949dbe09cc28676de24b101e4792da24bdb1b15c1b4fbd2699cba9432f2be0258d2b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc179f49a027efe2102cf4a931d9ecaed9b9c57d6d1b6546b62008e8bd4e11247336710e44a6c91245c77ba4ecf8c24f8d49ffb3ec0a186089eaeafa378e2a6d444a80869ebd20b4ae012d1a4009aacae451e3282eddd705b8c93e23027c7d949bd976773d7bf846245;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7e6ff8bb22b248ccb553bf3ccbab621835e27f21438017acca3967f1369e13752887253bea0c220e3a47c96af13346a943cfa8df856919912f155510e9589816b7f1d18c65bf23b86e7cd26ca7b920c4b506afbff637f7cbc4a41d7875d495a86fac92fc2fe7e28e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7584b3f1f5b114eadbb75c7e78f2b62effe1bee5b750d4808af7618d9b9730552921a3e0b9ef5ec1fe3553306460b03b3a8ec137d9e19deb146542325bbf20c3c134dde210c8cff087cef7f3683bd41a48c203671c04431015d8ef2e357fc619a9dc1c1575cce29e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec1864a98c56e5fd569db04aad44b13cd771e22d29997545ee7fb3caaefe825166712df85386231bdbf7a078e889b0850e8fe8709dd763254b937bfdeae48fe78707847714440f338ce6c4691e90814b3dd93439bbd8a12a0241025b2aa1b28553709ad688da1ff2e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119ba2f39d3574deea274cb990f485ce01d97437db4bcbc51d74e1a8e0401281e04f822f7100fc0e2a3885d054a4c698e8b61297136e538decf159552d754925f21697cb0cf1190309ee00291f53363b152417b55c884fa747bbc685663f118981b9ee5890cb6890b04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdca005afc6149d6c3958f9d5e1b1869300a571ea206837b2c91a0db660ad249ae701c4ec63559afd0b280b5dfa0a679360d8a878c00af1887b009ebfa3287c5e73777a9ac12a77ba976568520b47783424216742bf39a1db1b81fe33410b7abbe0b0d13ee2ee25f927;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44e0011f809b81c52089b6403c0a62ed64ed437099465706a8ee44a7c414e17166bbee0e8ef68faa9132c4d909ef097a5ac1e987c231894dedf23a05f227037efc22bc5806ffd2deb9e12656f31f333ea1cd031b3417c2fc677901b6b2f627d6a6aca7b7932bee9123;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be8c9665f3bb15bc5d7426c29fb90cc118baa64c5835f2cee8964699f2ee00f7f08679bc2377f5d2530f383fce94f504a3add7036595fa33f813160beb7cd233722fe9a8281d9649b6dafdb087e015e12c37a5eb4f0d70773941d877fafafc223eba32ad79dc0f9a05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa07a13208ee0130511f5b25d7c89a4791bb4eb8dc807236b2413d4a9f1071d632c33dc03611b970e0fa371ccf79847802430b2a5cb4e9950dfc2d0a076954ca916cbd8f5d3aa8b666425a2cb347bf0b7ae3003283c3dde1e433d2f1501b308a8c91f2b011746da460;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d9528a897ad116cfe077e20044642c37ff0b2c886c3395691725923e1bc7149d33f7054e78b4c0cda969716be90ad5fabc6f4cad9300d035c54c7dec2abeb53f220c28fe91825b8ca295b01ad9c48a423727c1a1af641f6bd7c0e514697e510f716249d220620c5d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca0367481f53742bd9623c23546f2e8b6d5061d6a9e1ef5929b8523f25b9674f26ea88e7d4b80075d3e5c54a8b9e85da75b9bb848bc4f1fee460fda3a9f793721d66f215acc7532ea917d7d3cebb7065c1b35baf6d89c1e2c1fec42bba486ba16f2fc381d83f444596;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h222b81e637ae1a19cc483500826959946c99012e91060c8d5ad5f1c407082219facc2d1618bd4baac6bebce958471c8fe5b64f4aca2e2bc90a055d58ae6d367f70d82cae2400748c9159ac1171e83ee789bf08318edf9e010722acfc9d13f98a69b8343134b9f3b9dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5340fdbf7ad883094fc73e43a0d18104ebbcbc12513595c2fa04e63a9a22c3aba98d68e2713a67558643ff03e3215f96f0da5d31808f3e02f61bb5d2026247b76da557b26014d13df37056b9d6670d0fdc2b53c160b77016f1c0662244230251b92456d8467be0a44;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c2069cb87cf7fd420e4958bd42c9ecff8fd46cb9244b042f23b1469492afc595c038c52fbef724d48167483934e6dcc853ffb0fa84f6daa10295fcab6e3a81955335fae71a300363d08c883862123ec3e409641a3688d0fff05bc816c78f0c7bb77b26f6d3f0bf143;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd637f7f83ecdae9f9c375c3054aaea500ad111d4cce9b9056fa4e3a3450f973c5c9fce9875e5a0b847518271f780bfaf5fae89bb7b380f23c3133ef5fb01de5a8cd860e99763f3c5a7b2da649de67c9da86913988ff2cad2dfb362f93c80784db67181622ad2427652;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdc188ec8063b20b83588b70962567b0903d144c51f7d4d29ce23ec9f77e670c93611c61998ea5062a25c84c72ac69c8cfa1ada81d9abe7d019357575a752daa95625c105e8462923e8a7fd69c49ff0ff2da915af35eb841f909aa9c53ee1c47eaa047682f40f7980b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14be58dfd01f1dbc2486160e7f7044bc16ee5f6c0f5af96f2d6ba6de06fe8c59a4871fa1752ac8bb0332ae92047d5a591c7b436e8e4ad928e02695a3ff1a0c581c665f24f32551f39d857bcb26447b05ffa9af422c5512dc5285e809f3e507eb1824da821acbfc2da20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8f8579be2a42f0de80bed77cca60c328447145feda6e86a7facf82c0501f11a63e1394bc60bec1fd7c97dac258fcd7fcd1a5d700cfb7ac9cded0a6fda5955a6d1c33f6bbb3ad258119dd4ef348926b6d5e5fb57702039632894059234b19fba2d2896737d6a49604e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c91821a506639fe4c31514b53d2fee75c2b66c94aabbec0bec67108fb09f004d99aaf033d7806427249b044cecafec3c9d26f82b59a2201a069788e2580c51b00ea363253bc55b7264934bcaf9870d1bd5767da754755fe6775b0042d720979451d5132436c4e69a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha235a57fd8e5c21cf815b0d95edd11176d43c1901cd38a4bc5870306f26e5c0d9990f711b4faed8f2c19f9749b38fb62683ca1ca7cdd288bf085856bb2154898f0cdbc1f91f5bebc4073d4f63d4d763072719dea8de69508eac4242aa8ac3c9797f6d0e107acdf9ea1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2e0b3845eed4d3ee4f1d021853068ef6660c2228873d18973897ea2eca9fe0b237ff3dcf294a054a9aafdddff2b0574cd549156cf89d68f1bd062ef8490d9fb750c87181ee692bf4c987518fdcb04b259142e6cdaa75c6244e77505b19319f666f50bde6946a9f2ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f063de34de16fc0bcb00abe02dc9c590b3e95917dcde1510b220ca07ade98c3a22d3b30441418f86c3ee8e2d2cf18aa0f56bee4fda1d21ff9950af842c2d180b442c3443447059ae42b5a22a4642beab42665dea7189eae164571bc34823e3be3a93951955423eb2fe;
        #1
        $finish();
    end
endmodule
